module dtc_split05_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node14;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node23;
	wire [4-1:0] node27;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node37;
	wire [4-1:0] node39;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node58;
	wire [4-1:0] node59;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node65;
	wire [4-1:0] node68;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node91;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node99;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node115;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node137;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node164;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node171;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node186;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node193;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node204;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node234;
	wire [4-1:0] node237;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node242;
	wire [4-1:0] node244;
	wire [4-1:0] node247;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node255;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node272;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node287;
	wire [4-1:0] node289;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node307;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node331;
	wire [4-1:0] node334;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node365;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node387;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node397;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node403;
	wire [4-1:0] node406;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node430;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node447;
	wire [4-1:0] node449;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node461;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node474;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node488;
	wire [4-1:0] node490;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node505;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node511;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node528;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node533;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node549;
	wire [4-1:0] node550;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node574;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node584;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node600;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node631;
	wire [4-1:0] node633;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node643;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node655;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node661;
	wire [4-1:0] node664;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node669;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node682;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node695;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node702;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node735;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node747;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node763;
	wire [4-1:0] node765;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node794;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node813;
	wire [4-1:0] node815;
	wire [4-1:0] node818;
	wire [4-1:0] node820;
	wire [4-1:0] node822;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node840;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node854;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node878;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node887;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node897;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node927;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node953;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node969;
	wire [4-1:0] node972;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node990;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1004;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1032;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1041;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1048;
	wire [4-1:0] node1050;
	wire [4-1:0] node1052;
	wire [4-1:0] node1054;
	wire [4-1:0] node1057;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1073;
	wire [4-1:0] node1076;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1117;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1124;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1171;
	wire [4-1:0] node1174;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1187;
	wire [4-1:0] node1191;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1202;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1211;
	wire [4-1:0] node1213;
	wire [4-1:0] node1215;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1223;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1254;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1262;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1274;
	wire [4-1:0] node1277;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1312;
	wire [4-1:0] node1315;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1336;
	wire [4-1:0] node1338;
	wire [4-1:0] node1340;
	wire [4-1:0] node1343;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1357;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1389;
	wire [4-1:0] node1391;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1415;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1448;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1459;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1537;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1546;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1555;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1564;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1590;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1605;
	wire [4-1:0] node1607;
	wire [4-1:0] node1610;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1625;
	wire [4-1:0] node1627;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1633;
	wire [4-1:0] node1636;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1670;
	wire [4-1:0] node1673;
	wire [4-1:0] node1674;
	wire [4-1:0] node1676;
	wire [4-1:0] node1678;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1691;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1697;
	wire [4-1:0] node1699;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1721;
	wire [4-1:0] node1722;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1732;
	wire [4-1:0] node1734;
	wire [4-1:0] node1736;
	wire [4-1:0] node1739;
	wire [4-1:0] node1740;
	wire [4-1:0] node1743;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1749;
	wire [4-1:0] node1750;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1762;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1771;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1785;
	wire [4-1:0] node1788;
	wire [4-1:0] node1792;
	wire [4-1:0] node1794;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1805;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1810;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1817;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1835;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1859;
	wire [4-1:0] node1861;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1883;
	wire [4-1:0] node1885;
	wire [4-1:0] node1888;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1895;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1907;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1920;
	wire [4-1:0] node1923;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1940;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1947;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1954;
	wire [4-1:0] node1956;
	wire [4-1:0] node1959;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1982;
	wire [4-1:0] node1985;
	wire [4-1:0] node1987;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1999;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2006;
	wire [4-1:0] node2008;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2016;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2024;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2036;
	wire [4-1:0] node2037;
	wire [4-1:0] node2038;
	wire [4-1:0] node2042;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2053;
	wire [4-1:0] node2054;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2062;
	wire [4-1:0] node2066;
	wire [4-1:0] node2067;
	wire [4-1:0] node2068;
	wire [4-1:0] node2072;
	wire [4-1:0] node2074;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2086;
	wire [4-1:0] node2089;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2103;
	wire [4-1:0] node2105;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2113;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2120;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2128;
	wire [4-1:0] node2130;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2141;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2150;
	wire [4-1:0] node2153;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2166;
	wire [4-1:0] node2167;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2178;
	wire [4-1:0] node2179;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2187;
	wire [4-1:0] node2189;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2199;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2207;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2231;
	wire [4-1:0] node2233;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2268;
	wire [4-1:0] node2270;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2282;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2288;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2293;
	wire [4-1:0] node2295;
	wire [4-1:0] node2298;
	wire [4-1:0] node2301;
	wire [4-1:0] node2303;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2328;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2332;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2339;
	wire [4-1:0] node2342;
	wire [4-1:0] node2343;
	wire [4-1:0] node2346;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2360;
	wire [4-1:0] node2362;
	wire [4-1:0] node2364;
	wire [4-1:0] node2368;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2376;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2382;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2388;
	wire [4-1:0] node2391;
	wire [4-1:0] node2394;
	wire [4-1:0] node2395;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2401;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2408;
	wire [4-1:0] node2410;
	wire [4-1:0] node2413;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2416;
	wire [4-1:0] node2418;
	wire [4-1:0] node2421;
	wire [4-1:0] node2424;
	wire [4-1:0] node2426;
	wire [4-1:0] node2429;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2437;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2444;
	wire [4-1:0] node2447;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2453;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2466;
	wire [4-1:0] node2467;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2474;
	wire [4-1:0] node2475;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2487;
	wire [4-1:0] node2488;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2494;
	wire [4-1:0] node2495;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2506;
	wire [4-1:0] node2508;
	wire [4-1:0] node2510;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2517;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2537;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2544;
	wire [4-1:0] node2547;
	wire [4-1:0] node2549;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2568;
	wire [4-1:0] node2570;
	wire [4-1:0] node2573;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2578;
	wire [4-1:0] node2580;
	wire [4-1:0] node2582;
	wire [4-1:0] node2585;
	wire [4-1:0] node2586;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2593;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2601;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2614;
	wire [4-1:0] node2617;
	wire [4-1:0] node2618;
	wire [4-1:0] node2619;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2625;
	wire [4-1:0] node2627;
	wire [4-1:0] node2630;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2635;
	wire [4-1:0] node2636;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2644;
	wire [4-1:0] node2646;
	wire [4-1:0] node2649;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2657;
	wire [4-1:0] node2659;
	wire [4-1:0] node2661;
	wire [4-1:0] node2663;
	wire [4-1:0] node2665;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2673;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2685;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2691;
	wire [4-1:0] node2694;
	wire [4-1:0] node2695;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2706;
	wire [4-1:0] node2709;
	wire [4-1:0] node2710;
	wire [4-1:0] node2711;
	wire [4-1:0] node2716;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2728;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2734;
	wire [4-1:0] node2736;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2742;
	wire [4-1:0] node2744;
	wire [4-1:0] node2747;
	wire [4-1:0] node2748;
	wire [4-1:0] node2751;
	wire [4-1:0] node2752;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2763;
	wire [4-1:0] node2764;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2770;
	wire [4-1:0] node2771;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2784;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2789;
	wire [4-1:0] node2791;
	wire [4-1:0] node2794;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2801;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2808;
	wire [4-1:0] node2811;
	wire [4-1:0] node2813;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2820;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2828;
	wire [4-1:0] node2830;
	wire [4-1:0] node2832;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2838;
	wire [4-1:0] node2839;
	wire [4-1:0] node2840;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2847;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2855;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2861;
	wire [4-1:0] node2863;
	wire [4-1:0] node2865;
	wire [4-1:0] node2868;
	wire [4-1:0] node2869;
	wire [4-1:0] node2871;
	wire [4-1:0] node2874;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2880;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2886;
	wire [4-1:0] node2888;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2902;
	wire [4-1:0] node2905;
	wire [4-1:0] node2909;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2916;
	wire [4-1:0] node2917;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2930;
	wire [4-1:0] node2933;
	wire [4-1:0] node2936;
	wire [4-1:0] node2938;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2948;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2959;
	wire [4-1:0] node2960;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2980;
	wire [4-1:0] node2984;
	wire [4-1:0] node2985;
	wire [4-1:0] node2986;
	wire [4-1:0] node2987;
	wire [4-1:0] node2988;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2996;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3002;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3010;
	wire [4-1:0] node3011;
	wire [4-1:0] node3012;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3034;
	wire [4-1:0] node3037;
	wire [4-1:0] node3039;
	wire [4-1:0] node3040;
	wire [4-1:0] node3044;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3054;
	wire [4-1:0] node3055;
	wire [4-1:0] node3056;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3064;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3074;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3080;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3099;
	wire [4-1:0] node3101;
	wire [4-1:0] node3104;
	wire [4-1:0] node3106;
	wire [4-1:0] node3109;
	wire [4-1:0] node3110;
	wire [4-1:0] node3114;
	wire [4-1:0] node3115;
	wire [4-1:0] node3117;
	wire [4-1:0] node3118;
	wire [4-1:0] node3119;
	wire [4-1:0] node3123;
	wire [4-1:0] node3125;
	wire [4-1:0] node3127;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3146;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3152;
	wire [4-1:0] node3154;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3171;
	wire [4-1:0] node3173;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3179;
	wire [4-1:0] node3180;
	wire [4-1:0] node3182;
	wire [4-1:0] node3185;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3191;
	wire [4-1:0] node3192;
	wire [4-1:0] node3194;
	wire [4-1:0] node3196;
	wire [4-1:0] node3200;
	wire [4-1:0] node3202;
	wire [4-1:0] node3205;
	wire [4-1:0] node3206;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3214;
	wire [4-1:0] node3216;
	wire [4-1:0] node3218;
	wire [4-1:0] node3221;
	wire [4-1:0] node3224;
	wire [4-1:0] node3225;
	wire [4-1:0] node3226;
	wire [4-1:0] node3227;
	wire [4-1:0] node3231;
	wire [4-1:0] node3234;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3256;
	wire [4-1:0] node3257;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3281;
	wire [4-1:0] node3282;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3296;
	wire [4-1:0] node3297;
	wire [4-1:0] node3298;
	wire [4-1:0] node3300;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3305;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3313;
	wire [4-1:0] node3314;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3324;
	wire [4-1:0] node3325;
	wire [4-1:0] node3326;
	wire [4-1:0] node3331;
	wire [4-1:0] node3332;
	wire [4-1:0] node3333;
	wire [4-1:0] node3334;
	wire [4-1:0] node3336;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3343;
	wire [4-1:0] node3346;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3350;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3365;
	wire [4-1:0] node3366;
	wire [4-1:0] node3369;
	wire [4-1:0] node3372;
	wire [4-1:0] node3373;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3379;
	wire [4-1:0] node3381;
	wire [4-1:0] node3385;
	wire [4-1:0] node3386;
	wire [4-1:0] node3387;
	wire [4-1:0] node3388;
	wire [4-1:0] node3392;
	wire [4-1:0] node3395;
	wire [4-1:0] node3396;
	wire [4-1:0] node3399;
	wire [4-1:0] node3400;
	wire [4-1:0] node3402;
	wire [4-1:0] node3405;
	wire [4-1:0] node3407;
	wire [4-1:0] node3410;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3413;
	wire [4-1:0] node3414;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3418;
	wire [4-1:0] node3422;
	wire [4-1:0] node3425;
	wire [4-1:0] node3426;
	wire [4-1:0] node3428;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3436;
	wire [4-1:0] node3437;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3457;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3465;
	wire [4-1:0] node3466;
	wire [4-1:0] node3469;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3475;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3485;
	wire [4-1:0] node3487;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3492;
	wire [4-1:0] node3493;
	wire [4-1:0] node3494;
	wire [4-1:0] node3498;
	wire [4-1:0] node3500;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3505;
	wire [4-1:0] node3510;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3513;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3524;
	wire [4-1:0] node3530;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3536;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3545;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3552;
	wire [4-1:0] node3556;
	wire [4-1:0] node3557;
	wire [4-1:0] node3559;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3570;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3581;
	wire [4-1:0] node3582;
	wire [4-1:0] node3586;
	wire [4-1:0] node3587;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3595;
	wire [4-1:0] node3596;
	wire [4-1:0] node3597;
	wire [4-1:0] node3598;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3611;
	wire [4-1:0] node3613;
	wire [4-1:0] node3615;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3638;
	wire [4-1:0] node3640;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3646;
	wire [4-1:0] node3649;
	wire [4-1:0] node3651;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3659;
	wire [4-1:0] node3664;
	wire [4-1:0] node3666;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3672;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3677;
	wire [4-1:0] node3680;
	wire [4-1:0] node3683;
	wire [4-1:0] node3684;
	wire [4-1:0] node3687;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3702;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3716;
	wire [4-1:0] node3719;
	wire [4-1:0] node3721;
	wire [4-1:0] node3724;
	wire [4-1:0] node3726;
	wire [4-1:0] node3728;
	wire [4-1:0] node3729;
	wire [4-1:0] node3733;
	wire [4-1:0] node3734;
	wire [4-1:0] node3735;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3744;
	wire [4-1:0] node3745;
	wire [4-1:0] node3746;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3757;
	wire [4-1:0] node3758;
	wire [4-1:0] node3762;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3773;
	wire [4-1:0] node3775;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3784;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3791;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3797;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3808;
	wire [4-1:0] node3809;
	wire [4-1:0] node3814;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3826;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3833;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3837;
	wire [4-1:0] node3839;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3848;
	wire [4-1:0] node3849;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3854;
	wire [4-1:0] node3862;
	wire [4-1:0] node3863;
	wire [4-1:0] node3865;
	wire [4-1:0] node3867;
	wire [4-1:0] node3870;
	wire [4-1:0] node3871;
	wire [4-1:0] node3873;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3882;
	wire [4-1:0] node3886;
	wire [4-1:0] node3888;
	wire [4-1:0] node3891;
	wire [4-1:0] node3892;
	wire [4-1:0] node3894;
	wire [4-1:0] node3897;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3910;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3918;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3929;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3940;
	wire [4-1:0] node3944;
	wire [4-1:0] node3947;
	wire [4-1:0] node3950;
	wire [4-1:0] node3951;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3959;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3966;
	wire [4-1:0] node3970;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3978;
	wire [4-1:0] node3979;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3985;
	wire [4-1:0] node3987;
	wire [4-1:0] node3990;
	wire [4-1:0] node3992;
	wire [4-1:0] node3994;
	wire [4-1:0] node3997;
	wire [4-1:0] node3998;
	wire [4-1:0] node3999;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4006;
	wire [4-1:0] node4009;
	wire [4-1:0] node4012;
	wire [4-1:0] node4014;
	wire [4-1:0] node4017;
	wire [4-1:0] node4020;
	wire [4-1:0] node4021;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4037;
	wire [4-1:0] node4041;
	wire [4-1:0] node4043;
	wire [4-1:0] node4046;
	wire [4-1:0] node4048;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4060;
	wire [4-1:0] node4061;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4068;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4076;
	wire [4-1:0] node4077;
	wire [4-1:0] node4081;
	wire [4-1:0] node4082;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4090;
	wire [4-1:0] node4091;
	wire [4-1:0] node4093;
	wire [4-1:0] node4095;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4106;
	wire [4-1:0] node4108;
	wire [4-1:0] node4109;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4115;
	wire [4-1:0] node4117;
	wire [4-1:0] node4120;
	wire [4-1:0] node4123;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4129;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4136;
	wire [4-1:0] node4138;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4144;
	wire [4-1:0] node4150;
	wire [4-1:0] node4151;

	assign outp = (inp[6]) ? node2172 : node1;
		assign node1 = (inp[3]) ? node1129 : node2;
			assign node2 = (inp[14]) ? node538 : node3;
				assign node3 = (inp[8]) ? node275 : node4;
					assign node4 = (inp[11]) ? node142 : node5;
						assign node5 = (inp[12]) ? node71 : node6;
							assign node6 = (inp[7]) ? node42 : node7;
								assign node7 = (inp[5]) ? node27 : node8;
									assign node8 = (inp[9]) ? node18 : node9;
										assign node9 = (inp[0]) ? 4'b0110 : node10;
											assign node10 = (inp[2]) ? node14 : node11;
												assign node11 = (inp[13]) ? 4'b0011 : 4'b0001;
												assign node14 = (inp[4]) ? 4'b0001 : 4'b0000;
										assign node18 = (inp[2]) ? node20 : 4'b0100;
											assign node20 = (inp[1]) ? 4'b0010 : node21;
												assign node21 = (inp[15]) ? node23 : 4'b0001;
													assign node23 = (inp[13]) ? 4'b0000 : 4'b0100;
									assign node27 = (inp[2]) ? node35 : node28;
										assign node28 = (inp[1]) ? node32 : node29;
											assign node29 = (inp[15]) ? 4'b0001 : 4'b0101;
											assign node32 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node35 = (inp[15]) ? node37 : 4'b0101;
											assign node37 = (inp[0]) ? node39 : 4'b0101;
												assign node39 = (inp[10]) ? 4'b0111 : 4'b0011;
								assign node42 = (inp[15]) ? node54 : node43;
									assign node43 = (inp[13]) ? node49 : node44;
										assign node44 = (inp[0]) ? 4'b0010 : node45;
											assign node45 = (inp[2]) ? 4'b0111 : 4'b0011;
										assign node49 = (inp[9]) ? 4'b0110 : node50;
											assign node50 = (inp[4]) ? 4'b0010 : 4'b0110;
									assign node54 = (inp[4]) ? node58 : node55;
										assign node55 = (inp[5]) ? 4'b0110 : 4'b0010;
										assign node58 = (inp[0]) ? node62 : node59;
											assign node59 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node62 = (inp[2]) ? node68 : node63;
												assign node63 = (inp[1]) ? node65 : 4'b0000;
													assign node65 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node68 = (inp[9]) ? 4'b0101 : 4'b0100;
							assign node71 = (inp[7]) ? node109 : node72;
								assign node72 = (inp[15]) ? node94 : node73;
									assign node73 = (inp[5]) ? node79 : node74;
										assign node74 = (inp[1]) ? 4'b0010 : node75;
											assign node75 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node79 = (inp[13]) ? node85 : node80;
											assign node80 = (inp[4]) ? 4'b0010 : node81;
												assign node81 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node85 = (inp[10]) ? node89 : node86;
												assign node86 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node89 = (inp[4]) ? node91 : 4'b0010;
													assign node91 = (inp[0]) ? 4'b0110 : 4'b0111;
									assign node94 = (inp[4]) ? node102 : node95;
										assign node95 = (inp[10]) ? node99 : node96;
											assign node96 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node99 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node102 = (inp[5]) ? node104 : 4'b0001;
											assign node104 = (inp[9]) ? 4'b0000 : node105;
												assign node105 = (inp[2]) ? 4'b0101 : 4'b0000;
								assign node109 = (inp[4]) ? node123 : node110;
									assign node110 = (inp[1]) ? node112 : 4'b0000;
										assign node112 = (inp[13]) ? node118 : node113;
											assign node113 = (inp[2]) ? node115 : 4'b0001;
												assign node115 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node118 = (inp[2]) ? 4'b0001 : node119;
												assign node119 = (inp[10]) ? 4'b0101 : 4'b0100;
									assign node123 = (inp[15]) ? node131 : node124;
										assign node124 = (inp[1]) ? 4'b0000 : node125;
											assign node125 = (inp[13]) ? node127 : 4'b0100;
												assign node127 = (inp[0]) ? 4'b0001 : 4'b0100;
										assign node131 = (inp[5]) ? node135 : node132;
											assign node132 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node135 = (inp[9]) ? node137 : 4'b0010;
												assign node137 = (inp[13]) ? node139 : 4'b0010;
													assign node139 = (inp[1]) ? 4'b0011 : 4'b0111;
						assign node142 = (inp[7]) ? node196 : node143;
							assign node143 = (inp[12]) ? node167 : node144;
								assign node144 = (inp[4]) ? node154 : node145;
									assign node145 = (inp[9]) ? node149 : node146;
										assign node146 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node149 = (inp[15]) ? 4'b0001 : node150;
											assign node150 = (inp[10]) ? 4'b0001 : 4'b0000;
									assign node154 = (inp[15]) ? node160 : node155;
										assign node155 = (inp[2]) ? node157 : 4'b0100;
											assign node157 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node160 = (inp[0]) ? node164 : node161;
											assign node161 = (inp[5]) ? 4'b0011 : 4'b0110;
											assign node164 = (inp[10]) ? 4'b0111 : 4'b0110;
								assign node167 = (inp[15]) ? node179 : node168;
									assign node168 = (inp[0]) ? node174 : node169;
										assign node169 = (inp[2]) ? node171 : 4'b0111;
											assign node171 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node174 = (inp[1]) ? 4'b0011 : node175;
											assign node175 = (inp[5]) ? 4'b0010 : 4'b0110;
									assign node179 = (inp[4]) ? node189 : node180;
										assign node180 = (inp[1]) ? node186 : node181;
											assign node181 = (inp[13]) ? 4'b0011 : node182;
												assign node182 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node186 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node189 = (inp[13]) ? node193 : node190;
											assign node190 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node193 = (inp[9]) ? 4'b0001 : 4'b0000;
							assign node196 = (inp[15]) ? node222 : node197;
								assign node197 = (inp[12]) ? node207 : node198;
									assign node198 = (inp[1]) ? node200 : 4'b0011;
										assign node200 = (inp[10]) ? node204 : node201;
											assign node201 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node204 = (inp[9]) ? 4'b0010 : 4'b0011;
									assign node207 = (inp[4]) ? node217 : node208;
										assign node208 = (inp[1]) ? node212 : node209;
											assign node209 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node212 = (inp[9]) ? 4'b0101 : node213;
												assign node213 = (inp[2]) ? 4'b0000 : 4'b0100;
										assign node217 = (inp[0]) ? node219 : 4'b0001;
											assign node219 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node222 = (inp[0]) ? node250 : node223;
									assign node223 = (inp[4]) ? node237 : node224;
										assign node224 = (inp[12]) ? node234 : node225;
											assign node225 = (inp[1]) ? node227 : 4'b0110;
												assign node227 = (inp[9]) ? 4'b0110 : node228;
													assign node228 = (inp[5]) ? node230 : 4'b0010;
														assign node230 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node234 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node237 = (inp[12]) ? node239 : 4'b0101;
											assign node239 = (inp[5]) ? node247 : node240;
												assign node240 = (inp[1]) ? node242 : 4'b0110;
													assign node242 = (inp[13]) ? node244 : 4'b0111;
														assign node244 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node247 = (inp[13]) ? 4'b0110 : 4'b0010;
									assign node250 = (inp[2]) ? node264 : node251;
										assign node251 = (inp[9]) ? node255 : node252;
											assign node252 = (inp[12]) ? 4'b0110 : 4'b0100;
											assign node255 = (inp[10]) ? node259 : node256;
												assign node256 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node259 = (inp[4]) ? 4'b0111 : node260;
													assign node260 = (inp[12]) ? 4'b0001 : 4'b0011;
										assign node264 = (inp[13]) ? node268 : node265;
											assign node265 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node268 = (inp[4]) ? node272 : node269;
												assign node269 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node272 = (inp[12]) ? 4'b0011 : 4'b0001;
					assign node275 = (inp[1]) ? node409 : node276;
						assign node276 = (inp[2]) ? node338 : node277;
							assign node277 = (inp[10]) ? node311 : node278;
								assign node278 = (inp[4]) ? node292 : node279;
									assign node279 = (inp[12]) ? node283 : node280;
										assign node280 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node283 = (inp[13]) ? node287 : node284;
											assign node284 = (inp[15]) ? 4'b1011 : 4'b1010;
											assign node287 = (inp[15]) ? node289 : 4'b1011;
												assign node289 = (inp[5]) ? 4'b1011 : 4'b1110;
									assign node292 = (inp[12]) ? 4'b1001 : node293;
										assign node293 = (inp[9]) ? node301 : node294;
											assign node294 = (inp[5]) ? node296 : 4'b1011;
												assign node296 = (inp[11]) ? node298 : 4'b1111;
													assign node298 = (inp[15]) ? 4'b1111 : 4'b1011;
											assign node301 = (inp[7]) ? node307 : node302;
												assign node302 = (inp[15]) ? 4'b1010 : node303;
													assign node303 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node307 = (inp[0]) ? 4'b1011 : 4'b1010;
								assign node311 = (inp[13]) ? node327 : node312;
									assign node312 = (inp[5]) ? node322 : node313;
										assign node313 = (inp[0]) ? node317 : node314;
											assign node314 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node317 = (inp[4]) ? 4'b1100 : node318;
												assign node318 = (inp[12]) ? 4'b1010 : 4'b1100;
										assign node322 = (inp[7]) ? 4'b1000 : node323;
											assign node323 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node327 = (inp[15]) ? 4'b1010 : node328;
										assign node328 = (inp[5]) ? node334 : node329;
											assign node329 = (inp[9]) ? node331 : 4'b1000;
												assign node331 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node334 = (inp[12]) ? 4'b1111 : 4'b1100;
							assign node338 = (inp[7]) ? node376 : node339;
								assign node339 = (inp[12]) ? node357 : node340;
									assign node340 = (inp[4]) ? node348 : node341;
										assign node341 = (inp[10]) ? node343 : 4'b1101;
											assign node343 = (inp[11]) ? 4'b1100 : node344;
												assign node344 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node348 = (inp[5]) ? node354 : node349;
											assign node349 = (inp[13]) ? 4'b1111 : node350;
												assign node350 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node354 = (inp[15]) ? 4'b1011 : 4'b1111;
									assign node357 = (inp[4]) ? node359 : 4'b1111;
										assign node359 = (inp[5]) ? node365 : node360;
											assign node360 = (inp[10]) ? node362 : 4'b1000;
												assign node362 = (inp[15]) ? 4'b1101 : 4'b1001;
											assign node365 = (inp[13]) ? node367 : 4'b1101;
												assign node367 = (inp[9]) ? 4'b1100 : node368;
													assign node368 = (inp[0]) ? 4'b1101 : node369;
														assign node369 = (inp[10]) ? 4'b1100 : node370;
															assign node370 = (inp[15]) ? 4'b1100 : 4'b1101;
								assign node376 = (inp[0]) ? node390 : node377;
									assign node377 = (inp[10]) ? node383 : node378;
										assign node378 = (inp[4]) ? node380 : 4'b1010;
											assign node380 = (inp[15]) ? 4'b1000 : 4'b1100;
										assign node383 = (inp[4]) ? node387 : node384;
											assign node384 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node387 = (inp[5]) ? 4'b1101 : 4'b1110;
									assign node390 = (inp[15]) ? node400 : node391;
										assign node391 = (inp[5]) ? node395 : node392;
											assign node392 = (inp[10]) ? 4'b1111 : 4'b1100;
											assign node395 = (inp[10]) ? node397 : 4'b1011;
												assign node397 = (inp[4]) ? 4'b1011 : 4'b1000;
										assign node400 = (inp[9]) ? node406 : node401;
											assign node401 = (inp[5]) ? node403 : 4'b1110;
												assign node403 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node406 = (inp[5]) ? 4'b1100 : 4'b1010;
						assign node409 = (inp[2]) ? node461 : node410;
							assign node410 = (inp[7]) ? node438 : node411;
								assign node411 = (inp[13]) ? node425 : node412;
									assign node412 = (inp[4]) ? node418 : node413;
										assign node413 = (inp[12]) ? 4'b1111 : node414;
											assign node414 = (inp[5]) ? 4'b1101 : 4'b1100;
										assign node418 = (inp[12]) ? 4'b1101 : node419;
											assign node419 = (inp[15]) ? node421 : 4'b1111;
												assign node421 = (inp[9]) ? 4'b1010 : 4'b1110;
									assign node425 = (inp[11]) ? node433 : node426;
										assign node426 = (inp[12]) ? node430 : node427;
											assign node427 = (inp[4]) ? 4'b1110 : 4'b1100;
											assign node430 = (inp[5]) ? 4'b1100 : 4'b1001;
										assign node433 = (inp[12]) ? 4'b1110 : node434;
											assign node434 = (inp[4]) ? 4'b1110 : 4'b1100;
								assign node438 = (inp[4]) ? node452 : node439;
									assign node439 = (inp[12]) ? node443 : node440;
										assign node440 = (inp[13]) ? 4'b1101 : 4'b1000;
										assign node443 = (inp[5]) ? node447 : node444;
											assign node444 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node447 = (inp[15]) ? node449 : 4'b1011;
												assign node449 = (inp[13]) ? 4'b1110 : 4'b1111;
									assign node452 = (inp[12]) ? node456 : node453;
										assign node453 = (inp[11]) ? 4'b1111 : 4'b1010;
										assign node456 = (inp[9]) ? 4'b1100 : node457;
											assign node457 = (inp[0]) ? 4'b1101 : 4'b1100;
							assign node461 = (inp[7]) ? node499 : node462;
								assign node462 = (inp[5]) ? node480 : node463;
									assign node463 = (inp[9]) ? node471 : node464;
										assign node464 = (inp[12]) ? 4'b1010 : node465;
											assign node465 = (inp[13]) ? 4'b1001 : node466;
												assign node466 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node471 = (inp[15]) ? node477 : node472;
											assign node472 = (inp[12]) ? node474 : 4'b1000;
												assign node474 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node477 = (inp[13]) ? 4'b1010 : 4'b1000;
									assign node480 = (inp[15]) ? node488 : node481;
										assign node481 = (inp[12]) ? node485 : node482;
											assign node482 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node485 = (inp[4]) ? 4'b1001 : 4'b1011;
										assign node488 = (inp[12]) ? node490 : 4'b1000;
											assign node490 = (inp[4]) ? node492 : 4'b1011;
												assign node492 = (inp[10]) ? node494 : 4'b1000;
													assign node494 = (inp[11]) ? 4'b1001 : node495;
														assign node495 = (inp[9]) ? 4'b1000 : 4'b1001;
								assign node499 = (inp[5]) ? node519 : node500;
									assign node500 = (inp[15]) ? node508 : node501;
										assign node501 = (inp[13]) ? node505 : node502;
											assign node502 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node505 = (inp[4]) ? 4'b1001 : 4'b1011;
										assign node508 = (inp[12]) ? node514 : node509;
											assign node509 = (inp[4]) ? node511 : 4'b1101;
												assign node511 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node514 = (inp[0]) ? 4'b1101 : node515;
												assign node515 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node519 = (inp[15]) ? node531 : node520;
										assign node520 = (inp[11]) ? node528 : node521;
											assign node521 = (inp[9]) ? 4'b1000 : node522;
												assign node522 = (inp[12]) ? 4'b1110 : node523;
													assign node523 = (inp[13]) ? 4'b1100 : 4'b1110;
											assign node528 = (inp[4]) ? 4'b1111 : 4'b1101;
										assign node531 = (inp[11]) ? 4'b1010 : node532;
											assign node532 = (inp[4]) ? 4'b1001 : node533;
												assign node533 = (inp[12]) ? 4'b1010 : 4'b1000;
				assign node538 = (inp[12]) ? node804 : node539;
					assign node539 = (inp[4]) ? node689 : node540;
						assign node540 = (inp[8]) ? node620 : node541;
							assign node541 = (inp[7]) ? node579 : node542;
								assign node542 = (inp[15]) ? node564 : node543;
									assign node543 = (inp[2]) ? node549 : node544;
										assign node544 = (inp[5]) ? 4'b1000 : node545;
											assign node545 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node549 = (inp[10]) ? node555 : node550;
											assign node550 = (inp[5]) ? node552 : 4'b1000;
												assign node552 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node555 = (inp[13]) ? node559 : node556;
												assign node556 = (inp[11]) ? 4'b1000 : 4'b1100;
												assign node559 = (inp[11]) ? 4'b1001 : node560;
													assign node560 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node564 = (inp[10]) ? node574 : node565;
										assign node565 = (inp[2]) ? node569 : node566;
											assign node566 = (inp[5]) ? 4'b1010 : 4'b1111;
											assign node569 = (inp[1]) ? 4'b1010 : node570;
												assign node570 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node574 = (inp[0]) ? node576 : 4'b1011;
											assign node576 = (inp[11]) ? 4'b1111 : 4'b1110;
								assign node579 = (inp[15]) ? node605 : node580;
									assign node580 = (inp[10]) ? node588 : node581;
										assign node581 = (inp[9]) ? 4'b1110 : node582;
											assign node582 = (inp[13]) ? node584 : 4'b1111;
												assign node584 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node588 = (inp[2]) ? node596 : node589;
											assign node589 = (inp[11]) ? 4'b1011 : node590;
												assign node590 = (inp[5]) ? 4'b1111 : node591;
													assign node591 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node596 = (inp[0]) ? 4'b1011 : node597;
												assign node597 = (inp[1]) ? 4'b1010 : node598;
													assign node598 = (inp[5]) ? node600 : 4'b1010;
														assign node600 = (inp[13]) ? 4'b1111 : 4'b1010;
									assign node605 = (inp[10]) ? node613 : node606;
										assign node606 = (inp[9]) ? 4'b1101 : node607;
											assign node607 = (inp[0]) ? 4'b1001 : node608;
												assign node608 = (inp[1]) ? 4'b1001 : 4'b1101;
										assign node613 = (inp[5]) ? node617 : node614;
											assign node614 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node617 = (inp[1]) ? 4'b1101 : 4'b1001;
							assign node620 = (inp[2]) ? node664 : node621;
								assign node621 = (inp[1]) ? node643 : node622;
									assign node622 = (inp[9]) ? node636 : node623;
										assign node623 = (inp[7]) ? node631 : node624;
											assign node624 = (inp[0]) ? node626 : 4'b1000;
												assign node626 = (inp[15]) ? 4'b1001 : node627;
													assign node627 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node631 = (inp[0]) ? node633 : 4'b1001;
												assign node633 = (inp[10]) ? 4'b1000 : 4'b1001;
										assign node636 = (inp[15]) ? 4'b1101 : node637;
											assign node637 = (inp[13]) ? node639 : 4'b1101;
												assign node639 = (inp[7]) ? 4'b1000 : 4'b1100;
									assign node643 = (inp[5]) ? node655 : node644;
										assign node644 = (inp[13]) ? 4'b1101 : node645;
											assign node645 = (inp[11]) ? node651 : node646;
												assign node646 = (inp[0]) ? node648 : 4'b1101;
													assign node648 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node651 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node655 = (inp[11]) ? node657 : 4'b1101;
											assign node657 = (inp[10]) ? node659 : 4'b1100;
												assign node659 = (inp[13]) ? node661 : 4'b1000;
													assign node661 = (inp[15]) ? 4'b1000 : 4'b1100;
								assign node664 = (inp[9]) ? node682 : node665;
									assign node665 = (inp[13]) ? node673 : node666;
										assign node666 = (inp[0]) ? 4'b1100 : node667;
											assign node667 = (inp[5]) ? node669 : 4'b1101;
												assign node669 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node673 = (inp[1]) ? 4'b1000 : node674;
											assign node674 = (inp[5]) ? 4'b1001 : node675;
												assign node675 = (inp[11]) ? 4'b1100 : node676;
													assign node676 = (inp[15]) ? 4'b1100 : 4'b1101;
									assign node682 = (inp[5]) ? node684 : 4'b1001;
										assign node684 = (inp[1]) ? 4'b1100 : node685;
											assign node685 = (inp[15]) ? 4'b1100 : 4'b1000;
						assign node689 = (inp[7]) ? node759 : node690;
							assign node690 = (inp[8]) ? node730 : node691;
								assign node691 = (inp[13]) ? node711 : node692;
									assign node692 = (inp[5]) ? node702 : node693;
										assign node693 = (inp[0]) ? node695 : 4'b1101;
											assign node695 = (inp[9]) ? node697 : 4'b1001;
												assign node697 = (inp[10]) ? 4'b1100 : node698;
													assign node698 = (inp[1]) ? 4'b1001 : 4'b1101;
										assign node702 = (inp[11]) ? node704 : 4'b1000;
											assign node704 = (inp[0]) ? 4'b1100 : node705;
												assign node705 = (inp[2]) ? 4'b1100 : node706;
													assign node706 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node711 = (inp[0]) ? node717 : node712;
										assign node712 = (inp[15]) ? node714 : 4'b1000;
											assign node714 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node717 = (inp[10]) ? node727 : node718;
											assign node718 = (inp[2]) ? node720 : 4'b1100;
												assign node720 = (inp[9]) ? 4'b1100 : node721;
													assign node721 = (inp[11]) ? 4'b1000 : node722;
														assign node722 = (inp[15]) ? 4'b1100 : 4'b1000;
											assign node727 = (inp[1]) ? 4'b1000 : 4'b1001;
								assign node730 = (inp[11]) ? node740 : node731;
									assign node731 = (inp[13]) ? 4'b1110 : node732;
										assign node732 = (inp[15]) ? 4'b1111 : node733;
											assign node733 = (inp[2]) ? node735 : 4'b1111;
												assign node735 = (inp[10]) ? 4'b1110 : 4'b1010;
									assign node740 = (inp[10]) ? node752 : node741;
										assign node741 = (inp[9]) ? node747 : node742;
											assign node742 = (inp[2]) ? 4'b1011 : node743;
												assign node743 = (inp[5]) ? 4'b1011 : 4'b1110;
											assign node747 = (inp[13]) ? node749 : 4'b1111;
												assign node749 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node752 = (inp[0]) ? 4'b1110 : node753;
											assign node753 = (inp[2]) ? 4'b1110 : node754;
												assign node754 = (inp[1]) ? 4'b1011 : 4'b1010;
							assign node759 = (inp[2]) ? node775 : node760;
								assign node760 = (inp[13]) ? node770 : node761;
									assign node761 = (inp[11]) ? node763 : 4'b1010;
										assign node763 = (inp[10]) ? node765 : 4'b1110;
											assign node765 = (inp[8]) ? node767 : 4'b1010;
												assign node767 = (inp[1]) ? 4'b1110 : 4'b1010;
									assign node770 = (inp[8]) ? 4'b1010 : node771;
										assign node771 = (inp[0]) ? 4'b1111 : 4'b1110;
								assign node775 = (inp[1]) ? node787 : node776;
									assign node776 = (inp[8]) ? 4'b1111 : node777;
										assign node777 = (inp[0]) ? node783 : node778;
											assign node778 = (inp[10]) ? 4'b1010 : node779;
												assign node779 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node783 = (inp[5]) ? 4'b1110 : 4'b1111;
									assign node787 = (inp[9]) ? node797 : node788;
										assign node788 = (inp[15]) ? node790 : 4'b1010;
											assign node790 = (inp[10]) ? node792 : 4'b1011;
												assign node792 = (inp[5]) ? node794 : 4'b1010;
													assign node794 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node797 = (inp[8]) ? 4'b1011 : node798;
											assign node798 = (inp[5]) ? 4'b1011 : node799;
												assign node799 = (inp[10]) ? 4'b1111 : 4'b1110;
					assign node804 = (inp[4]) ? node996 : node805;
						assign node805 = (inp[8]) ? node921 : node806;
							assign node806 = (inp[0]) ? node866 : node807;
								assign node807 = (inp[5]) ? node835 : node808;
									assign node808 = (inp[7]) ? node826 : node809;
										assign node809 = (inp[15]) ? 4'b1101 : node810;
											assign node810 = (inp[10]) ? node818 : node811;
												assign node811 = (inp[11]) ? node813 : 4'b1010;
													assign node813 = (inp[9]) ? node815 : 4'b1110;
														assign node815 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node818 = (inp[9]) ? node820 : 4'b1111;
													assign node820 = (inp[13]) ? node822 : 4'b1010;
														assign node822 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node826 = (inp[15]) ? 4'b1010 : node827;
											assign node827 = (inp[2]) ? node829 : 4'b1000;
												assign node829 = (inp[13]) ? 4'b1101 : node830;
													assign node830 = (inp[10]) ? 4'b1000 : 4'b1001;
									assign node835 = (inp[11]) ? node851 : node836;
										assign node836 = (inp[10]) ? node844 : node837;
											assign node837 = (inp[15]) ? 4'b1110 : node838;
												assign node838 = (inp[2]) ? node840 : 4'b1001;
													assign node840 = (inp[13]) ? 4'b1001 : 4'b1100;
											assign node844 = (inp[2]) ? 4'b1111 : node845;
												assign node845 = (inp[7]) ? 4'b1111 : node846;
													assign node846 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node851 = (inp[2]) ? node857 : node852;
											assign node852 = (inp[1]) ? node854 : 4'b1111;
												assign node854 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node857 = (inp[7]) ? node863 : node858;
												assign node858 = (inp[10]) ? 4'b1000 : node859;
													assign node859 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node863 = (inp[1]) ? 4'b1100 : 4'b1001;
								assign node866 = (inp[10]) ? node882 : node867;
									assign node867 = (inp[1]) ? node875 : node868;
										assign node868 = (inp[5]) ? node872 : node869;
											assign node869 = (inp[2]) ? 4'b1001 : 4'b1010;
											assign node872 = (inp[2]) ? 4'b1010 : 4'b1110;
										assign node875 = (inp[15]) ? 4'b1100 : node876;
											assign node876 = (inp[9]) ? node878 : 4'b1110;
												assign node878 = (inp[2]) ? 4'b1111 : 4'b1010;
									assign node882 = (inp[9]) ? node908 : node883;
										assign node883 = (inp[11]) ? node901 : node884;
											assign node884 = (inp[7]) ? node890 : node885;
												assign node885 = (inp[5]) ? node887 : 4'b1101;
													assign node887 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node890 = (inp[13]) ? 4'b1101 : node891;
													assign node891 = (inp[2]) ? node897 : node892;
														assign node892 = (inp[5]) ? 4'b1001 : node893;
															assign node893 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node897 = (inp[5]) ? 4'b1100 : 4'b1000;
											assign node901 = (inp[5]) ? node905 : node902;
												assign node902 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node905 = (inp[1]) ? 4'b1011 : 4'b1010;
										assign node908 = (inp[13]) ? node916 : node909;
											assign node909 = (inp[1]) ? node911 : 4'b1110;
												assign node911 = (inp[5]) ? 4'b1010 : node912;
													assign node912 = (inp[15]) ? 4'b1111 : 4'b1010;
											assign node916 = (inp[1]) ? 4'b1100 : node917;
												assign node917 = (inp[15]) ? 4'b1110 : 4'b1100;
							assign node921 = (inp[13]) ? node961 : node922;
								assign node922 = (inp[10]) ? node938 : node923;
									assign node923 = (inp[15]) ? node931 : node924;
										assign node924 = (inp[7]) ? 4'b1010 : node925;
											assign node925 = (inp[11]) ? node927 : 4'b1010;
												assign node927 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node931 = (inp[2]) ? 4'b1011 : node932;
											assign node932 = (inp[5]) ? 4'b1010 : node933;
												assign node933 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node938 = (inp[1]) ? node950 : node939;
										assign node939 = (inp[2]) ? 4'b1111 : node940;
											assign node940 = (inp[7]) ? node944 : node941;
												assign node941 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node944 = (inp[15]) ? 4'b1010 : node945;
													assign node945 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node950 = (inp[11]) ? node956 : node951;
											assign node951 = (inp[15]) ? node953 : 4'b1010;
												assign node953 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node956 = (inp[5]) ? 4'b1111 : node957;
												assign node957 = (inp[0]) ? 4'b1110 : 4'b1010;
								assign node961 = (inp[11]) ? node975 : node962;
									assign node962 = (inp[1]) ? node966 : node963;
										assign node963 = (inp[2]) ? 4'b1111 : 4'b1011;
										assign node966 = (inp[2]) ? node972 : node967;
											assign node967 = (inp[0]) ? node969 : 4'b1111;
												assign node969 = (inp[15]) ? 4'b1010 : 4'b1110;
											assign node972 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node975 = (inp[15]) ? node981 : node976;
										assign node976 = (inp[1]) ? node978 : 4'b1010;
											assign node978 = (inp[2]) ? 4'b1010 : 4'b1110;
										assign node981 = (inp[2]) ? node985 : node982;
											assign node982 = (inp[5]) ? 4'b1111 : 4'b1010;
											assign node985 = (inp[7]) ? 4'b1110 : node986;
												assign node986 = (inp[0]) ? 4'b1010 : node987;
													assign node987 = (inp[10]) ? 4'b1110 : node988;
														assign node988 = (inp[5]) ? node990 : 4'b1010;
															assign node990 = (inp[1]) ? 4'b1010 : 4'b1110;
						assign node996 = (inp[7]) ? node1066 : node997;
							assign node997 = (inp[8]) ? node1035 : node998;
								assign node998 = (inp[1]) ? node1018 : node999;
									assign node999 = (inp[9]) ? node1009 : node1000;
										assign node1000 = (inp[11]) ? node1004 : node1001;
											assign node1001 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node1004 = (inp[0]) ? node1006 : 4'b1011;
												assign node1006 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node1009 = (inp[10]) ? node1013 : node1010;
											assign node1010 = (inp[15]) ? 4'b1110 : 4'b1010;
											assign node1013 = (inp[13]) ? 4'b1111 : node1014;
												assign node1014 = (inp[5]) ? 4'b1010 : 4'b1011;
									assign node1018 = (inp[5]) ? node1024 : node1019;
										assign node1019 = (inp[11]) ? 4'b1110 : node1020;
											assign node1020 = (inp[9]) ? 4'b1110 : 4'b1010;
										assign node1024 = (inp[9]) ? node1032 : node1025;
											assign node1025 = (inp[2]) ? node1027 : 4'b1110;
												assign node1027 = (inp[11]) ? node1029 : 4'b1010;
													assign node1029 = (inp[0]) ? 4'b1010 : 4'b1111;
											assign node1032 = (inp[11]) ? 4'b1010 : 4'b1011;
								assign node1035 = (inp[13]) ? node1057 : node1036;
									assign node1036 = (inp[11]) ? node1048 : node1037;
										assign node1037 = (inp[15]) ? node1041 : node1038;
											assign node1038 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node1041 = (inp[9]) ? node1043 : 4'b1001;
												assign node1043 = (inp[10]) ? 4'b1000 : node1044;
													assign node1044 = (inp[5]) ? 4'b1000 : 4'b1001;
										assign node1048 = (inp[9]) ? node1050 : 4'b1000;
											assign node1050 = (inp[0]) ? node1052 : 4'b1001;
												assign node1052 = (inp[15]) ? node1054 : 4'b1101;
													assign node1054 = (inp[2]) ? 4'b1101 : 4'b1001;
									assign node1057 = (inp[0]) ? node1059 : 4'b1101;
										assign node1059 = (inp[1]) ? 4'b1100 : node1060;
											assign node1060 = (inp[11]) ? 4'b1001 : node1061;
												assign node1061 = (inp[2]) ? 4'b1100 : 4'b1101;
							assign node1066 = (inp[1]) ? node1094 : node1067;
								assign node1067 = (inp[10]) ? node1081 : node1068;
									assign node1068 = (inp[15]) ? node1076 : node1069;
										assign node1069 = (inp[2]) ? node1073 : node1070;
											assign node1070 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node1073 = (inp[5]) ? 4'b1000 : 4'b1100;
										assign node1076 = (inp[0]) ? node1078 : 4'b1001;
											assign node1078 = (inp[9]) ? 4'b1000 : 4'b1001;
									assign node1081 = (inp[8]) ? node1091 : node1082;
										assign node1082 = (inp[13]) ? node1084 : 4'b1101;
											assign node1084 = (inp[11]) ? node1086 : 4'b1000;
												assign node1086 = (inp[9]) ? node1088 : 4'b1101;
													assign node1088 = (inp[15]) ? 4'b1000 : 4'b1100;
										assign node1091 = (inp[2]) ? 4'b1100 : 4'b1000;
								assign node1094 = (inp[0]) ? node1120 : node1095;
									assign node1095 = (inp[15]) ? node1113 : node1096;
										assign node1096 = (inp[8]) ? node1106 : node1097;
											assign node1097 = (inp[13]) ? node1103 : node1098;
												assign node1098 = (inp[10]) ? 4'b1101 : node1099;
													assign node1099 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node1103 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node1106 = (inp[2]) ? node1108 : 4'b1101;
												assign node1108 = (inp[11]) ? 4'b1001 : node1109;
													assign node1109 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node1113 = (inp[13]) ? node1117 : node1114;
											assign node1114 = (inp[5]) ? 4'b1000 : 4'b1100;
											assign node1117 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node1120 = (inp[5]) ? 4'b1001 : node1121;
										assign node1121 = (inp[13]) ? 4'b1000 : node1122;
											assign node1122 = (inp[10]) ? node1124 : 4'b1001;
												assign node1124 = (inp[15]) ? 4'b1000 : 4'b1001;
			assign node1129 = (inp[8]) ? node1715 : node1130;
				assign node1130 = (inp[14]) ? node1420 : node1131;
					assign node1131 = (inp[2]) ? node1245 : node1132;
						assign node1132 = (inp[13]) ? node1194 : node1133;
							assign node1133 = (inp[11]) ? node1159 : node1134;
								assign node1134 = (inp[4]) ? node1146 : node1135;
									assign node1135 = (inp[10]) ? node1139 : node1136;
										assign node1136 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node1139 = (inp[15]) ? 4'b1011 : node1140;
											assign node1140 = (inp[0]) ? 4'b1010 : node1141;
												assign node1141 = (inp[12]) ? 4'b1111 : 4'b1010;
									assign node1146 = (inp[1]) ? node1150 : node1147;
										assign node1147 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node1150 = (inp[9]) ? 4'b1111 : node1151;
											assign node1151 = (inp[0]) ? node1153 : 4'b1110;
												assign node1153 = (inp[12]) ? 4'b1010 : node1154;
													assign node1154 = (inp[7]) ? 4'b1011 : 4'b1101;
								assign node1159 = (inp[5]) ? node1183 : node1160;
									assign node1160 = (inp[1]) ? node1174 : node1161;
										assign node1161 = (inp[4]) ? node1165 : node1162;
											assign node1162 = (inp[9]) ? 4'b1010 : 4'b1000;
											assign node1165 = (inp[12]) ? node1171 : node1166;
												assign node1166 = (inp[15]) ? 4'b1100 : node1167;
													assign node1167 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node1171 = (inp[9]) ? 4'b1100 : 4'b1010;
										assign node1174 = (inp[10]) ? node1176 : 4'b1001;
											assign node1176 = (inp[4]) ? node1180 : node1177;
												assign node1177 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node1180 = (inp[15]) ? 4'b1001 : 4'b1101;
									assign node1183 = (inp[15]) ? node1191 : node1184;
										assign node1184 = (inp[9]) ? 4'b1101 : node1185;
											assign node1185 = (inp[10]) ? node1187 : 4'b1111;
												assign node1187 = (inp[1]) ? 4'b1010 : 4'b1100;
										assign node1191 = (inp[0]) ? 4'b1011 : 4'b1001;
							assign node1194 = (inp[4]) ? node1218 : node1195;
								assign node1195 = (inp[1]) ? node1211 : node1196;
									assign node1196 = (inp[9]) ? node1198 : 4'b1001;
										assign node1198 = (inp[7]) ? node1206 : node1199;
											assign node1199 = (inp[0]) ? 4'b1101 : node1200;
												assign node1200 = (inp[11]) ? node1202 : 4'b1100;
													assign node1202 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node1206 = (inp[15]) ? 4'b1100 : node1207;
												assign node1207 = (inp[10]) ? 4'b1111 : 4'b1110;
									assign node1211 = (inp[12]) ? node1213 : 4'b1000;
										assign node1213 = (inp[7]) ? node1215 : 4'b1110;
											assign node1215 = (inp[15]) ? 4'b1101 : 4'b1100;
								assign node1218 = (inp[15]) ? node1236 : node1219;
									assign node1219 = (inp[5]) ? node1227 : node1220;
										assign node1220 = (inp[11]) ? 4'b1110 : node1221;
											assign node1221 = (inp[7]) ? node1223 : 4'b1110;
												assign node1223 = (inp[12]) ? 4'b1111 : 4'b1001;
										assign node1227 = (inp[0]) ? node1231 : node1228;
											assign node1228 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node1231 = (inp[1]) ? 4'b1001 : node1232;
												assign node1232 = (inp[12]) ? 4'b1111 : 4'b1001;
									assign node1236 = (inp[1]) ? node1240 : node1237;
										assign node1237 = (inp[7]) ? 4'b1101 : 4'b1110;
										assign node1240 = (inp[7]) ? 4'b1110 : node1241;
											assign node1241 = (inp[11]) ? 4'b1111 : 4'b1011;
						assign node1245 = (inp[13]) ? node1329 : node1246;
							assign node1246 = (inp[1]) ? node1280 : node1247;
								assign node1247 = (inp[9]) ? node1265 : node1248;
									assign node1248 = (inp[5]) ? node1254 : node1249;
										assign node1249 = (inp[4]) ? node1251 : 4'b1111;
											assign node1251 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node1254 = (inp[0]) ? node1256 : 4'b1111;
											assign node1256 = (inp[15]) ? node1262 : node1257;
												assign node1257 = (inp[12]) ? 4'b1001 : node1258;
													assign node1258 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node1262 = (inp[4]) ? 4'b1011 : 4'b1111;
									assign node1265 = (inp[11]) ? node1277 : node1266;
										assign node1266 = (inp[12]) ? node1274 : node1267;
											assign node1267 = (inp[7]) ? node1271 : node1268;
												assign node1268 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node1271 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node1274 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node1277 = (inp[7]) ? 4'b1101 : 4'b1111;
								assign node1280 = (inp[5]) ? node1306 : node1281;
									assign node1281 = (inp[7]) ? node1291 : node1282;
										assign node1282 = (inp[12]) ? node1286 : node1283;
											assign node1283 = (inp[15]) ? 4'b1000 : 4'b1001;
											assign node1286 = (inp[9]) ? 4'b1010 : node1287;
												assign node1287 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node1291 = (inp[0]) ? node1301 : node1292;
											assign node1292 = (inp[9]) ? 4'b1001 : node1293;
												assign node1293 = (inp[10]) ? 4'b1101 : node1294;
													assign node1294 = (inp[12]) ? 4'b1011 : node1295;
														assign node1295 = (inp[11]) ? 4'b1111 : 4'b1101;
											assign node1301 = (inp[9]) ? 4'b1111 : node1302;
												assign node1302 = (inp[15]) ? 4'b1010 : 4'b1110;
									assign node1306 = (inp[0]) ? node1320 : node1307;
										assign node1307 = (inp[4]) ? node1309 : 4'b1110;
											assign node1309 = (inp[11]) ? node1315 : node1310;
												assign node1310 = (inp[15]) ? node1312 : 4'b1111;
													assign node1312 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node1315 = (inp[10]) ? node1317 : 4'b1000;
													assign node1317 = (inp[12]) ? 4'b1100 : 4'b1111;
										assign node1320 = (inp[11]) ? node1324 : node1321;
											assign node1321 = (inp[15]) ? 4'b1100 : 4'b1000;
											assign node1324 = (inp[7]) ? 4'b1110 : node1325;
												assign node1325 = (inp[12]) ? 4'b1110 : 4'b1101;
							assign node1329 = (inp[5]) ? node1373 : node1330;
								assign node1330 = (inp[1]) ? node1350 : node1331;
									assign node1331 = (inp[7]) ? node1343 : node1332;
										assign node1332 = (inp[15]) ? node1336 : node1333;
											assign node1333 = (inp[10]) ? 4'b1011 : 4'b1101;
											assign node1336 = (inp[4]) ? node1338 : 4'b1011;
												assign node1338 = (inp[10]) ? node1340 : 4'b1010;
													assign node1340 = (inp[9]) ? 4'b1011 : 4'b1010;
										assign node1343 = (inp[15]) ? node1345 : 4'b1010;
											assign node1345 = (inp[12]) ? 4'b1000 : node1346;
												assign node1346 = (inp[11]) ? 4'b1011 : 4'b1110;
									assign node1350 = (inp[9]) ? node1364 : node1351;
										assign node1351 = (inp[10]) ? node1357 : node1352;
											assign node1352 = (inp[15]) ? 4'b1100 : node1353;
												assign node1353 = (inp[7]) ? 4'b1010 : 4'b1110;
											assign node1357 = (inp[11]) ? node1359 : 4'b1110;
												assign node1359 = (inp[15]) ? 4'b1101 : node1360;
													assign node1360 = (inp[0]) ? 4'b1111 : 4'b1101;
										assign node1364 = (inp[7]) ? node1366 : 4'b1111;
											assign node1366 = (inp[12]) ? 4'b1000 : node1367;
												assign node1367 = (inp[10]) ? 4'b1010 : node1368;
													assign node1368 = (inp[4]) ? 4'b1011 : 4'b1010;
								assign node1373 = (inp[15]) ? node1399 : node1374;
									assign node1374 = (inp[11]) ? node1384 : node1375;
										assign node1375 = (inp[1]) ? 4'b1011 : node1376;
											assign node1376 = (inp[7]) ? 4'b1101 : node1377;
												assign node1377 = (inp[12]) ? 4'b1001 : node1378;
													assign node1378 = (inp[4]) ? 4'b1010 : 4'b1000;
										assign node1384 = (inp[9]) ? node1394 : node1385;
											assign node1385 = (inp[12]) ? node1389 : node1386;
												assign node1386 = (inp[7]) ? 4'b1100 : 4'b1010;
												assign node1389 = (inp[4]) ? node1391 : 4'b1011;
													assign node1391 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node1394 = (inp[4]) ? 4'b1011 : node1395;
												assign node1395 = (inp[12]) ? 4'b1010 : 4'b1011;
									assign node1399 = (inp[4]) ? node1413 : node1400;
										assign node1400 = (inp[0]) ? node1404 : node1401;
											assign node1401 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node1404 = (inp[10]) ? 4'b1000 : node1405;
												assign node1405 = (inp[11]) ? node1407 : 4'b1011;
													assign node1407 = (inp[9]) ? node1409 : 4'b1000;
														assign node1409 = (inp[1]) ? 4'b1011 : 4'b1010;
										assign node1413 = (inp[7]) ? 4'b1000 : node1414;
											assign node1414 = (inp[0]) ? 4'b1010 : node1415;
												assign node1415 = (inp[11]) ? 4'b1010 : 4'b1011;
					assign node1420 = (inp[1]) ? node1582 : node1421;
						assign node1421 = (inp[4]) ? node1525 : node1422;
							assign node1422 = (inp[0]) ? node1464 : node1423;
								assign node1423 = (inp[12]) ? node1445 : node1424;
									assign node1424 = (inp[9]) ? node1432 : node1425;
										assign node1425 = (inp[5]) ? 4'b0100 : node1426;
											assign node1426 = (inp[11]) ? 4'b0010 : node1427;
												assign node1427 = (inp[2]) ? 4'b0111 : 4'b0011;
										assign node1432 = (inp[10]) ? node1436 : node1433;
											assign node1433 = (inp[13]) ? 4'b0100 : 4'b0110;
											assign node1436 = (inp[13]) ? node1440 : node1437;
												assign node1437 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node1440 = (inp[15]) ? 4'b0101 : node1441;
													assign node1441 = (inp[7]) ? 4'b0101 : 4'b0011;
									assign node1445 = (inp[15]) ? node1455 : node1446;
										assign node1446 = (inp[7]) ? node1452 : node1447;
											assign node1447 = (inp[9]) ? 4'b0000 : node1448;
												assign node1448 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node1452 = (inp[2]) ? 4'b0110 : 4'b0010;
										assign node1455 = (inp[10]) ? node1459 : node1456;
											assign node1456 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node1459 = (inp[9]) ? node1461 : 4'b0001;
												assign node1461 = (inp[5]) ? 4'b0100 : 4'b0101;
								assign node1464 = (inp[9]) ? node1482 : node1465;
									assign node1465 = (inp[5]) ? node1473 : node1466;
										assign node1466 = (inp[11]) ? node1468 : 4'b0111;
											assign node1468 = (inp[7]) ? 4'b0000 : node1469;
												assign node1469 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node1473 = (inp[10]) ? node1477 : node1474;
											assign node1474 = (inp[11]) ? 4'b0011 : 4'b0111;
											assign node1477 = (inp[13]) ? node1479 : 4'b0100;
												assign node1479 = (inp[2]) ? 4'b0001 : 4'b0101;
									assign node1482 = (inp[12]) ? node1506 : node1483;
										assign node1483 = (inp[10]) ? node1497 : node1484;
											assign node1484 = (inp[11]) ? node1490 : node1485;
												assign node1485 = (inp[13]) ? 4'b0011 : node1486;
													assign node1486 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node1490 = (inp[13]) ? node1494 : node1491;
													assign node1491 = (inp[7]) ? 4'b0010 : 4'b0000;
													assign node1494 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node1497 = (inp[7]) ? node1503 : node1498;
												assign node1498 = (inp[15]) ? 4'b0101 : node1499;
													assign node1499 = (inp[5]) ? 4'b0010 : 4'b0111;
												assign node1503 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node1506 = (inp[15]) ? node1516 : node1507;
											assign node1507 = (inp[7]) ? node1511 : node1508;
												assign node1508 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node1511 = (inp[13]) ? 4'b0011 : node1512;
													assign node1512 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node1516 = (inp[13]) ? node1520 : node1517;
												assign node1517 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node1520 = (inp[10]) ? 4'b0111 : node1521;
													assign node1521 = (inp[2]) ? 4'b0110 : 4'b0010;
							assign node1525 = (inp[7]) ? node1549 : node1526;
								assign node1526 = (inp[12]) ? node1534 : node1527;
									assign node1527 = (inp[5]) ? 4'b0000 : node1528;
										assign node1528 = (inp[13]) ? 4'b0001 : node1529;
											assign node1529 = (inp[0]) ? 4'b0000 : 4'b0001;
									assign node1534 = (inp[9]) ? node1540 : node1535;
										assign node1535 = (inp[13]) ? node1537 : 4'b0110;
											assign node1537 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node1540 = (inp[15]) ? node1546 : node1541;
											assign node1541 = (inp[10]) ? 4'b0110 : node1542;
												assign node1542 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node1546 = (inp[5]) ? 4'b0011 : 4'b0111;
								assign node1549 = (inp[12]) ? node1567 : node1550;
									assign node1550 = (inp[2]) ? node1564 : node1551;
										assign node1551 = (inp[13]) ? node1555 : node1552;
											assign node1552 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node1555 = (inp[5]) ? node1557 : 4'b0010;
												assign node1557 = (inp[0]) ? node1559 : 4'b0111;
													assign node1559 = (inp[10]) ? 4'b0110 : node1560;
														assign node1560 = (inp[15]) ? 4'b0111 : 4'b0110;
										assign node1564 = (inp[9]) ? 4'b0111 : 4'b0110;
									assign node1567 = (inp[0]) ? node1573 : node1568;
										assign node1568 = (inp[2]) ? 4'b0000 : node1569;
											assign node1569 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node1573 = (inp[13]) ? node1579 : node1574;
											assign node1574 = (inp[5]) ? node1576 : 4'b0101;
												assign node1576 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node1579 = (inp[11]) ? 4'b0100 : 4'b0101;
						assign node1582 = (inp[15]) ? node1658 : node1583;
							assign node1583 = (inp[2]) ? node1621 : node1584;
								assign node1584 = (inp[11]) ? node1598 : node1585;
									assign node1585 = (inp[0]) ? node1593 : node1586;
										assign node1586 = (inp[4]) ? node1590 : node1587;
											assign node1587 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node1590 = (inp[5]) ? 4'b0000 : 4'b0110;
										assign node1593 = (inp[9]) ? 4'b0110 : node1594;
											assign node1594 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node1598 = (inp[0]) ? node1610 : node1599;
										assign node1599 = (inp[13]) ? node1605 : node1600;
											assign node1600 = (inp[5]) ? node1602 : 4'b0001;
												assign node1602 = (inp[10]) ? 4'b0010 : 4'b0111;
											assign node1605 = (inp[5]) ? node1607 : 4'b0100;
												assign node1607 = (inp[12]) ? 4'b0100 : 4'b0001;
										assign node1610 = (inp[9]) ? node1612 : 4'b0111;
											assign node1612 = (inp[10]) ? 4'b0010 : node1613;
												assign node1613 = (inp[13]) ? 4'b0011 : node1614;
													assign node1614 = (inp[4]) ? 4'b0000 : node1615;
														assign node1615 = (inp[7]) ? 4'b0011 : 4'b0000;
								assign node1621 = (inp[10]) ? node1639 : node1622;
									assign node1622 = (inp[12]) ? node1630 : node1623;
										assign node1623 = (inp[0]) ? node1625 : 4'b0111;
											assign node1625 = (inp[7]) ? node1627 : 4'b0010;
												assign node1627 = (inp[13]) ? 4'b0010 : 4'b0111;
										assign node1630 = (inp[9]) ? node1636 : node1631;
											assign node1631 = (inp[4]) ? node1633 : 4'b0101;
												assign node1633 = (inp[13]) ? 4'b0111 : 4'b0011;
											assign node1636 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1639 = (inp[0]) ? node1645 : node1640;
										assign node1640 = (inp[12]) ? 4'b0101 : node1641;
											assign node1641 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node1645 = (inp[9]) ? node1651 : node1646;
											assign node1646 = (inp[7]) ? node1648 : 4'b0100;
												assign node1648 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node1651 = (inp[11]) ? node1653 : 4'b0111;
												assign node1653 = (inp[4]) ? 4'b0111 : node1654;
													assign node1654 = (inp[12]) ? 4'b0111 : 4'b0101;
							assign node1658 = (inp[4]) ? node1686 : node1659;
								assign node1659 = (inp[12]) ? node1673 : node1660;
									assign node1660 = (inp[7]) ? node1664 : node1661;
										assign node1661 = (inp[2]) ? 4'b0100 : 4'b0000;
										assign node1664 = (inp[11]) ? node1670 : node1665;
											assign node1665 = (inp[2]) ? 4'b0010 : node1666;
												assign node1666 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node1670 = (inp[2]) ? 4'b0110 : 4'b0010;
									assign node1673 = (inp[7]) ? node1681 : node1674;
										assign node1674 = (inp[9]) ? node1676 : 4'b0111;
											assign node1676 = (inp[5]) ? node1678 : 4'b0010;
												assign node1678 = (inp[13]) ? 4'b0010 : 4'b0111;
										assign node1681 = (inp[10]) ? 4'b0101 : node1682;
											assign node1682 = (inp[2]) ? 4'b0000 : 4'b0101;
								assign node1686 = (inp[9]) ? node1702 : node1687;
									assign node1687 = (inp[5]) ? node1691 : node1688;
										assign node1688 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node1691 = (inp[2]) ? node1697 : node1692;
											assign node1692 = (inp[13]) ? node1694 : 4'b0010;
												assign node1694 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node1697 = (inp[13]) ? node1699 : 4'b0101;
												assign node1699 = (inp[10]) ? 4'b0011 : 4'b0010;
									assign node1702 = (inp[10]) ? node1710 : node1703;
										assign node1703 = (inp[7]) ? 4'b0001 : node1704;
											assign node1704 = (inp[5]) ? 4'b0111 : node1705;
												assign node1705 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node1710 = (inp[7]) ? 4'b0110 : node1711;
											assign node1711 = (inp[2]) ? 4'b0010 : 4'b0110;
				assign node1715 = (inp[12]) ? node1975 : node1716;
					assign node1716 = (inp[15]) ? node1846 : node1717;
						assign node1717 = (inp[14]) ? node1797 : node1718;
							assign node1718 = (inp[4]) ? node1746 : node1719;
								assign node1719 = (inp[9]) ? node1739 : node1720;
									assign node1720 = (inp[0]) ? node1732 : node1721;
										assign node1721 = (inp[10]) ? 4'b0001 : node1722;
											assign node1722 = (inp[5]) ? 4'b0100 : node1723;
												assign node1723 = (inp[11]) ? 4'b0000 : node1724;
													assign node1724 = (inp[13]) ? 4'b0001 : node1725;
														assign node1725 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node1732 = (inp[1]) ? node1734 : 4'b0001;
											assign node1734 = (inp[7]) ? node1736 : 4'b0101;
												assign node1736 = (inp[2]) ? 4'b0001 : 4'b0101;
									assign node1739 = (inp[1]) ? node1743 : node1740;
										assign node1740 = (inp[2]) ? 4'b0100 : 4'b0000;
										assign node1743 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node1746 = (inp[9]) ? node1780 : node1747;
									assign node1747 = (inp[1]) ? node1755 : node1748;
										assign node1748 = (inp[10]) ? 4'b0000 : node1749;
											assign node1749 = (inp[0]) ? 4'b0000 : node1750;
												assign node1750 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node1755 = (inp[13]) ? node1771 : node1756;
											assign node1756 = (inp[11]) ? node1762 : node1757;
												assign node1757 = (inp[5]) ? 4'b0100 : node1758;
													assign node1758 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node1762 = (inp[7]) ? node1764 : 4'b0101;
													assign node1764 = (inp[10]) ? 4'b0000 : node1765;
														assign node1765 = (inp[2]) ? 4'b0000 : node1766;
															assign node1766 = (inp[5]) ? 4'b0001 : 4'b0101;
											assign node1771 = (inp[7]) ? 4'b0001 : node1772;
												assign node1772 = (inp[10]) ? 4'b0000 : node1773;
													assign node1773 = (inp[2]) ? 4'b0100 : node1774;
														assign node1774 = (inp[0]) ? 4'b0100 : 4'b0001;
									assign node1780 = (inp[5]) ? node1792 : node1781;
										assign node1781 = (inp[10]) ? 4'b0001 : node1782;
											assign node1782 = (inp[13]) ? node1788 : node1783;
												assign node1783 = (inp[0]) ? node1785 : 4'b0101;
													assign node1785 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node1788 = (inp[1]) ? 4'b0001 : 4'b0101;
										assign node1792 = (inp[11]) ? node1794 : 4'b0101;
											assign node1794 = (inp[13]) ? 4'b0100 : 4'b0101;
							assign node1797 = (inp[7]) ? node1823 : node1798;
								assign node1798 = (inp[2]) ? node1808 : node1799;
									assign node1799 = (inp[5]) ? node1805 : node1800;
										assign node1800 = (inp[9]) ? 4'b0010 : node1801;
											assign node1801 = (inp[4]) ? 4'b0011 : 4'b0010;
										assign node1805 = (inp[4]) ? 4'b0010 : 4'b0110;
									assign node1808 = (inp[0]) ? node1814 : node1809;
										assign node1809 = (inp[4]) ? 4'b0111 : node1810;
											assign node1810 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node1814 = (inp[5]) ? node1820 : node1815;
											assign node1815 = (inp[9]) ? node1817 : 4'b0110;
												assign node1817 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node1820 = (inp[4]) ? 4'b0111 : 4'b0010;
								assign node1823 = (inp[2]) ? node1835 : node1824;
									assign node1824 = (inp[13]) ? node1830 : node1825;
										assign node1825 = (inp[4]) ? 4'b0111 : node1826;
											assign node1826 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node1830 = (inp[11]) ? 4'b0010 : node1831;
											assign node1831 = (inp[4]) ? 4'b0110 : 4'b0111;
									assign node1835 = (inp[5]) ? node1843 : node1836;
										assign node1836 = (inp[1]) ? 4'b0011 : node1837;
											assign node1837 = (inp[4]) ? 4'b0010 : node1838;
												assign node1838 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node1843 = (inp[4]) ? 4'b0011 : 4'b0111;
						assign node1846 = (inp[9]) ? node1910 : node1847;
							assign node1847 = (inp[14]) ? node1879 : node1848;
								assign node1848 = (inp[7]) ? node1866 : node1849;
									assign node1849 = (inp[4]) ? node1855 : node1850;
										assign node1850 = (inp[0]) ? 4'b0110 : node1851;
											assign node1851 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node1855 = (inp[2]) ? node1859 : node1856;
											assign node1856 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node1859 = (inp[13]) ? node1861 : 4'b0010;
												assign node1861 = (inp[10]) ? node1863 : 4'b0011;
													assign node1863 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node1866 = (inp[4]) ? node1872 : node1867;
										assign node1867 = (inp[2]) ? 4'b0111 : node1868;
											assign node1868 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node1872 = (inp[2]) ? node1876 : node1873;
											assign node1873 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node1876 = (inp[13]) ? 4'b0011 : 4'b0010;
								assign node1879 = (inp[7]) ? node1891 : node1880;
									assign node1880 = (inp[11]) ? node1888 : node1881;
										assign node1881 = (inp[2]) ? node1883 : 4'b0011;
											assign node1883 = (inp[5]) ? node1885 : 4'b0011;
												assign node1885 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node1888 = (inp[0]) ? 4'b0110 : 4'b0010;
									assign node1891 = (inp[5]) ? node1901 : node1892;
										assign node1892 = (inp[0]) ? node1898 : node1893;
											assign node1893 = (inp[4]) ? node1895 : 4'b0110;
												assign node1895 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node1898 = (inp[4]) ? 4'b0110 : 4'b0111;
										assign node1901 = (inp[0]) ? node1907 : node1902;
											assign node1902 = (inp[4]) ? 4'b0110 : node1903;
												assign node1903 = (inp[11]) ? 4'b0110 : 4'b0010;
											assign node1907 = (inp[1]) ? 4'b0011 : 4'b0010;
							assign node1910 = (inp[13]) ? node1950 : node1911;
								assign node1911 = (inp[11]) ? node1923 : node1912;
									assign node1912 = (inp[0]) ? node1920 : node1913;
										assign node1913 = (inp[10]) ? node1915 : 4'b0011;
											assign node1915 = (inp[1]) ? 4'b0110 : node1916;
												assign node1916 = (inp[14]) ? 4'b0011 : 4'b0111;
										assign node1920 = (inp[14]) ? 4'b0111 : 4'b0011;
									assign node1923 = (inp[2]) ? node1937 : node1924;
										assign node1924 = (inp[4]) ? node1932 : node1925;
											assign node1925 = (inp[7]) ? 4'b0011 : node1926;
												assign node1926 = (inp[1]) ? 4'b0010 : node1927;
													assign node1927 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node1932 = (inp[10]) ? 4'b0110 : node1933;
												assign node1933 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node1937 = (inp[4]) ? node1947 : node1938;
											assign node1938 = (inp[5]) ? node1940 : 4'b0111;
												assign node1940 = (inp[7]) ? 4'b0111 : node1941;
													assign node1941 = (inp[10]) ? 4'b0110 : node1942;
														assign node1942 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node1947 = (inp[1]) ? 4'b0011 : 4'b0010;
								assign node1950 = (inp[4]) ? node1966 : node1951;
									assign node1951 = (inp[2]) ? node1959 : node1952;
										assign node1952 = (inp[0]) ? node1954 : 4'b0011;
											assign node1954 = (inp[7]) ? node1956 : 4'b0010;
												assign node1956 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node1959 = (inp[11]) ? node1961 : 4'b0110;
											assign node1961 = (inp[0]) ? 4'b0111 : node1962;
												assign node1962 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node1966 = (inp[2]) ? node1970 : node1967;
										assign node1967 = (inp[14]) ? 4'b0111 : 4'b0110;
										assign node1970 = (inp[7]) ? node1972 : 4'b0011;
											assign node1972 = (inp[5]) ? 4'b0011 : 4'b0010;
					assign node1975 = (inp[14]) ? node2077 : node1976;
						assign node1976 = (inp[15]) ? node2034 : node1977;
							assign node1977 = (inp[4]) ? node2011 : node1978;
								assign node1978 = (inp[9]) ? node1990 : node1979;
									assign node1979 = (inp[7]) ? node1985 : node1980;
										assign node1980 = (inp[2]) ? node1982 : 4'b0011;
											assign node1982 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node1985 = (inp[2]) ? node1987 : 4'b0111;
											assign node1987 = (inp[11]) ? 4'b0011 : 4'b0010;
									assign node1990 = (inp[7]) ? node2002 : node1991;
										assign node1991 = (inp[2]) ? node1999 : node1992;
											assign node1992 = (inp[5]) ? 4'b0010 : node1993;
												assign node1993 = (inp[11]) ? 4'b0011 : node1994;
													assign node1994 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node1999 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node2002 = (inp[5]) ? node2006 : node2003;
											assign node2003 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node2006 = (inp[0]) ? node2008 : 4'b0111;
												assign node2008 = (inp[1]) ? 4'b0111 : 4'b0110;
								assign node2011 = (inp[5]) ? node2021 : node2012;
									assign node2012 = (inp[11]) ? 4'b0111 : node2013;
										assign node2013 = (inp[1]) ? 4'b0110 : node2014;
											assign node2014 = (inp[9]) ? node2016 : 4'b0010;
												assign node2016 = (inp[2]) ? 4'b0010 : 4'b0111;
									assign node2021 = (inp[13]) ? node2027 : node2022;
										assign node2022 = (inp[7]) ? node2024 : 4'b0010;
											assign node2024 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node2027 = (inp[7]) ? node2031 : node2028;
											assign node2028 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node2031 = (inp[10]) ? 4'b0010 : 4'b0110;
							assign node2034 = (inp[4]) ? node2058 : node2035;
								assign node2035 = (inp[0]) ? node2049 : node2036;
									assign node2036 = (inp[10]) ? node2042 : node2037;
										assign node2037 = (inp[9]) ? 4'b0000 : node2038;
											assign node2038 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node2042 = (inp[7]) ? node2044 : 4'b0101;
											assign node2044 = (inp[1]) ? 4'b0101 : node2045;
												assign node2045 = (inp[11]) ? 4'b0000 : 4'b0100;
									assign node2049 = (inp[5]) ? node2053 : node2050;
										assign node2050 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node2053 = (inp[2]) ? 4'b0000 : node2054;
											assign node2054 = (inp[1]) ? 4'b0101 : 4'b0100;
								assign node2058 = (inp[13]) ? node2066 : node2059;
									assign node2059 = (inp[10]) ? 4'b0100 : node2060;
										assign node2060 = (inp[11]) ? node2062 : 4'b0101;
											assign node2062 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node2066 = (inp[5]) ? node2072 : node2067;
										assign node2067 = (inp[2]) ? 4'b0101 : node2068;
											assign node2068 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node2072 = (inp[2]) ? node2074 : 4'b0101;
											assign node2074 = (inp[9]) ? 4'b0000 : 4'b0001;
						assign node2077 = (inp[2]) ? node2125 : node2078;
							assign node2078 = (inp[15]) ? node2108 : node2079;
								assign node2079 = (inp[7]) ? node2089 : node2080;
									assign node2080 = (inp[4]) ? node2086 : node2081;
										assign node2081 = (inp[5]) ? 4'b0000 : node2082;
											assign node2082 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node2086 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node2089 = (inp[5]) ? node2095 : node2090;
										assign node2090 = (inp[4]) ? 4'b0100 : node2091;
											assign node2091 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node2095 = (inp[0]) ? node2103 : node2096;
											assign node2096 = (inp[1]) ? node2098 : 4'b0101;
												assign node2098 = (inp[10]) ? 4'b0100 : node2099;
													assign node2099 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node2103 = (inp[4]) ? node2105 : 4'b0100;
												assign node2105 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node2108 = (inp[7]) ? node2120 : node2109;
									assign node2109 = (inp[11]) ? node2113 : node2110;
										assign node2110 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node2113 = (inp[10]) ? node2115 : 4'b0100;
											assign node2115 = (inp[4]) ? 4'b0100 : node2116;
												assign node2116 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node2120 = (inp[10]) ? node2122 : 4'b0101;
										assign node2122 = (inp[5]) ? 4'b0101 : 4'b0100;
							assign node2125 = (inp[15]) ? node2153 : node2126;
								assign node2126 = (inp[7]) ? node2144 : node2127;
									assign node2127 = (inp[5]) ? node2133 : node2128;
										assign node2128 = (inp[4]) ? node2130 : 4'b0001;
											assign node2130 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node2133 = (inp[4]) ? node2139 : node2134;
											assign node2134 = (inp[1]) ? node2136 : 4'b0100;
												assign node2136 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node2139 = (inp[0]) ? node2141 : 4'b0101;
												assign node2141 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node2144 = (inp[5]) ? node2150 : node2145;
										assign node2145 = (inp[13]) ? 4'b0101 : node2146;
											assign node2146 = (inp[4]) ? 4'b0001 : 4'b0100;
										assign node2150 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node2153 = (inp[10]) ? node2163 : node2154;
									assign node2154 = (inp[7]) ? 4'b0001 : node2155;
										assign node2155 = (inp[5]) ? 4'b0001 : node2156;
											assign node2156 = (inp[11]) ? 4'b0000 : node2157;
												assign node2157 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node2163 = (inp[5]) ? 4'b0000 : node2164;
										assign node2164 = (inp[7]) ? node2166 : 4'b0001;
											assign node2166 = (inp[0]) ? 4'b0000 : node2167;
												assign node2167 = (inp[1]) ? 4'b0000 : 4'b0001;
		assign node2172 = (inp[14]) ? node3262 : node2173;
			assign node2173 = (inp[8]) ? node2781 : node2174;
				assign node2174 = (inp[1]) ? node2500 : node2175;
					assign node2175 = (inp[2]) ? node2325 : node2176;
						assign node2176 = (inp[9]) ? node2254 : node2177;
							assign node2177 = (inp[11]) ? node2223 : node2178;
								assign node2178 = (inp[4]) ? node2194 : node2179;
									assign node2179 = (inp[3]) ? node2185 : node2180;
										assign node2180 = (inp[5]) ? 4'b1010 : node2181;
											assign node2181 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node2185 = (inp[0]) ? 4'b1100 : node2186;
											assign node2186 = (inp[13]) ? 4'b1001 : node2187;
												assign node2187 = (inp[12]) ? node2189 : 4'b1010;
													assign node2189 = (inp[15]) ? 4'b1100 : 4'b1000;
									assign node2194 = (inp[3]) ? node2210 : node2195;
										assign node2195 = (inp[7]) ? node2207 : node2196;
											assign node2196 = (inp[15]) ? node2202 : node2197;
												assign node2197 = (inp[0]) ? node2199 : 4'b1100;
													assign node2199 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node2202 = (inp[10]) ? 4'b1110 : node2203;
													assign node2203 = (inp[13]) ? 4'b1110 : 4'b1010;
											assign node2207 = (inp[13]) ? 4'b1100 : 4'b1001;
										assign node2210 = (inp[10]) ? node2214 : node2211;
											assign node2211 = (inp[13]) ? 4'b1110 : 4'b1010;
											assign node2214 = (inp[0]) ? 4'b1111 : node2215;
												assign node2215 = (inp[5]) ? 4'b1110 : node2216;
													assign node2216 = (inp[13]) ? 4'b1100 : node2217;
														assign node2217 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node2223 = (inp[13]) ? node2243 : node2224;
									assign node2224 = (inp[0]) ? node2236 : node2225;
										assign node2225 = (inp[10]) ? node2231 : node2226;
											assign node2226 = (inp[12]) ? 4'b1111 : node2227;
												assign node2227 = (inp[5]) ? 4'b1001 : 4'b1111;
											assign node2231 = (inp[3]) ? node2233 : 4'b1000;
												assign node2233 = (inp[5]) ? 4'b1111 : 4'b1010;
										assign node2236 = (inp[12]) ? 4'b1000 : node2237;
											assign node2237 = (inp[7]) ? 4'b1110 : node2238;
												assign node2238 = (inp[5]) ? 4'b1100 : 4'b1000;
									assign node2243 = (inp[5]) ? node2247 : node2244;
										assign node2244 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node2247 = (inp[7]) ? 4'b1111 : node2248;
											assign node2248 = (inp[12]) ? 4'b1100 : node2249;
												assign node2249 = (inp[15]) ? 4'b1010 : 4'b1000;
							assign node2254 = (inp[4]) ? node2286 : node2255;
								assign node2255 = (inp[13]) ? node2273 : node2256;
									assign node2256 = (inp[5]) ? node2268 : node2257;
										assign node2257 = (inp[11]) ? 4'b1000 : node2258;
											assign node2258 = (inp[10]) ? node2262 : node2259;
												assign node2259 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node2262 = (inp[12]) ? 4'b1010 : node2263;
													assign node2263 = (inp[3]) ? 4'b1010 : 4'b1011;
										assign node2268 = (inp[7]) ? node2270 : 4'b1111;
											assign node2270 = (inp[10]) ? 4'b1000 : 4'b1110;
									assign node2273 = (inp[0]) ? 4'b1111 : node2274;
										assign node2274 = (inp[15]) ? node2282 : node2275;
											assign node2275 = (inp[12]) ? node2277 : 4'b1000;
												assign node2277 = (inp[3]) ? 4'b1001 : node2278;
													assign node2278 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node2282 = (inp[10]) ? 4'b1011 : 4'b1001;
								assign node2286 = (inp[7]) ? node2308 : node2287;
									assign node2287 = (inp[15]) ? node2291 : node2288;
										assign node2288 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node2291 = (inp[11]) ? node2301 : node2292;
											assign node2292 = (inp[0]) ? node2298 : node2293;
												assign node2293 = (inp[5]) ? node2295 : 4'b1111;
													assign node2295 = (inp[3]) ? 4'b1110 : 4'b1111;
												assign node2298 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node2301 = (inp[10]) ? node2303 : 4'b1111;
												assign node2303 = (inp[13]) ? node2305 : 4'b1010;
													assign node2305 = (inp[3]) ? 4'b1011 : 4'b1010;
									assign node2308 = (inp[15]) ? node2314 : node2309;
										assign node2309 = (inp[12]) ? 4'b1111 : node2310;
											assign node2310 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node2314 = (inp[12]) ? node2320 : node2315;
											assign node2315 = (inp[5]) ? 4'b1100 : node2316;
												assign node2316 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node2320 = (inp[10]) ? 4'b1100 : node2321;
												assign node2321 = (inp[11]) ? 4'b1100 : 4'b1000;
						assign node2325 = (inp[3]) ? node2399 : node2326;
							assign node2326 = (inp[10]) ? node2368 : node2327;
								assign node2327 = (inp[9]) ? node2349 : node2328;
									assign node2328 = (inp[11]) ? node2342 : node2329;
										assign node2329 = (inp[7]) ? node2337 : node2330;
											assign node2330 = (inp[15]) ? node2332 : 4'b1101;
												assign node2332 = (inp[5]) ? node2334 : 4'b1111;
													assign node2334 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node2337 = (inp[15]) ? node2339 : 4'b1111;
												assign node2339 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node2342 = (inp[12]) ? node2346 : node2343;
											assign node2343 = (inp[13]) ? 4'b1111 : 4'b1010;
											assign node2346 = (inp[0]) ? 4'b1100 : 4'b1001;
									assign node2349 = (inp[15]) ? node2357 : node2350;
										assign node2350 = (inp[7]) ? node2354 : node2351;
											assign node2351 = (inp[13]) ? 4'b1001 : 4'b1100;
											assign node2354 = (inp[5]) ? 4'b1111 : 4'b1011;
										assign node2357 = (inp[7]) ? 4'b1000 : node2358;
											assign node2358 = (inp[4]) ? node2360 : 4'b1111;
												assign node2360 = (inp[13]) ? node2362 : 4'b1110;
													assign node2362 = (inp[11]) ? node2364 : 4'b1010;
														assign node2364 = (inp[12]) ? 4'b1010 : 4'b1011;
								assign node2368 = (inp[11]) ? node2394 : node2369;
									assign node2369 = (inp[5]) ? node2379 : node2370;
										assign node2370 = (inp[13]) ? node2376 : node2371;
											assign node2371 = (inp[7]) ? 4'b1011 : node2372;
												assign node2372 = (inp[4]) ? 4'b1000 : 4'b1011;
											assign node2376 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node2379 = (inp[13]) ? node2385 : node2380;
											assign node2380 = (inp[4]) ? node2382 : 4'b1110;
												assign node2382 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node2385 = (inp[12]) ? node2391 : node2386;
												assign node2386 = (inp[9]) ? node2388 : 4'b1010;
													assign node2388 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node2391 = (inp[15]) ? 4'b1011 : 4'b1010;
									assign node2394 = (inp[4]) ? 4'b1110 : node2395;
										assign node2395 = (inp[13]) ? 4'b1011 : 4'b1111;
							assign node2399 = (inp[9]) ? node2447 : node2400;
								assign node2400 = (inp[4]) ? node2432 : node2401;
									assign node2401 = (inp[15]) ? node2413 : node2402;
										assign node2402 = (inp[7]) ? node2408 : node2403;
											assign node2403 = (inp[13]) ? 4'b1101 : node2404;
												assign node2404 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node2408 = (inp[12]) ? node2410 : 4'b1011;
												assign node2410 = (inp[13]) ? 4'b1011 : 4'b1110;
										assign node2413 = (inp[7]) ? node2429 : node2414;
											assign node2414 = (inp[11]) ? node2424 : node2415;
												assign node2415 = (inp[10]) ? node2421 : node2416;
													assign node2416 = (inp[0]) ? node2418 : 4'b1110;
														assign node2418 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node2421 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node2424 = (inp[10]) ? node2426 : 4'b1111;
													assign node2426 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node2429 = (inp[10]) ? 4'b1000 : 4'b1001;
									assign node2432 = (inp[15]) ? node2440 : node2433;
										assign node2433 = (inp[13]) ? node2437 : node2434;
											assign node2434 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node2437 = (inp[12]) ? 4'b1101 : 4'b1001;
										assign node2440 = (inp[11]) ? node2444 : node2441;
											assign node2441 = (inp[5]) ? 4'b1000 : 4'b1100;
											assign node2444 = (inp[13]) ? 4'b1001 : 4'b1000;
								assign node2447 = (inp[0]) ? node2479 : node2448;
									assign node2448 = (inp[15]) ? node2464 : node2449;
										assign node2449 = (inp[12]) ? node2457 : node2450;
											assign node2450 = (inp[7]) ? 4'b1110 : node2451;
												assign node2451 = (inp[5]) ? node2453 : 4'b1100;
													assign node2453 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node2457 = (inp[10]) ? node2461 : node2458;
												assign node2458 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node2461 = (inp[5]) ? 4'b1100 : 4'b1000;
										assign node2464 = (inp[7]) ? node2466 : 4'b1010;
											assign node2466 = (inp[12]) ? node2474 : node2467;
												assign node2467 = (inp[11]) ? node2469 : 4'b1001;
													assign node2469 = (inp[10]) ? 4'b1001 : node2470;
														assign node2470 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node2474 = (inp[13]) ? 4'b1000 : node2475;
													assign node2475 = (inp[5]) ? 4'b1100 : 4'b1000;
									assign node2479 = (inp[13]) ? node2487 : node2480;
										assign node2480 = (inp[15]) ? node2482 : 4'b1100;
											assign node2482 = (inp[5]) ? 4'b1110 : node2483;
												assign node2483 = (inp[11]) ? 4'b1010 : 4'b1110;
										assign node2487 = (inp[5]) ? 4'b1000 : node2488;
											assign node2488 = (inp[10]) ? node2492 : node2489;
												assign node2489 = (inp[12]) ? 4'b1101 : 4'b1000;
												assign node2492 = (inp[11]) ? node2494 : 4'b1111;
													assign node2494 = (inp[7]) ? 4'b1100 : node2495;
														assign node2495 = (inp[12]) ? 4'b1100 : 4'b1111;
					assign node2500 = (inp[0]) ? node2652 : node2501;
						assign node2501 = (inp[13]) ? node2573 : node2502;
							assign node2502 = (inp[5]) ? node2542 : node2503;
								assign node2503 = (inp[15]) ? node2527 : node2504;
									assign node2504 = (inp[7]) ? node2524 : node2505;
										assign node2505 = (inp[10]) ? node2515 : node2506;
											assign node2506 = (inp[3]) ? node2508 : 4'b1001;
												assign node2508 = (inp[9]) ? node2510 : 4'b1000;
													assign node2510 = (inp[12]) ? node2512 : 4'b1001;
														assign node2512 = (inp[11]) ? 4'b1001 : 4'b1100;
											assign node2515 = (inp[11]) ? node2517 : 4'b1101;
												assign node2517 = (inp[2]) ? 4'b1000 : node2518;
													assign node2518 = (inp[3]) ? 4'b1001 : node2519;
														assign node2519 = (inp[12]) ? 4'b1100 : 4'b1001;
										assign node2524 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node2527 = (inp[7]) ? node2537 : node2528;
										assign node2528 = (inp[12]) ? node2530 : 4'b1111;
											assign node2530 = (inp[4]) ? 4'b1011 : node2531;
												assign node2531 = (inp[2]) ? 4'b1011 : node2532;
													assign node2532 = (inp[3]) ? 4'b1010 : 4'b1110;
										assign node2537 = (inp[11]) ? node2539 : 4'b1001;
											assign node2539 = (inp[9]) ? 4'b1001 : 4'b1000;
								assign node2542 = (inp[12]) ? node2552 : node2543;
									assign node2543 = (inp[2]) ? node2547 : node2544;
										assign node2544 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node2547 = (inp[10]) ? node2549 : 4'b1111;
											assign node2549 = (inp[3]) ? 4'b1001 : 4'b1101;
									assign node2552 = (inp[3]) ? node2562 : node2553;
										assign node2553 = (inp[4]) ? node2559 : node2554;
											assign node2554 = (inp[7]) ? node2556 : 4'b1001;
												assign node2556 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node2559 = (inp[7]) ? 4'b1110 : 4'b1100;
										assign node2562 = (inp[9]) ? node2568 : node2563;
											assign node2563 = (inp[2]) ? 4'b1111 : node2564;
												assign node2564 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node2568 = (inp[15]) ? node2570 : 4'b1111;
												assign node2570 = (inp[2]) ? 4'b1101 : 4'b1100;
							assign node2573 = (inp[11]) ? node2617 : node2574;
								assign node2574 = (inp[9]) ? node2590 : node2575;
									assign node2575 = (inp[15]) ? node2585 : node2576;
										assign node2576 = (inp[7]) ? node2578 : 4'b1101;
											assign node2578 = (inp[4]) ? node2580 : 4'b1010;
												assign node2580 = (inp[5]) ? node2582 : 4'b1111;
													assign node2582 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node2585 = (inp[7]) ? 4'b1001 : node2586;
											assign node2586 = (inp[5]) ? 4'b1010 : 4'b1011;
									assign node2590 = (inp[7]) ? node2604 : node2591;
										assign node2591 = (inp[15]) ? node2601 : node2592;
											assign node2592 = (inp[5]) ? 4'b1001 : node2593;
												assign node2593 = (inp[12]) ? node2595 : 4'b1000;
													assign node2595 = (inp[4]) ? 4'b1001 : node2596;
														assign node2596 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node2601 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node2604 = (inp[15]) ? node2614 : node2605;
											assign node2605 = (inp[2]) ? node2609 : node2606;
												assign node2606 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node2609 = (inp[3]) ? 4'b1110 : node2610;
													assign node2610 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node2614 = (inp[5]) ? 4'b1000 : 4'b1100;
								assign node2617 = (inp[5]) ? node2633 : node2618;
									assign node2618 = (inp[7]) ? node2630 : node2619;
										assign node2619 = (inp[15]) ? node2625 : node2620;
											assign node2620 = (inp[12]) ? 4'b1001 : node2621;
												assign node2621 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node2625 = (inp[2]) ? node2627 : 4'b1110;
												assign node2627 = (inp[10]) ? 4'b1111 : 4'b1110;
										assign node2630 = (inp[3]) ? 4'b1001 : 4'b1101;
									assign node2633 = (inp[3]) ? node2649 : node2634;
										assign node2634 = (inp[9]) ? node2640 : node2635;
											assign node2635 = (inp[4]) ? 4'b1111 : node2636;
												assign node2636 = (inp[2]) ? 4'b1110 : 4'b1010;
											assign node2640 = (inp[4]) ? node2644 : node2641;
												assign node2641 = (inp[12]) ? 4'b1111 : 4'b1010;
												assign node2644 = (inp[10]) ? node2646 : 4'b1010;
													assign node2646 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node2649 = (inp[7]) ? 4'b1000 : 4'b1100;
						assign node2652 = (inp[15]) ? node2716 : node2653;
							assign node2653 = (inp[7]) ? node2673 : node2654;
								assign node2654 = (inp[11]) ? node2668 : node2655;
									assign node2655 = (inp[13]) ? node2657 : 4'b1000;
										assign node2657 = (inp[2]) ? node2659 : 4'b1101;
											assign node2659 = (inp[3]) ? node2661 : 4'b1101;
												assign node2661 = (inp[10]) ? node2663 : 4'b1001;
													assign node2663 = (inp[12]) ? node2665 : 4'b1001;
														assign node2665 = (inp[4]) ? 4'b1100 : 4'b1001;
									assign node2668 = (inp[3]) ? 4'b1101 : node2669;
										assign node2669 = (inp[4]) ? 4'b1101 : 4'b1001;
								assign node2673 = (inp[4]) ? node2699 : node2674;
									assign node2674 = (inp[2]) ? node2688 : node2675;
										assign node2675 = (inp[13]) ? node2681 : node2676;
											assign node2676 = (inp[9]) ? 4'b1011 : node2677;
												assign node2677 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node2681 = (inp[9]) ? node2685 : node2682;
												assign node2682 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node2685 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node2688 = (inp[5]) ? node2694 : node2689;
											assign node2689 = (inp[13]) ? node2691 : 4'b1010;
												assign node2691 = (inp[3]) ? 4'b1110 : 4'b1010;
											assign node2694 = (inp[3]) ? 4'b1011 : node2695;
												assign node2695 = (inp[13]) ? 4'b1111 : 4'b1011;
									assign node2699 = (inp[12]) ? node2709 : node2700;
										assign node2700 = (inp[13]) ? node2706 : node2701;
											assign node2701 = (inp[10]) ? 4'b1110 : node2702;
												assign node2702 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node2706 = (inp[5]) ? 4'b1011 : 4'b1110;
										assign node2709 = (inp[5]) ? 4'b1111 : node2710;
											assign node2710 = (inp[13]) ? 4'b1111 : node2711;
												assign node2711 = (inp[11]) ? 4'b1011 : 4'b1010;
							assign node2716 = (inp[7]) ? node2756 : node2717;
								assign node2717 = (inp[5]) ? node2739 : node2718;
									assign node2718 = (inp[4]) ? node2728 : node2719;
										assign node2719 = (inp[2]) ? node2721 : 4'b1110;
											assign node2721 = (inp[12]) ? 4'b1111 : node2722;
												assign node2722 = (inp[10]) ? 4'b1110 : node2723;
													assign node2723 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node2728 = (inp[13]) ? node2730 : 4'b1011;
											assign node2730 = (inp[3]) ? node2734 : node2731;
												assign node2731 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node2734 = (inp[9]) ? node2736 : 4'b1111;
													assign node2736 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node2739 = (inp[4]) ? node2747 : node2740;
										assign node2740 = (inp[11]) ? node2742 : 4'b1010;
											assign node2742 = (inp[12]) ? node2744 : 4'b1111;
												assign node2744 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node2747 = (inp[11]) ? node2751 : node2748;
											assign node2748 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node2751 = (inp[12]) ? 4'b1011 : node2752;
												assign node2752 = (inp[13]) ? 4'b1110 : 4'b1011;
								assign node2756 = (inp[12]) ? node2768 : node2757;
									assign node2757 = (inp[13]) ? node2759 : 4'b1001;
										assign node2759 = (inp[5]) ? node2763 : node2760;
											assign node2760 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node2763 = (inp[4]) ? 4'b1000 : node2764;
												assign node2764 = (inp[3]) ? 4'b1100 : 4'b1000;
									assign node2768 = (inp[2]) ? node2776 : node2769;
										assign node2769 = (inp[9]) ? 4'b1101 : node2770;
											assign node2770 = (inp[4]) ? 4'b1001 : node2771;
												assign node2771 = (inp[5]) ? 4'b1101 : 4'b1001;
										assign node2776 = (inp[3]) ? 4'b1100 : node2777;
											assign node2777 = (inp[10]) ? 4'b1001 : 4'b1000;
				assign node2781 = (inp[15]) ? node3023 : node2782;
					assign node2782 = (inp[3]) ? node2892 : node2783;
						assign node2783 = (inp[4]) ? node2835 : node2784;
							assign node2784 = (inp[1]) ? node2816 : node2785;
								assign node2785 = (inp[5]) ? node2797 : node2786;
									assign node2786 = (inp[12]) ? node2794 : node2787;
										assign node2787 = (inp[0]) ? node2789 : 4'b0000;
											assign node2789 = (inp[11]) ? node2791 : 4'b0001;
												assign node2791 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node2794 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node2797 = (inp[12]) ? node2811 : node2798;
										assign node2798 = (inp[0]) ? node2806 : node2799;
											assign node2799 = (inp[7]) ? node2801 : 4'b0101;
												assign node2801 = (inp[13]) ? node2803 : 4'b0101;
													assign node2803 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node2806 = (inp[7]) ? node2808 : 4'b0100;
												assign node2808 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node2811 = (inp[7]) ? node2813 : 4'b0100;
											assign node2813 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node2816 = (inp[5]) ? node2828 : node2817;
									assign node2817 = (inp[12]) ? node2823 : node2818;
										assign node2818 = (inp[13]) ? node2820 : 4'b0100;
											assign node2820 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node2823 = (inp[9]) ? 4'b0000 : node2824;
											assign node2824 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node2828 = (inp[7]) ? node2830 : 4'b0000;
										assign node2830 = (inp[12]) ? node2832 : 4'b0000;
											assign node2832 = (inp[2]) ? 4'b0101 : 4'b0100;
							assign node2835 = (inp[12]) ? node2859 : node2836;
								assign node2836 = (inp[11]) ? node2852 : node2837;
									assign node2837 = (inp[0]) ? node2845 : node2838;
										assign node2838 = (inp[5]) ? 4'b0111 : node2839;
											assign node2839 = (inp[10]) ? 4'b0110 : node2840;
												assign node2840 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node2845 = (inp[9]) ? 4'b0011 : node2846;
											assign node2846 = (inp[13]) ? 4'b0111 : node2847;
												assign node2847 = (inp[2]) ? 4'b0110 : 4'b0111;
									assign node2852 = (inp[0]) ? 4'b0010 : node2853;
										assign node2853 = (inp[10]) ? node2855 : 4'b0011;
											assign node2855 = (inp[9]) ? 4'b0111 : 4'b0010;
								assign node2859 = (inp[11]) ? node2877 : node2860;
									assign node2860 = (inp[9]) ? node2868 : node2861;
										assign node2861 = (inp[0]) ? node2863 : 4'b0110;
											assign node2863 = (inp[5]) ? node2865 : 4'b0111;
												assign node2865 = (inp[2]) ? 4'b0111 : 4'b0011;
										assign node2868 = (inp[0]) ? node2874 : node2869;
											assign node2869 = (inp[1]) ? node2871 : 4'b0011;
												assign node2871 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node2874 = (inp[1]) ? 4'b0010 : 4'b0110;
									assign node2877 = (inp[7]) ? node2883 : node2878;
										assign node2878 = (inp[1]) ? node2880 : 4'b0111;
											assign node2880 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node2883 = (inp[13]) ? 4'b0010 : node2884;
											assign node2884 = (inp[0]) ? node2886 : 4'b0111;
												assign node2886 = (inp[9]) ? node2888 : 4'b0011;
													assign node2888 = (inp[1]) ? 4'b0111 : 4'b0011;
						assign node2892 = (inp[9]) ? node2956 : node2893;
							assign node2893 = (inp[2]) ? node2925 : node2894;
								assign node2894 = (inp[10]) ? node2916 : node2895;
									assign node2895 = (inp[12]) ? node2909 : node2896;
										assign node2896 = (inp[7]) ? node2900 : node2897;
											assign node2897 = (inp[0]) ? 4'b0111 : 4'b0011;
											assign node2900 = (inp[5]) ? 4'b0010 : node2901;
												assign node2901 = (inp[11]) ? node2905 : node2902;
													assign node2902 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node2905 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node2909 = (inp[0]) ? node2911 : 4'b0110;
											assign node2911 = (inp[11]) ? 4'b0110 : node2912;
												assign node2912 = (inp[1]) ? 4'b0011 : 4'b0010;
									assign node2916 = (inp[4]) ? 4'b0010 : node2917;
										assign node2917 = (inp[12]) ? 4'b0110 : node2918;
											assign node2918 = (inp[7]) ? 4'b0010 : node2919;
												assign node2919 = (inp[5]) ? 4'b0110 : 4'b0010;
								assign node2925 = (inp[10]) ? node2941 : node2926;
									assign node2926 = (inp[4]) ? node2936 : node2927;
										assign node2927 = (inp[0]) ? node2933 : node2928;
											assign node2928 = (inp[11]) ? node2930 : 4'b0111;
												assign node2930 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node2933 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node2936 = (inp[5]) ? node2938 : 4'b0010;
											assign node2938 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node2941 = (inp[13]) ? node2945 : node2942;
										assign node2942 = (inp[12]) ? 4'b0010 : 4'b0111;
										assign node2945 = (inp[0]) ? node2951 : node2946;
											assign node2946 = (inp[4]) ? node2948 : 4'b0010;
												assign node2948 = (inp[5]) ? 4'b0010 : 4'b0111;
											assign node2951 = (inp[12]) ? 4'b0111 : node2952;
												assign node2952 = (inp[4]) ? 4'b0111 : 4'b0110;
							assign node2956 = (inp[12]) ? node2984 : node2957;
								assign node2957 = (inp[4]) ? node2967 : node2958;
									assign node2958 = (inp[5]) ? node2964 : node2959;
										assign node2959 = (inp[0]) ? 4'b0010 : node2960;
											assign node2960 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node2964 = (inp[7]) ? 4'b0010 : 4'b0110;
									assign node2967 = (inp[13]) ? node2977 : node2968;
										assign node2968 = (inp[11]) ? 4'b0111 : node2969;
											assign node2969 = (inp[10]) ? 4'b0110 : node2970;
												assign node2970 = (inp[2]) ? 4'b0011 : node2971;
													assign node2971 = (inp[5]) ? 4'b0110 : 4'b0010;
										assign node2977 = (inp[11]) ? 4'b0010 : node2978;
											assign node2978 = (inp[0]) ? node2980 : 4'b0111;
												assign node2980 = (inp[10]) ? 4'b0011 : 4'b0010;
								assign node2984 = (inp[2]) ? node3010 : node2985;
									assign node2985 = (inp[13]) ? node2999 : node2986;
										assign node2986 = (inp[11]) ? node2992 : node2987;
											assign node2987 = (inp[5]) ? 4'b0110 : node2988;
												assign node2988 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node2992 = (inp[5]) ? node2996 : node2993;
												assign node2993 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node2996 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node2999 = (inp[11]) ? node3007 : node3000;
											assign node3000 = (inp[0]) ? node3002 : 4'b0111;
												assign node3002 = (inp[7]) ? node3004 : 4'b0011;
													assign node3004 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node3007 = (inp[10]) ? 4'b0111 : 4'b0011;
									assign node3010 = (inp[11]) ? node3018 : node3011;
										assign node3011 = (inp[13]) ? node3015 : node3012;
											assign node3012 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node3015 = (inp[1]) ? 4'b0111 : 4'b0011;
										assign node3018 = (inp[13]) ? 4'b0010 : node3019;
											assign node3019 = (inp[4]) ? 4'b0010 : 4'b0011;
					assign node3023 = (inp[4]) ? node3133 : node3024;
						assign node3024 = (inp[3]) ? node3090 : node3025;
							assign node3025 = (inp[12]) ? node3053 : node3026;
								assign node3026 = (inp[7]) ? node3044 : node3027;
									assign node3027 = (inp[13]) ? node3037 : node3028;
										assign node3028 = (inp[1]) ? node3032 : node3029;
											assign node3029 = (inp[5]) ? 4'b0110 : 4'b0010;
											assign node3032 = (inp[0]) ? node3034 : 4'b0111;
												assign node3034 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node3037 = (inp[1]) ? node3039 : 4'b0011;
											assign node3039 = (inp[11]) ? 4'b0110 : node3040;
												assign node3040 = (inp[2]) ? 4'b0111 : 4'b0011;
									assign node3044 = (inp[11]) ? node3048 : node3045;
										assign node3045 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node3048 = (inp[0]) ? node3050 : 4'b0010;
											assign node3050 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node3053 = (inp[9]) ? node3077 : node3054;
									assign node3054 = (inp[11]) ? node3068 : node3055;
										assign node3055 = (inp[5]) ? node3061 : node3056;
											assign node3056 = (inp[1]) ? node3058 : 4'b0011;
												assign node3058 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node3061 = (inp[1]) ? 4'b0011 : node3062;
												assign node3062 = (inp[10]) ? node3064 : 4'b0111;
													assign node3064 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node3068 = (inp[10]) ? node3074 : node3069;
											assign node3069 = (inp[5]) ? 4'b0011 : node3070;
												assign node3070 = (inp[7]) ? 4'b0111 : 4'b0011;
											assign node3074 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node3077 = (inp[13]) ? 4'b0011 : node3078;
										assign node3078 = (inp[10]) ? node3080 : 4'b0010;
											assign node3080 = (inp[11]) ? 4'b0111 : node3081;
												assign node3081 = (inp[0]) ? 4'b0111 : node3082;
													assign node3082 = (inp[1]) ? 4'b0010 : node3083;
														assign node3083 = (inp[5]) ? 4'b0110 : 4'b0010;
							assign node3090 = (inp[12]) ? node3114 : node3091;
								assign node3091 = (inp[5]) ? node3109 : node3092;
									assign node3092 = (inp[7]) ? node3104 : node3093;
										assign node3093 = (inp[13]) ? node3099 : node3094;
											assign node3094 = (inp[1]) ? 4'b0001 : node3095;
												assign node3095 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node3099 = (inp[10]) ? node3101 : 4'b0000;
												assign node3101 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node3104 = (inp[2]) ? node3106 : 4'b0000;
											assign node3106 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node3109 = (inp[11]) ? 4'b0100 : node3110;
										assign node3110 = (inp[7]) ? 4'b0101 : 4'b0100;
								assign node3114 = (inp[5]) ? node3130 : node3115;
									assign node3115 = (inp[9]) ? node3117 : 4'b0101;
										assign node3117 = (inp[0]) ? node3123 : node3118;
											assign node3118 = (inp[7]) ? 4'b0101 : node3119;
												assign node3119 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node3123 = (inp[1]) ? node3125 : 4'b0101;
												assign node3125 = (inp[2]) ? node3127 : 4'b0100;
													assign node3127 = (inp[13]) ? 4'b0101 : 4'b0100;
									assign node3130 = (inp[0]) ? 4'b0001 : 4'b0000;
						assign node3133 = (inp[5]) ? node3205 : node3134;
							assign node3134 = (inp[3]) ? node3164 : node3135;
								assign node3135 = (inp[9]) ? node3157 : node3136;
									assign node3136 = (inp[1]) ? node3146 : node3137;
										assign node3137 = (inp[12]) ? 4'b0000 : node3138;
											assign node3138 = (inp[7]) ? node3142 : node3139;
												assign node3139 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node3142 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node3146 = (inp[7]) ? node3152 : node3147;
											assign node3147 = (inp[12]) ? 4'b0101 : node3148;
												assign node3148 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node3152 = (inp[0]) ? node3154 : 4'b0100;
												assign node3154 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node3157 = (inp[13]) ? node3161 : node3158;
										assign node3158 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node3161 = (inp[2]) ? 4'b0001 : 4'b0101;
								assign node3164 = (inp[2]) ? node3176 : node3165;
									assign node3165 = (inp[11]) ? node3171 : node3166;
										assign node3166 = (inp[1]) ? 4'b0101 : node3167;
											assign node3167 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node3171 = (inp[7]) ? node3173 : 4'b0101;
											assign node3173 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node3176 = (inp[10]) ? node3188 : node3177;
										assign node3177 = (inp[12]) ? node3179 : 4'b0100;
											assign node3179 = (inp[9]) ? node3185 : node3180;
												assign node3180 = (inp[11]) ? node3182 : 4'b0100;
													assign node3182 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node3185 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node3188 = (inp[13]) ? node3200 : node3189;
											assign node3189 = (inp[12]) ? node3191 : 4'b0101;
												assign node3191 = (inp[1]) ? 4'b0101 : node3192;
													assign node3192 = (inp[0]) ? node3194 : 4'b0100;
														assign node3194 = (inp[9]) ? node3196 : 4'b0101;
															assign node3196 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node3200 = (inp[0]) ? node3202 : 4'b0100;
												assign node3202 = (inp[1]) ? 4'b0100 : 4'b0101;
							assign node3205 = (inp[3]) ? node3243 : node3206;
								assign node3206 = (inp[1]) ? node3224 : node3207;
									assign node3207 = (inp[12]) ? node3211 : node3208;
										assign node3208 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node3211 = (inp[2]) ? node3221 : node3212;
											assign node3212 = (inp[0]) ? node3214 : 4'b0100;
												assign node3214 = (inp[7]) ? node3216 : 4'b0101;
													assign node3216 = (inp[11]) ? node3218 : 4'b0100;
														assign node3218 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node3221 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node3224 = (inp[7]) ? node3234 : node3225;
										assign node3225 = (inp[12]) ? node3231 : node3226;
											assign node3226 = (inp[11]) ? 4'b0100 : node3227;
												assign node3227 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node3231 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node3234 = (inp[12]) ? 4'b0001 : node3235;
											assign node3235 = (inp[0]) ? 4'b0000 : node3236;
												assign node3236 = (inp[10]) ? 4'b0001 : node3237;
													assign node3237 = (inp[13]) ? 4'b0001 : 4'b0000;
								assign node3243 = (inp[11]) ? node3249 : node3244;
									assign node3244 = (inp[12]) ? 4'b0001 : node3245;
										assign node3245 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node3249 = (inp[12]) ? 4'b0000 : node3250;
										assign node3250 = (inp[13]) ? node3256 : node3251;
											assign node3251 = (inp[9]) ? 4'b0001 : node3252;
												assign node3252 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node3256 = (inp[7]) ? 4'b0000 : node3257;
												assign node3257 = (inp[10]) ? 4'b0001 : 4'b0000;
			assign node3262 = (inp[3]) ? node3744 : node3263;
				assign node3263 = (inp[4]) ? node3543 : node3264;
					assign node3264 = (inp[8]) ? node3410 : node3265;
						assign node3265 = (inp[7]) ? node3331 : node3266;
							assign node3266 = (inp[2]) ? node3296 : node3267;
								assign node3267 = (inp[13]) ? node3281 : node3268;
									assign node3268 = (inp[9]) ? node3272 : node3269;
										assign node3269 = (inp[15]) ? 4'b0100 : 4'b0000;
										assign node3272 = (inp[10]) ? node3276 : node3273;
											assign node3273 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node3276 = (inp[1]) ? 4'b0100 : node3277;
												assign node3277 = (inp[12]) ? 4'b0101 : 4'b0001;
									assign node3281 = (inp[12]) ? node3291 : node3282;
										assign node3282 = (inp[15]) ? node3286 : node3283;
											assign node3283 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node3286 = (inp[11]) ? 4'b0001 : node3287;
												assign node3287 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node3291 = (inp[1]) ? 4'b0000 : node3292;
											assign node3292 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node3296 = (inp[13]) ? node3310 : node3297;
									assign node3297 = (inp[9]) ? node3303 : node3298;
										assign node3298 = (inp[15]) ? node3300 : 4'b0000;
											assign node3300 = (inp[11]) ? 4'b0100 : 4'b0000;
										assign node3303 = (inp[11]) ? 4'b0000 : node3304;
											assign node3304 = (inp[15]) ? 4'b0101 : node3305;
												assign node3305 = (inp[0]) ? 4'b0101 : 4'b0100;
									assign node3310 = (inp[1]) ? node3320 : node3311;
										assign node3311 = (inp[12]) ? 4'b0001 : node3312;
											assign node3312 = (inp[10]) ? 4'b0101 : node3313;
												assign node3313 = (inp[5]) ? 4'b0101 : node3314;
													assign node3314 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node3320 = (inp[11]) ? node3324 : node3321;
											assign node3321 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node3324 = (inp[0]) ? 4'b0101 : node3325;
												assign node3325 = (inp[12]) ? 4'b0100 : node3326;
													assign node3326 = (inp[5]) ? 4'b0000 : 4'b0001;
							assign node3331 = (inp[5]) ? node3361 : node3332;
								assign node3332 = (inp[11]) ? node3346 : node3333;
									assign node3333 = (inp[1]) ? node3339 : node3334;
										assign node3334 = (inp[2]) ? node3336 : 4'b0111;
											assign node3336 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node3339 = (inp[13]) ? node3343 : node3340;
											assign node3340 = (inp[15]) ? 4'b0010 : 4'b0011;
											assign node3343 = (inp[2]) ? 4'b0010 : 4'b0110;
									assign node3346 = (inp[12]) ? node3354 : node3347;
										assign node3347 = (inp[2]) ? 4'b0011 : node3348;
											assign node3348 = (inp[9]) ? node3350 : 4'b0011;
												assign node3350 = (inp[15]) ? 4'b0010 : 4'b0011;
										assign node3354 = (inp[0]) ? 4'b0111 : node3355;
											assign node3355 = (inp[13]) ? 4'b0010 : node3356;
												assign node3356 = (inp[15]) ? 4'b0010 : 4'b0110;
								assign node3361 = (inp[15]) ? node3385 : node3362;
									assign node3362 = (inp[11]) ? node3372 : node3363;
										assign node3363 = (inp[2]) ? node3365 : 4'b0011;
											assign node3365 = (inp[10]) ? node3369 : node3366;
												assign node3366 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node3369 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node3372 = (inp[2]) ? node3376 : node3373;
											assign node3373 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node3376 = (inp[9]) ? 4'b0111 : node3377;
												assign node3377 = (inp[0]) ? node3379 : 4'b0010;
													assign node3379 = (inp[12]) ? node3381 : 4'b0111;
														assign node3381 = (inp[1]) ? 4'b0011 : 4'b0010;
									assign node3385 = (inp[9]) ? node3395 : node3386;
										assign node3386 = (inp[0]) ? node3392 : node3387;
											assign node3387 = (inp[12]) ? 4'b0111 : node3388;
												assign node3388 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node3392 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node3395 = (inp[10]) ? node3399 : node3396;
											assign node3396 = (inp[0]) ? 4'b0110 : 4'b0010;
											assign node3399 = (inp[1]) ? node3405 : node3400;
												assign node3400 = (inp[0]) ? node3402 : 4'b0110;
													assign node3402 = (inp[13]) ? 4'b0111 : 4'b0010;
												assign node3405 = (inp[2]) ? node3407 : 4'b0111;
													assign node3407 = (inp[12]) ? 4'b0110 : 4'b0111;
						assign node3410 = (inp[7]) ? node3490 : node3411;
							assign node3411 = (inp[5]) ? node3461 : node3412;
								assign node3412 = (inp[2]) ? node3436 : node3413;
									assign node3413 = (inp[9]) ? node3425 : node3414;
										assign node3414 = (inp[11]) ? node3416 : 4'b0110;
											assign node3416 = (inp[13]) ? node3422 : node3417;
												assign node3417 = (inp[1]) ? 4'b0110 : node3418;
													assign node3418 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node3422 = (inp[15]) ? 4'b0010 : 4'b0111;
										assign node3425 = (inp[12]) ? node3431 : node3426;
											assign node3426 = (inp[0]) ? node3428 : 4'b0110;
												assign node3428 = (inp[1]) ? 4'b0111 : 4'b0011;
											assign node3431 = (inp[1]) ? 4'b0010 : node3432;
												assign node3432 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node3436 = (inp[13]) ? node3450 : node3437;
										assign node3437 = (inp[10]) ? node3439 : 4'b0011;
											assign node3439 = (inp[0]) ? 4'b0110 : node3440;
												assign node3440 = (inp[15]) ? node3442 : 4'b0111;
													assign node3442 = (inp[9]) ? 4'b0111 : node3443;
														assign node3443 = (inp[1]) ? 4'b0011 : node3444;
															assign node3444 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node3450 = (inp[15]) ? 4'b0010 : node3451;
											assign node3451 = (inp[10]) ? node3457 : node3452;
												assign node3452 = (inp[12]) ? 4'b0011 : node3453;
													assign node3453 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node3457 = (inp[11]) ? 4'b0010 : 4'b0110;
								assign node3461 = (inp[13]) ? node3481 : node3462;
									assign node3462 = (inp[1]) ? node3472 : node3463;
										assign node3463 = (inp[12]) ? node3465 : 4'b0010;
											assign node3465 = (inp[0]) ? node3469 : node3466;
												assign node3466 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node3469 = (inp[15]) ? 4'b0110 : 4'b0111;
										assign node3472 = (inp[12]) ? node3478 : node3473;
											assign node3473 = (inp[2]) ? node3475 : 4'b0111;
												assign node3475 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node3478 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node3481 = (inp[9]) ? node3485 : node3482;
										assign node3482 = (inp[11]) ? 4'b0111 : 4'b0011;
										assign node3485 = (inp[2]) ? node3487 : 4'b0011;
											assign node3487 = (inp[15]) ? 4'b0011 : 4'b0010;
							assign node3490 = (inp[12]) ? node3510 : node3491;
								assign node3491 = (inp[1]) ? node3503 : node3492;
									assign node3492 = (inp[0]) ? node3498 : node3493;
										assign node3493 = (inp[2]) ? 4'b0011 : node3494;
											assign node3494 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node3498 = (inp[15]) ? node3500 : 4'b0010;
											assign node3500 = (inp[13]) ? 4'b0010 : 4'b0011;
									assign node3503 = (inp[13]) ? 4'b0110 : node3504;
										assign node3504 = (inp[5]) ? 4'b0110 : node3505;
											assign node3505 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node3510 = (inp[1]) ? node3518 : node3511;
									assign node3511 = (inp[0]) ? 4'b0111 : node3512;
										assign node3512 = (inp[13]) ? 4'b0110 : node3513;
											assign node3513 = (inp[2]) ? 4'b0111 : 4'b0110;
									assign node3518 = (inp[9]) ? node3530 : node3519;
										assign node3519 = (inp[15]) ? 4'b0011 : node3520;
											assign node3520 = (inp[11]) ? 4'b0010 : node3521;
												assign node3521 = (inp[13]) ? 4'b0011 : node3522;
													assign node3522 = (inp[10]) ? node3524 : 4'b0010;
														assign node3524 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node3530 = (inp[13]) ? node3536 : node3531;
											assign node3531 = (inp[15]) ? 4'b0010 : node3532;
												assign node3532 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node3536 = (inp[10]) ? node3538 : 4'b0011;
												assign node3538 = (inp[0]) ? 4'b0010 : node3539;
													assign node3539 = (inp[2]) ? 4'b0011 : 4'b0010;
					assign node3543 = (inp[8]) ? node3669 : node3544;
						assign node3544 = (inp[7]) ? node3618 : node3545;
							assign node3545 = (inp[11]) ? node3573 : node3546;
								assign node3546 = (inp[1]) ? node3556 : node3547;
									assign node3547 = (inp[0]) ? 4'b0111 : node3548;
										assign node3548 = (inp[5]) ? node3552 : node3549;
											assign node3549 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node3552 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node3556 = (inp[10]) ? node3562 : node3557;
										assign node3557 = (inp[12]) ? node3559 : 4'b0011;
											assign node3559 = (inp[13]) ? 4'b0111 : 4'b0010;
										assign node3562 = (inp[13]) ? node3570 : node3563;
											assign node3563 = (inp[15]) ? node3565 : 4'b0010;
												assign node3565 = (inp[12]) ? 4'b0111 : node3566;
													assign node3566 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node3570 = (inp[15]) ? 4'b0010 : 4'b0110;
								assign node3573 = (inp[12]) ? node3595 : node3574;
									assign node3574 = (inp[5]) ? node3586 : node3575;
										assign node3575 = (inp[2]) ? node3581 : node3576;
											assign node3576 = (inp[15]) ? 4'b0010 : node3577;
												assign node3577 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node3581 = (inp[0]) ? 4'b0010 : node3582;
												assign node3582 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node3586 = (inp[10]) ? node3592 : node3587;
											assign node3587 = (inp[9]) ? node3589 : 4'b0111;
												assign node3589 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node3592 = (inp[2]) ? 4'b0010 : 4'b0110;
									assign node3595 = (inp[5]) ? node3603 : node3596;
										assign node3596 = (inp[1]) ? 4'b0110 : node3597;
											assign node3597 = (inp[0]) ? 4'b0111 : node3598;
												assign node3598 = (inp[9]) ? 4'b0111 : 4'b0110;
										assign node3603 = (inp[13]) ? node3611 : node3604;
											assign node3604 = (inp[15]) ? 4'b0111 : node3605;
												assign node3605 = (inp[0]) ? 4'b0011 : node3606;
													assign node3606 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node3611 = (inp[2]) ? node3613 : 4'b0010;
												assign node3613 = (inp[10]) ? node3615 : 4'b0011;
													assign node3615 = (inp[1]) ? 4'b0010 : 4'b0011;
							assign node3618 = (inp[2]) ? node3634 : node3619;
								assign node3619 = (inp[15]) ? node3627 : node3620;
									assign node3620 = (inp[12]) ? 4'b0101 : node3621;
										assign node3621 = (inp[10]) ? 4'b0001 : node3622;
											assign node3622 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node3627 = (inp[12]) ? 4'b0000 : node3628;
										assign node3628 = (inp[1]) ? 4'b0100 : node3629;
											assign node3629 = (inp[0]) ? 4'b0000 : 4'b0100;
								assign node3634 = (inp[1]) ? node3654 : node3635;
									assign node3635 = (inp[13]) ? node3643 : node3636;
										assign node3636 = (inp[10]) ? node3638 : 4'b0000;
											assign node3638 = (inp[0]) ? node3640 : 4'b0001;
												assign node3640 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node3643 = (inp[5]) ? node3649 : node3644;
											assign node3644 = (inp[9]) ? node3646 : 4'b0100;
												assign node3646 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node3649 = (inp[10]) ? node3651 : 4'b0101;
												assign node3651 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node3654 = (inp[13]) ? node3664 : node3655;
										assign node3655 = (inp[10]) ? 4'b0101 : node3656;
											assign node3656 = (inp[0]) ? 4'b0100 : node3657;
												assign node3657 = (inp[9]) ? node3659 : 4'b0101;
													assign node3659 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node3664 = (inp[12]) ? node3666 : 4'b0001;
											assign node3666 = (inp[9]) ? 4'b0000 : 4'b0001;
						assign node3669 = (inp[1]) ? node3711 : node3670;
							assign node3670 = (inp[15]) ? node3690 : node3671;
								assign node3671 = (inp[7]) ? node3683 : node3672;
									assign node3672 = (inp[13]) ? node3674 : 4'b0001;
										assign node3674 = (inp[5]) ? node3680 : node3675;
											assign node3675 = (inp[0]) ? node3677 : 4'b0001;
												assign node3677 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node3680 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node3683 = (inp[12]) ? node3687 : node3684;
										assign node3684 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node3687 = (inp[0]) ? 4'b0100 : 4'b0101;
								assign node3690 = (inp[10]) ? node3700 : node3691;
									assign node3691 = (inp[0]) ? 4'b0101 : node3692;
										assign node3692 = (inp[12]) ? 4'b0101 : node3693;
											assign node3693 = (inp[5]) ? 4'b0100 : node3694;
												assign node3694 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node3700 = (inp[7]) ? node3706 : node3701;
										assign node3701 = (inp[12]) ? 4'b0100 : node3702;
											assign node3702 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node3706 = (inp[0]) ? 4'b0100 : node3707;
											assign node3707 = (inp[12]) ? 4'b0101 : 4'b0100;
							assign node3711 = (inp[7]) ? node3733 : node3712;
								assign node3712 = (inp[15]) ? node3724 : node3713;
									assign node3713 = (inp[11]) ? node3719 : node3714;
										assign node3714 = (inp[9]) ? node3716 : 4'b0101;
											assign node3716 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node3719 = (inp[10]) ? node3721 : 4'b0100;
											assign node3721 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node3724 = (inp[12]) ? node3726 : 4'b0000;
										assign node3726 = (inp[13]) ? node3728 : 4'b0001;
											assign node3728 = (inp[10]) ? 4'b0000 : node3729;
												assign node3729 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node3733 = (inp[0]) ? node3739 : node3734;
									assign node3734 = (inp[13]) ? 4'b0001 : node3735;
										assign node3735 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node3739 = (inp[15]) ? 4'b0000 : node3740;
										assign node3740 = (inp[13]) ? 4'b0000 : 4'b0001;
				assign node3744 = (inp[8]) ? node3978 : node3745;
					assign node3745 = (inp[7]) ? node3877 : node3746;
						assign node3746 = (inp[13]) ? node3814 : node3747;
							assign node3747 = (inp[15]) ? node3795 : node3748;
								assign node3748 = (inp[4]) ? node3778 : node3749;
									assign node3749 = (inp[0]) ? node3765 : node3750;
										assign node3750 = (inp[10]) ? node3762 : node3751;
											assign node3751 = (inp[5]) ? node3757 : node3752;
												assign node3752 = (inp[2]) ? 4'b0110 : node3753;
													assign node3753 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node3757 = (inp[2]) ? 4'b0111 : node3758;
													assign node3758 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node3762 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node3765 = (inp[10]) ? node3773 : node3766;
											assign node3766 = (inp[5]) ? 4'b0110 : node3767;
												assign node3767 = (inp[12]) ? 4'b0010 : node3768;
													assign node3768 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node3773 = (inp[2]) ? node3775 : 4'b0011;
												assign node3775 = (inp[1]) ? 4'b0011 : 4'b0110;
									assign node3778 = (inp[1]) ? node3788 : node3779;
										assign node3779 = (inp[2]) ? node3781 : 4'b0011;
											assign node3781 = (inp[10]) ? 4'b0011 : node3782;
												assign node3782 = (inp[0]) ? node3784 : 4'b0010;
													assign node3784 = (inp[12]) ? 4'b0011 : 4'b0010;
										assign node3788 = (inp[5]) ? 4'b0010 : node3789;
											assign node3789 = (inp[12]) ? node3791 : 4'b0011;
												assign node3791 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node3795 = (inp[12]) ? node3801 : node3796;
									assign node3796 = (inp[4]) ? 4'b0111 : node3797;
										assign node3797 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node3801 = (inp[2]) ? 4'b0110 : node3802;
										assign node3802 = (inp[4]) ? node3804 : 4'b0110;
											assign node3804 = (inp[10]) ? node3808 : node3805;
												assign node3805 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node3808 = (inp[0]) ? 4'b0110 : node3809;
													assign node3809 = (inp[9]) ? 4'b0110 : 4'b0111;
							assign node3814 = (inp[12]) ? node3848 : node3815;
								assign node3815 = (inp[1]) ? node3829 : node3816;
									assign node3816 = (inp[4]) ? node3822 : node3817;
										assign node3817 = (inp[0]) ? 4'b0110 : node3818;
											assign node3818 = (inp[15]) ? 4'b0110 : 4'b0111;
										assign node3822 = (inp[15]) ? node3826 : node3823;
											assign node3823 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node3826 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node3829 = (inp[0]) ? node3833 : node3830;
										assign node3830 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node3833 = (inp[2]) ? 4'b0111 : node3834;
											assign node3834 = (inp[9]) ? node3842 : node3835;
												assign node3835 = (inp[5]) ? node3837 : 4'b0110;
													assign node3837 = (inp[15]) ? node3839 : 4'b0011;
														assign node3839 = (inp[10]) ? 4'b0011 : 4'b0110;
												assign node3842 = (inp[15]) ? 4'b0011 : node3843;
													assign node3843 = (inp[11]) ? 4'b0011 : 4'b0111;
								assign node3848 = (inp[15]) ? node3862 : node3849;
									assign node3849 = (inp[1]) ? 4'b0111 : node3850;
										assign node3850 = (inp[4]) ? 4'b0110 : node3851;
											assign node3851 = (inp[11]) ? 4'b0010 : node3852;
												assign node3852 = (inp[5]) ? 4'b0011 : node3853;
													assign node3853 = (inp[2]) ? 4'b0010 : node3854;
														assign node3854 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node3862 = (inp[10]) ? node3870 : node3863;
										assign node3863 = (inp[1]) ? node3865 : 4'b0011;
											assign node3865 = (inp[4]) ? node3867 : 4'b0010;
												assign node3867 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node3870 = (inp[4]) ? 4'b0010 : node3871;
											assign node3871 = (inp[0]) ? node3873 : 4'b0011;
												assign node3873 = (inp[9]) ? 4'b0011 : 4'b0010;
						assign node3877 = (inp[13]) ? node3923 : node3878;
							assign node3878 = (inp[4]) ? node3902 : node3879;
								assign node3879 = (inp[12]) ? node3891 : node3880;
									assign node3880 = (inp[15]) ? node3886 : node3881;
										assign node3881 = (inp[1]) ? 4'b0000 : node3882;
											assign node3882 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node3886 = (inp[10]) ? node3888 : 4'b0000;
											assign node3888 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node3891 = (inp[9]) ? node3897 : node3892;
										assign node3892 = (inp[2]) ? node3894 : 4'b0100;
											assign node3894 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node3897 = (inp[15]) ? node3899 : 4'b0001;
											assign node3899 = (inp[0]) ? 4'b0101 : 4'b0100;
								assign node3902 = (inp[1]) ? node3914 : node3903;
									assign node3903 = (inp[2]) ? 4'b0101 : node3904;
										assign node3904 = (inp[12]) ? node3908 : node3905;
											assign node3905 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node3908 = (inp[15]) ? node3910 : 4'b0101;
												assign node3910 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node3914 = (inp[2]) ? 4'b0100 : node3915;
										assign node3915 = (inp[11]) ? 4'b0101 : node3916;
											assign node3916 = (inp[12]) ? node3918 : 4'b0100;
												assign node3918 = (inp[9]) ? 4'b0100 : 4'b0101;
							assign node3923 = (inp[4]) ? node3955 : node3924;
								assign node3924 = (inp[9]) ? node3932 : node3925;
									assign node3925 = (inp[10]) ? node3929 : node3926;
										assign node3926 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node3929 = (inp[0]) ? 4'b0001 : 4'b0101;
									assign node3932 = (inp[5]) ? node3950 : node3933;
										assign node3933 = (inp[1]) ? node3947 : node3934;
											assign node3934 = (inp[10]) ? node3944 : node3935;
												assign node3935 = (inp[2]) ? 4'b0100 : node3936;
													assign node3936 = (inp[15]) ? node3940 : node3937;
														assign node3937 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node3940 = (inp[12]) ? 4'b0001 : 4'b0100;
												assign node3944 = (inp[0]) ? 4'b0100 : 4'b0001;
											assign node3947 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node3950 = (inp[0]) ? 4'b0101 : node3951;
											assign node3951 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node3955 = (inp[9]) ? node3963 : node3956;
									assign node3956 = (inp[10]) ? 4'b0001 : node3957;
										assign node3957 = (inp[0]) ? node3959 : 4'b0001;
											assign node3959 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node3963 = (inp[1]) ? 4'b0000 : node3964;
										assign node3964 = (inp[10]) ? node3970 : node3965;
											assign node3965 = (inp[5]) ? 4'b0001 : node3966;
												assign node3966 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node3970 = (inp[11]) ? node3972 : 4'b0000;
												assign node3972 = (inp[0]) ? 4'b0000 : node3973;
													assign node3973 = (inp[15]) ? 4'b0000 : 4'b0001;
					assign node3978 = (inp[12]) ? node4086 : node3979;
						assign node3979 = (inp[4]) ? node4051 : node3980;
							assign node3980 = (inp[7]) ? node4020 : node3981;
								assign node3981 = (inp[15]) ? node3997 : node3982;
									assign node3982 = (inp[10]) ? node3990 : node3983;
										assign node3983 = (inp[13]) ? node3985 : 4'b0001;
											assign node3985 = (inp[2]) ? node3987 : 4'b0001;
												assign node3987 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node3990 = (inp[13]) ? node3992 : 4'b0000;
											assign node3992 = (inp[2]) ? node3994 : 4'b0001;
												assign node3994 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node3997 = (inp[10]) ? node4003 : node3998;
										assign node3998 = (inp[5]) ? 4'b0101 : node3999;
											assign node3999 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node4003 = (inp[13]) ? node4017 : node4004;
											assign node4004 = (inp[0]) ? node4012 : node4005;
												assign node4005 = (inp[11]) ? node4009 : node4006;
													assign node4006 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node4009 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node4012 = (inp[1]) ? node4014 : 4'b0100;
													assign node4014 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node4017 = (inp[1]) ? 4'b0100 : 4'b0101;
								assign node4020 = (inp[13]) ? node4032 : node4021;
									assign node4021 = (inp[2]) ? node4023 : 4'b0100;
										assign node4023 = (inp[15]) ? node4029 : node4024;
											assign node4024 = (inp[1]) ? 4'b0101 : node4025;
												assign node4025 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node4029 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node4032 = (inp[0]) ? node4046 : node4033;
										assign node4033 = (inp[11]) ? node4035 : 4'b0100;
											assign node4035 = (inp[15]) ? node4041 : node4036;
												assign node4036 = (inp[2]) ? 4'b0101 : node4037;
													assign node4037 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node4041 = (inp[10]) ? node4043 : 4'b0100;
													assign node4043 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node4046 = (inp[1]) ? node4048 : 4'b0101;
											assign node4048 = (inp[2]) ? 4'b0100 : 4'b0101;
							assign node4051 = (inp[7]) ? node4073 : node4052;
								assign node4052 = (inp[15]) ? node4060 : node4053;
									assign node4053 = (inp[5]) ? node4057 : node4054;
										assign node4054 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node4057 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node4060 = (inp[2]) ? node4064 : node4061;
										assign node4061 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node4064 = (inp[9]) ? 4'b0001 : node4065;
											assign node4065 = (inp[11]) ? 4'b0000 : node4066;
												assign node4066 = (inp[5]) ? node4068 : 4'b0001;
													assign node4068 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node4073 = (inp[1]) ? node4081 : node4074;
									assign node4074 = (inp[0]) ? node4076 : 4'b0001;
										assign node4076 = (inp[13]) ? 4'b0001 : node4077;
											assign node4077 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node4081 = (inp[13]) ? 4'b0000 : node4082;
										assign node4082 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node4086 = (inp[15]) ? node4134 : node4087;
							assign node4087 = (inp[7]) ? node4113 : node4088;
								assign node4088 = (inp[2]) ? node4106 : node4089;
									assign node4089 = (inp[11]) ? 4'b0100 : node4090;
										assign node4090 = (inp[4]) ? node4098 : node4091;
											assign node4091 = (inp[13]) ? node4093 : 4'b0100;
												assign node4093 = (inp[9]) ? node4095 : 4'b0101;
													assign node4095 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node4098 = (inp[10]) ? 4'b0101 : node4099;
												assign node4099 = (inp[13]) ? 4'b0100 : node4100;
													assign node4100 = (inp[5]) ? 4'b0101 : 4'b0100;
									assign node4106 = (inp[4]) ? node4108 : 4'b0101;
										assign node4108 = (inp[5]) ? 4'b0100 : node4109;
											assign node4109 = (inp[13]) ? 4'b0101 : 4'b0100;
								assign node4113 = (inp[13]) ? node4123 : node4114;
									assign node4114 = (inp[0]) ? node4120 : node4115;
										assign node4115 = (inp[11]) ? node4117 : 4'b0001;
											assign node4117 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node4120 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node4123 = (inp[4]) ? 4'b0000 : node4124;
										assign node4124 = (inp[11]) ? 4'b0001 : node4125;
											assign node4125 = (inp[1]) ? node4129 : node4126;
												assign node4126 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node4129 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node4134 = (inp[5]) ? node4150 : node4135;
								assign node4135 = (inp[9]) ? node4141 : node4136;
									assign node4136 = (inp[7]) ? node4138 : 4'b0001;
										assign node4138 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node4141 = (inp[0]) ? 4'b0000 : node4142;
										assign node4142 = (inp[13]) ? 4'b0001 : node4143;
											assign node4143 = (inp[7]) ? 4'b0000 : node4144;
												assign node4144 = (inp[2]) ? 4'b0001 : 4'b0000;
								assign node4150 = (inp[4]) ? 4'b0000 : node4151;
									assign node4151 = (inp[2]) ? 4'b0000 : 4'b0001;

endmodule