module dtc_split75_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node12;
	wire [16-1:0] node15;
	wire [16-1:0] node16;
	wire [16-1:0] node19;
	wire [16-1:0] node22;
	wire [16-1:0] node23;
	wire [16-1:0] node24;
	wire [16-1:0] node27;
	wire [16-1:0] node30;
	wire [16-1:0] node31;
	wire [16-1:0] node34;
	wire [16-1:0] node37;
	wire [16-1:0] node38;
	wire [16-1:0] node39;
	wire [16-1:0] node40;
	wire [16-1:0] node43;
	wire [16-1:0] node46;
	wire [16-1:0] node47;
	wire [16-1:0] node50;
	wire [16-1:0] node53;
	wire [16-1:0] node54;
	wire [16-1:0] node55;
	wire [16-1:0] node58;
	wire [16-1:0] node61;
	wire [16-1:0] node62;
	wire [16-1:0] node65;
	wire [16-1:0] node68;
	wire [16-1:0] node69;
	wire [16-1:0] node70;
	wire [16-1:0] node71;
	wire [16-1:0] node72;
	wire [16-1:0] node75;
	wire [16-1:0] node78;
	wire [16-1:0] node79;
	wire [16-1:0] node82;
	wire [16-1:0] node85;
	wire [16-1:0] node86;
	wire [16-1:0] node87;
	wire [16-1:0] node90;
	wire [16-1:0] node93;
	wire [16-1:0] node94;
	wire [16-1:0] node97;
	wire [16-1:0] node100;
	wire [16-1:0] node101;
	wire [16-1:0] node102;
	wire [16-1:0] node103;
	wire [16-1:0] node106;
	wire [16-1:0] node109;
	wire [16-1:0] node110;
	wire [16-1:0] node113;
	wire [16-1:0] node116;
	wire [16-1:0] node117;
	wire [16-1:0] node118;
	wire [16-1:0] node121;
	wire [16-1:0] node124;
	wire [16-1:0] node125;
	wire [16-1:0] node128;
	wire [16-1:0] node131;
	wire [16-1:0] node132;
	wire [16-1:0] node133;
	wire [16-1:0] node134;
	wire [16-1:0] node135;
	wire [16-1:0] node136;
	wire [16-1:0] node139;
	wire [16-1:0] node142;
	wire [16-1:0] node143;
	wire [16-1:0] node146;
	wire [16-1:0] node149;
	wire [16-1:0] node150;
	wire [16-1:0] node151;
	wire [16-1:0] node154;
	wire [16-1:0] node157;
	wire [16-1:0] node158;
	wire [16-1:0] node161;
	wire [16-1:0] node164;
	wire [16-1:0] node165;
	wire [16-1:0] node166;
	wire [16-1:0] node167;
	wire [16-1:0] node170;
	wire [16-1:0] node173;
	wire [16-1:0] node174;
	wire [16-1:0] node177;
	wire [16-1:0] node180;
	wire [16-1:0] node181;
	wire [16-1:0] node182;
	wire [16-1:0] node185;
	wire [16-1:0] node188;
	wire [16-1:0] node189;
	wire [16-1:0] node192;
	wire [16-1:0] node195;
	wire [16-1:0] node196;
	wire [16-1:0] node197;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node202;
	wire [16-1:0] node205;
	wire [16-1:0] node206;
	wire [16-1:0] node209;
	wire [16-1:0] node212;
	wire [16-1:0] node213;
	wire [16-1:0] node214;
	wire [16-1:0] node217;
	wire [16-1:0] node220;
	wire [16-1:0] node221;
	wire [16-1:0] node224;
	wire [16-1:0] node227;
	wire [16-1:0] node228;
	wire [16-1:0] node229;
	wire [16-1:0] node230;
	wire [16-1:0] node233;
	wire [16-1:0] node236;
	wire [16-1:0] node237;
	wire [16-1:0] node240;
	wire [16-1:0] node243;
	wire [16-1:0] node244;
	wire [16-1:0] node245;
	wire [16-1:0] node248;
	wire [16-1:0] node251;
	wire [16-1:0] node252;
	wire [16-1:0] node255;
	wire [16-1:0] node258;
	wire [16-1:0] node259;
	wire [16-1:0] node260;
	wire [16-1:0] node261;
	wire [16-1:0] node262;
	wire [16-1:0] node263;
	wire [16-1:0] node264;
	wire [16-1:0] node267;
	wire [16-1:0] node270;
	wire [16-1:0] node271;
	wire [16-1:0] node274;
	wire [16-1:0] node277;
	wire [16-1:0] node278;
	wire [16-1:0] node279;
	wire [16-1:0] node282;
	wire [16-1:0] node285;
	wire [16-1:0] node286;
	wire [16-1:0] node289;
	wire [16-1:0] node292;
	wire [16-1:0] node293;
	wire [16-1:0] node294;
	wire [16-1:0] node295;
	wire [16-1:0] node298;
	wire [16-1:0] node301;
	wire [16-1:0] node302;
	wire [16-1:0] node305;
	wire [16-1:0] node308;
	wire [16-1:0] node309;
	wire [16-1:0] node310;
	wire [16-1:0] node313;
	wire [16-1:0] node316;
	wire [16-1:0] node317;
	wire [16-1:0] node320;
	wire [16-1:0] node323;
	wire [16-1:0] node324;
	wire [16-1:0] node325;
	wire [16-1:0] node326;
	wire [16-1:0] node327;
	wire [16-1:0] node330;
	wire [16-1:0] node333;
	wire [16-1:0] node334;
	wire [16-1:0] node337;
	wire [16-1:0] node340;
	wire [16-1:0] node341;
	wire [16-1:0] node342;
	wire [16-1:0] node345;
	wire [16-1:0] node348;
	wire [16-1:0] node349;
	wire [16-1:0] node352;
	wire [16-1:0] node355;
	wire [16-1:0] node356;
	wire [16-1:0] node357;
	wire [16-1:0] node358;
	wire [16-1:0] node361;
	wire [16-1:0] node364;
	wire [16-1:0] node365;
	wire [16-1:0] node368;
	wire [16-1:0] node371;
	wire [16-1:0] node372;
	wire [16-1:0] node373;
	wire [16-1:0] node376;
	wire [16-1:0] node379;
	wire [16-1:0] node380;
	wire [16-1:0] node383;
	wire [16-1:0] node386;
	wire [16-1:0] node387;
	wire [16-1:0] node388;
	wire [16-1:0] node389;
	wire [16-1:0] node390;
	wire [16-1:0] node391;
	wire [16-1:0] node394;
	wire [16-1:0] node397;
	wire [16-1:0] node398;
	wire [16-1:0] node401;
	wire [16-1:0] node404;
	wire [16-1:0] node405;
	wire [16-1:0] node406;
	wire [16-1:0] node409;
	wire [16-1:0] node412;
	wire [16-1:0] node413;
	wire [16-1:0] node416;
	wire [16-1:0] node419;
	wire [16-1:0] node420;
	wire [16-1:0] node421;
	wire [16-1:0] node422;
	wire [16-1:0] node425;
	wire [16-1:0] node428;
	wire [16-1:0] node429;
	wire [16-1:0] node432;
	wire [16-1:0] node435;
	wire [16-1:0] node436;
	wire [16-1:0] node437;
	wire [16-1:0] node440;
	wire [16-1:0] node443;
	wire [16-1:0] node444;
	wire [16-1:0] node447;
	wire [16-1:0] node450;
	wire [16-1:0] node451;
	wire [16-1:0] node452;
	wire [16-1:0] node453;
	wire [16-1:0] node454;
	wire [16-1:0] node457;
	wire [16-1:0] node460;
	wire [16-1:0] node461;
	wire [16-1:0] node464;
	wire [16-1:0] node467;
	wire [16-1:0] node468;
	wire [16-1:0] node469;
	wire [16-1:0] node472;
	wire [16-1:0] node475;
	wire [16-1:0] node476;
	wire [16-1:0] node479;
	wire [16-1:0] node482;
	wire [16-1:0] node483;
	wire [16-1:0] node484;
	wire [16-1:0] node485;
	wire [16-1:0] node488;
	wire [16-1:0] node491;
	wire [16-1:0] node492;
	wire [16-1:0] node495;
	wire [16-1:0] node498;
	wire [16-1:0] node499;
	wire [16-1:0] node500;
	wire [16-1:0] node503;
	wire [16-1:0] node506;
	wire [16-1:0] node507;
	wire [16-1:0] node510;
	wire [16-1:0] node513;
	wire [16-1:0] node514;
	wire [16-1:0] node515;
	wire [16-1:0] node516;
	wire [16-1:0] node517;
	wire [16-1:0] node518;
	wire [16-1:0] node519;
	wire [16-1:0] node520;
	wire [16-1:0] node523;
	wire [16-1:0] node526;
	wire [16-1:0] node527;
	wire [16-1:0] node530;
	wire [16-1:0] node533;
	wire [16-1:0] node534;
	wire [16-1:0] node535;
	wire [16-1:0] node538;
	wire [16-1:0] node541;
	wire [16-1:0] node542;
	wire [16-1:0] node545;
	wire [16-1:0] node548;
	wire [16-1:0] node549;
	wire [16-1:0] node550;
	wire [16-1:0] node551;
	wire [16-1:0] node554;
	wire [16-1:0] node557;
	wire [16-1:0] node558;
	wire [16-1:0] node561;
	wire [16-1:0] node564;
	wire [16-1:0] node565;
	wire [16-1:0] node566;
	wire [16-1:0] node569;
	wire [16-1:0] node572;
	wire [16-1:0] node573;
	wire [16-1:0] node576;
	wire [16-1:0] node579;
	wire [16-1:0] node580;
	wire [16-1:0] node581;
	wire [16-1:0] node582;
	wire [16-1:0] node583;
	wire [16-1:0] node586;
	wire [16-1:0] node589;
	wire [16-1:0] node590;
	wire [16-1:0] node593;
	wire [16-1:0] node596;
	wire [16-1:0] node597;
	wire [16-1:0] node598;
	wire [16-1:0] node601;
	wire [16-1:0] node604;
	wire [16-1:0] node605;
	wire [16-1:0] node608;
	wire [16-1:0] node611;
	wire [16-1:0] node612;
	wire [16-1:0] node613;
	wire [16-1:0] node614;
	wire [16-1:0] node617;
	wire [16-1:0] node620;
	wire [16-1:0] node621;
	wire [16-1:0] node624;
	wire [16-1:0] node627;
	wire [16-1:0] node628;
	wire [16-1:0] node629;
	wire [16-1:0] node632;
	wire [16-1:0] node635;
	wire [16-1:0] node636;
	wire [16-1:0] node639;
	wire [16-1:0] node642;
	wire [16-1:0] node643;
	wire [16-1:0] node644;
	wire [16-1:0] node645;
	wire [16-1:0] node646;
	wire [16-1:0] node647;
	wire [16-1:0] node650;
	wire [16-1:0] node653;
	wire [16-1:0] node654;
	wire [16-1:0] node657;
	wire [16-1:0] node660;
	wire [16-1:0] node661;
	wire [16-1:0] node662;
	wire [16-1:0] node665;
	wire [16-1:0] node668;
	wire [16-1:0] node669;
	wire [16-1:0] node672;
	wire [16-1:0] node675;
	wire [16-1:0] node676;
	wire [16-1:0] node677;
	wire [16-1:0] node678;
	wire [16-1:0] node681;
	wire [16-1:0] node684;
	wire [16-1:0] node685;
	wire [16-1:0] node688;
	wire [16-1:0] node691;
	wire [16-1:0] node692;
	wire [16-1:0] node693;
	wire [16-1:0] node696;
	wire [16-1:0] node699;
	wire [16-1:0] node700;
	wire [16-1:0] node703;
	wire [16-1:0] node706;
	wire [16-1:0] node707;
	wire [16-1:0] node708;
	wire [16-1:0] node709;
	wire [16-1:0] node710;
	wire [16-1:0] node713;
	wire [16-1:0] node716;
	wire [16-1:0] node717;
	wire [16-1:0] node720;
	wire [16-1:0] node723;
	wire [16-1:0] node724;
	wire [16-1:0] node725;
	wire [16-1:0] node728;
	wire [16-1:0] node731;
	wire [16-1:0] node732;
	wire [16-1:0] node735;
	wire [16-1:0] node738;
	wire [16-1:0] node739;
	wire [16-1:0] node740;
	wire [16-1:0] node741;
	wire [16-1:0] node744;
	wire [16-1:0] node747;
	wire [16-1:0] node748;
	wire [16-1:0] node751;
	wire [16-1:0] node754;
	wire [16-1:0] node755;
	wire [16-1:0] node756;
	wire [16-1:0] node759;
	wire [16-1:0] node762;
	wire [16-1:0] node763;
	wire [16-1:0] node766;
	wire [16-1:0] node769;
	wire [16-1:0] node770;
	wire [16-1:0] node771;
	wire [16-1:0] node772;
	wire [16-1:0] node773;
	wire [16-1:0] node774;
	wire [16-1:0] node775;
	wire [16-1:0] node778;
	wire [16-1:0] node781;
	wire [16-1:0] node782;
	wire [16-1:0] node785;
	wire [16-1:0] node788;
	wire [16-1:0] node789;
	wire [16-1:0] node790;
	wire [16-1:0] node793;
	wire [16-1:0] node796;
	wire [16-1:0] node797;
	wire [16-1:0] node800;
	wire [16-1:0] node803;
	wire [16-1:0] node804;
	wire [16-1:0] node805;
	wire [16-1:0] node806;
	wire [16-1:0] node809;
	wire [16-1:0] node812;
	wire [16-1:0] node813;
	wire [16-1:0] node816;
	wire [16-1:0] node819;
	wire [16-1:0] node820;
	wire [16-1:0] node821;
	wire [16-1:0] node824;
	wire [16-1:0] node827;
	wire [16-1:0] node828;
	wire [16-1:0] node831;
	wire [16-1:0] node834;
	wire [16-1:0] node835;
	wire [16-1:0] node836;
	wire [16-1:0] node837;
	wire [16-1:0] node838;
	wire [16-1:0] node841;
	wire [16-1:0] node844;
	wire [16-1:0] node845;
	wire [16-1:0] node848;
	wire [16-1:0] node851;
	wire [16-1:0] node852;
	wire [16-1:0] node853;
	wire [16-1:0] node856;
	wire [16-1:0] node859;
	wire [16-1:0] node860;
	wire [16-1:0] node863;
	wire [16-1:0] node866;
	wire [16-1:0] node867;
	wire [16-1:0] node868;
	wire [16-1:0] node869;
	wire [16-1:0] node872;
	wire [16-1:0] node875;
	wire [16-1:0] node876;
	wire [16-1:0] node879;
	wire [16-1:0] node882;
	wire [16-1:0] node883;
	wire [16-1:0] node884;
	wire [16-1:0] node887;
	wire [16-1:0] node890;
	wire [16-1:0] node891;
	wire [16-1:0] node894;
	wire [16-1:0] node897;
	wire [16-1:0] node898;
	wire [16-1:0] node899;
	wire [16-1:0] node900;
	wire [16-1:0] node901;
	wire [16-1:0] node902;
	wire [16-1:0] node905;
	wire [16-1:0] node908;
	wire [16-1:0] node909;
	wire [16-1:0] node912;
	wire [16-1:0] node915;
	wire [16-1:0] node916;
	wire [16-1:0] node917;
	wire [16-1:0] node920;
	wire [16-1:0] node923;
	wire [16-1:0] node924;
	wire [16-1:0] node927;
	wire [16-1:0] node930;
	wire [16-1:0] node931;
	wire [16-1:0] node932;
	wire [16-1:0] node933;
	wire [16-1:0] node936;
	wire [16-1:0] node939;
	wire [16-1:0] node940;
	wire [16-1:0] node943;
	wire [16-1:0] node946;
	wire [16-1:0] node947;
	wire [16-1:0] node948;
	wire [16-1:0] node951;
	wire [16-1:0] node954;
	wire [16-1:0] node955;
	wire [16-1:0] node958;
	wire [16-1:0] node961;
	wire [16-1:0] node962;
	wire [16-1:0] node963;
	wire [16-1:0] node964;
	wire [16-1:0] node965;
	wire [16-1:0] node968;
	wire [16-1:0] node971;
	wire [16-1:0] node972;
	wire [16-1:0] node975;
	wire [16-1:0] node978;
	wire [16-1:0] node979;
	wire [16-1:0] node980;
	wire [16-1:0] node983;
	wire [16-1:0] node986;
	wire [16-1:0] node987;
	wire [16-1:0] node990;
	wire [16-1:0] node993;
	wire [16-1:0] node994;
	wire [16-1:0] node995;
	wire [16-1:0] node996;
	wire [16-1:0] node999;
	wire [16-1:0] node1002;
	wire [16-1:0] node1003;
	wire [16-1:0] node1006;
	wire [16-1:0] node1009;
	wire [16-1:0] node1010;
	wire [16-1:0] node1011;
	wire [16-1:0] node1014;
	wire [16-1:0] node1017;
	wire [16-1:0] node1018;
	wire [16-1:0] node1021;
	wire [16-1:0] node1024;
	wire [16-1:0] node1025;
	wire [16-1:0] node1026;
	wire [16-1:0] node1027;
	wire [16-1:0] node1028;
	wire [16-1:0] node1029;
	wire [16-1:0] node1030;
	wire [16-1:0] node1031;
	wire [16-1:0] node1032;
	wire [16-1:0] node1035;
	wire [16-1:0] node1038;
	wire [16-1:0] node1039;
	wire [16-1:0] node1042;
	wire [16-1:0] node1045;
	wire [16-1:0] node1046;
	wire [16-1:0] node1047;
	wire [16-1:0] node1050;
	wire [16-1:0] node1053;
	wire [16-1:0] node1054;
	wire [16-1:0] node1057;
	wire [16-1:0] node1060;
	wire [16-1:0] node1061;
	wire [16-1:0] node1062;
	wire [16-1:0] node1063;
	wire [16-1:0] node1066;
	wire [16-1:0] node1069;
	wire [16-1:0] node1070;
	wire [16-1:0] node1073;
	wire [16-1:0] node1076;
	wire [16-1:0] node1077;
	wire [16-1:0] node1078;
	wire [16-1:0] node1081;
	wire [16-1:0] node1084;
	wire [16-1:0] node1085;
	wire [16-1:0] node1088;
	wire [16-1:0] node1091;
	wire [16-1:0] node1092;
	wire [16-1:0] node1093;
	wire [16-1:0] node1094;
	wire [16-1:0] node1095;
	wire [16-1:0] node1098;
	wire [16-1:0] node1101;
	wire [16-1:0] node1102;
	wire [16-1:0] node1105;
	wire [16-1:0] node1108;
	wire [16-1:0] node1109;
	wire [16-1:0] node1110;
	wire [16-1:0] node1113;
	wire [16-1:0] node1116;
	wire [16-1:0] node1117;
	wire [16-1:0] node1120;
	wire [16-1:0] node1123;
	wire [16-1:0] node1124;
	wire [16-1:0] node1125;
	wire [16-1:0] node1126;
	wire [16-1:0] node1129;
	wire [16-1:0] node1132;
	wire [16-1:0] node1133;
	wire [16-1:0] node1136;
	wire [16-1:0] node1139;
	wire [16-1:0] node1140;
	wire [16-1:0] node1141;
	wire [16-1:0] node1144;
	wire [16-1:0] node1147;
	wire [16-1:0] node1148;
	wire [16-1:0] node1151;
	wire [16-1:0] node1154;
	wire [16-1:0] node1155;
	wire [16-1:0] node1156;
	wire [16-1:0] node1157;
	wire [16-1:0] node1158;
	wire [16-1:0] node1159;
	wire [16-1:0] node1162;
	wire [16-1:0] node1165;
	wire [16-1:0] node1166;
	wire [16-1:0] node1169;
	wire [16-1:0] node1172;
	wire [16-1:0] node1173;
	wire [16-1:0] node1174;
	wire [16-1:0] node1177;
	wire [16-1:0] node1180;
	wire [16-1:0] node1181;
	wire [16-1:0] node1184;
	wire [16-1:0] node1187;
	wire [16-1:0] node1188;
	wire [16-1:0] node1189;
	wire [16-1:0] node1190;
	wire [16-1:0] node1193;
	wire [16-1:0] node1196;
	wire [16-1:0] node1197;
	wire [16-1:0] node1200;
	wire [16-1:0] node1203;
	wire [16-1:0] node1204;
	wire [16-1:0] node1205;
	wire [16-1:0] node1208;
	wire [16-1:0] node1211;
	wire [16-1:0] node1212;
	wire [16-1:0] node1215;
	wire [16-1:0] node1218;
	wire [16-1:0] node1219;
	wire [16-1:0] node1220;
	wire [16-1:0] node1221;
	wire [16-1:0] node1222;
	wire [16-1:0] node1225;
	wire [16-1:0] node1228;
	wire [16-1:0] node1229;
	wire [16-1:0] node1232;
	wire [16-1:0] node1235;
	wire [16-1:0] node1236;
	wire [16-1:0] node1237;
	wire [16-1:0] node1240;
	wire [16-1:0] node1243;
	wire [16-1:0] node1244;
	wire [16-1:0] node1247;
	wire [16-1:0] node1250;
	wire [16-1:0] node1251;
	wire [16-1:0] node1252;
	wire [16-1:0] node1253;
	wire [16-1:0] node1256;
	wire [16-1:0] node1259;
	wire [16-1:0] node1260;
	wire [16-1:0] node1263;
	wire [16-1:0] node1266;
	wire [16-1:0] node1267;
	wire [16-1:0] node1268;
	wire [16-1:0] node1271;
	wire [16-1:0] node1274;
	wire [16-1:0] node1275;
	wire [16-1:0] node1278;
	wire [16-1:0] node1281;
	wire [16-1:0] node1282;
	wire [16-1:0] node1283;
	wire [16-1:0] node1284;
	wire [16-1:0] node1285;
	wire [16-1:0] node1286;
	wire [16-1:0] node1287;
	wire [16-1:0] node1290;
	wire [16-1:0] node1293;
	wire [16-1:0] node1294;
	wire [16-1:0] node1297;
	wire [16-1:0] node1300;
	wire [16-1:0] node1301;
	wire [16-1:0] node1302;
	wire [16-1:0] node1305;
	wire [16-1:0] node1308;
	wire [16-1:0] node1309;
	wire [16-1:0] node1312;
	wire [16-1:0] node1315;
	wire [16-1:0] node1316;
	wire [16-1:0] node1317;
	wire [16-1:0] node1318;
	wire [16-1:0] node1321;
	wire [16-1:0] node1324;
	wire [16-1:0] node1325;
	wire [16-1:0] node1328;
	wire [16-1:0] node1331;
	wire [16-1:0] node1332;
	wire [16-1:0] node1333;
	wire [16-1:0] node1336;
	wire [16-1:0] node1339;
	wire [16-1:0] node1340;
	wire [16-1:0] node1343;
	wire [16-1:0] node1346;
	wire [16-1:0] node1347;
	wire [16-1:0] node1348;
	wire [16-1:0] node1349;
	wire [16-1:0] node1350;
	wire [16-1:0] node1353;
	wire [16-1:0] node1356;
	wire [16-1:0] node1357;
	wire [16-1:0] node1360;
	wire [16-1:0] node1363;
	wire [16-1:0] node1364;
	wire [16-1:0] node1365;
	wire [16-1:0] node1368;
	wire [16-1:0] node1371;
	wire [16-1:0] node1372;
	wire [16-1:0] node1375;
	wire [16-1:0] node1378;
	wire [16-1:0] node1379;
	wire [16-1:0] node1380;
	wire [16-1:0] node1381;
	wire [16-1:0] node1384;
	wire [16-1:0] node1387;
	wire [16-1:0] node1388;
	wire [16-1:0] node1391;
	wire [16-1:0] node1394;
	wire [16-1:0] node1395;
	wire [16-1:0] node1396;
	wire [16-1:0] node1399;
	wire [16-1:0] node1402;
	wire [16-1:0] node1403;
	wire [16-1:0] node1406;
	wire [16-1:0] node1409;
	wire [16-1:0] node1410;
	wire [16-1:0] node1411;
	wire [16-1:0] node1412;
	wire [16-1:0] node1413;
	wire [16-1:0] node1414;
	wire [16-1:0] node1417;
	wire [16-1:0] node1420;
	wire [16-1:0] node1421;
	wire [16-1:0] node1424;
	wire [16-1:0] node1427;
	wire [16-1:0] node1428;
	wire [16-1:0] node1429;
	wire [16-1:0] node1432;
	wire [16-1:0] node1435;
	wire [16-1:0] node1436;
	wire [16-1:0] node1439;
	wire [16-1:0] node1442;
	wire [16-1:0] node1443;
	wire [16-1:0] node1444;
	wire [16-1:0] node1445;
	wire [16-1:0] node1448;
	wire [16-1:0] node1451;
	wire [16-1:0] node1452;
	wire [16-1:0] node1455;
	wire [16-1:0] node1458;
	wire [16-1:0] node1459;
	wire [16-1:0] node1460;
	wire [16-1:0] node1463;
	wire [16-1:0] node1466;
	wire [16-1:0] node1467;
	wire [16-1:0] node1470;
	wire [16-1:0] node1473;
	wire [16-1:0] node1474;
	wire [16-1:0] node1475;
	wire [16-1:0] node1476;
	wire [16-1:0] node1477;
	wire [16-1:0] node1480;
	wire [16-1:0] node1483;
	wire [16-1:0] node1484;
	wire [16-1:0] node1487;
	wire [16-1:0] node1490;
	wire [16-1:0] node1491;
	wire [16-1:0] node1492;
	wire [16-1:0] node1495;
	wire [16-1:0] node1498;
	wire [16-1:0] node1499;
	wire [16-1:0] node1502;
	wire [16-1:0] node1505;
	wire [16-1:0] node1506;
	wire [16-1:0] node1507;
	wire [16-1:0] node1508;
	wire [16-1:0] node1511;
	wire [16-1:0] node1514;
	wire [16-1:0] node1515;
	wire [16-1:0] node1518;
	wire [16-1:0] node1521;
	wire [16-1:0] node1522;
	wire [16-1:0] node1523;
	wire [16-1:0] node1526;
	wire [16-1:0] node1529;
	wire [16-1:0] node1530;
	wire [16-1:0] node1533;
	wire [16-1:0] node1536;
	wire [16-1:0] node1537;
	wire [16-1:0] node1538;
	wire [16-1:0] node1539;
	wire [16-1:0] node1540;
	wire [16-1:0] node1541;
	wire [16-1:0] node1542;
	wire [16-1:0] node1543;
	wire [16-1:0] node1546;
	wire [16-1:0] node1549;
	wire [16-1:0] node1550;
	wire [16-1:0] node1553;
	wire [16-1:0] node1556;
	wire [16-1:0] node1557;
	wire [16-1:0] node1558;
	wire [16-1:0] node1561;
	wire [16-1:0] node1564;
	wire [16-1:0] node1565;
	wire [16-1:0] node1568;
	wire [16-1:0] node1571;
	wire [16-1:0] node1572;
	wire [16-1:0] node1573;
	wire [16-1:0] node1574;
	wire [16-1:0] node1577;
	wire [16-1:0] node1580;
	wire [16-1:0] node1581;
	wire [16-1:0] node1584;
	wire [16-1:0] node1587;
	wire [16-1:0] node1588;
	wire [16-1:0] node1589;
	wire [16-1:0] node1592;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1599;
	wire [16-1:0] node1602;
	wire [16-1:0] node1603;
	wire [16-1:0] node1604;
	wire [16-1:0] node1605;
	wire [16-1:0] node1606;
	wire [16-1:0] node1609;
	wire [16-1:0] node1612;
	wire [16-1:0] node1613;
	wire [16-1:0] node1616;
	wire [16-1:0] node1619;
	wire [16-1:0] node1620;
	wire [16-1:0] node1621;
	wire [16-1:0] node1624;
	wire [16-1:0] node1627;
	wire [16-1:0] node1628;
	wire [16-1:0] node1631;
	wire [16-1:0] node1634;
	wire [16-1:0] node1635;
	wire [16-1:0] node1636;
	wire [16-1:0] node1637;
	wire [16-1:0] node1640;
	wire [16-1:0] node1643;
	wire [16-1:0] node1644;
	wire [16-1:0] node1647;
	wire [16-1:0] node1650;
	wire [16-1:0] node1651;
	wire [16-1:0] node1652;
	wire [16-1:0] node1655;
	wire [16-1:0] node1658;
	wire [16-1:0] node1659;
	wire [16-1:0] node1662;
	wire [16-1:0] node1665;
	wire [16-1:0] node1666;
	wire [16-1:0] node1667;
	wire [16-1:0] node1668;
	wire [16-1:0] node1669;
	wire [16-1:0] node1670;
	wire [16-1:0] node1673;
	wire [16-1:0] node1676;
	wire [16-1:0] node1677;
	wire [16-1:0] node1680;
	wire [16-1:0] node1683;
	wire [16-1:0] node1684;
	wire [16-1:0] node1685;
	wire [16-1:0] node1688;
	wire [16-1:0] node1691;
	wire [16-1:0] node1692;
	wire [16-1:0] node1695;
	wire [16-1:0] node1698;
	wire [16-1:0] node1699;
	wire [16-1:0] node1700;
	wire [16-1:0] node1701;
	wire [16-1:0] node1704;
	wire [16-1:0] node1707;
	wire [16-1:0] node1708;
	wire [16-1:0] node1711;
	wire [16-1:0] node1714;
	wire [16-1:0] node1715;
	wire [16-1:0] node1716;
	wire [16-1:0] node1719;
	wire [16-1:0] node1722;
	wire [16-1:0] node1723;
	wire [16-1:0] node1726;
	wire [16-1:0] node1729;
	wire [16-1:0] node1730;
	wire [16-1:0] node1731;
	wire [16-1:0] node1732;
	wire [16-1:0] node1733;
	wire [16-1:0] node1736;
	wire [16-1:0] node1739;
	wire [16-1:0] node1740;
	wire [16-1:0] node1743;
	wire [16-1:0] node1746;
	wire [16-1:0] node1747;
	wire [16-1:0] node1748;
	wire [16-1:0] node1751;
	wire [16-1:0] node1754;
	wire [16-1:0] node1755;
	wire [16-1:0] node1758;
	wire [16-1:0] node1761;
	wire [16-1:0] node1762;
	wire [16-1:0] node1763;
	wire [16-1:0] node1764;
	wire [16-1:0] node1767;
	wire [16-1:0] node1770;
	wire [16-1:0] node1771;
	wire [16-1:0] node1774;
	wire [16-1:0] node1777;
	wire [16-1:0] node1778;
	wire [16-1:0] node1779;
	wire [16-1:0] node1782;
	wire [16-1:0] node1785;
	wire [16-1:0] node1786;
	wire [16-1:0] node1789;
	wire [16-1:0] node1792;
	wire [16-1:0] node1793;
	wire [16-1:0] node1794;
	wire [16-1:0] node1795;
	wire [16-1:0] node1796;
	wire [16-1:0] node1797;
	wire [16-1:0] node1798;
	wire [16-1:0] node1801;
	wire [16-1:0] node1804;
	wire [16-1:0] node1805;
	wire [16-1:0] node1808;
	wire [16-1:0] node1811;
	wire [16-1:0] node1812;
	wire [16-1:0] node1813;
	wire [16-1:0] node1816;
	wire [16-1:0] node1819;
	wire [16-1:0] node1820;
	wire [16-1:0] node1823;
	wire [16-1:0] node1826;
	wire [16-1:0] node1827;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1832;
	wire [16-1:0] node1835;
	wire [16-1:0] node1836;
	wire [16-1:0] node1839;
	wire [16-1:0] node1842;
	wire [16-1:0] node1843;
	wire [16-1:0] node1844;
	wire [16-1:0] node1847;
	wire [16-1:0] node1850;
	wire [16-1:0] node1851;
	wire [16-1:0] node1854;
	wire [16-1:0] node1857;
	wire [16-1:0] node1858;
	wire [16-1:0] node1859;
	wire [16-1:0] node1860;
	wire [16-1:0] node1861;
	wire [16-1:0] node1864;
	wire [16-1:0] node1867;
	wire [16-1:0] node1868;
	wire [16-1:0] node1871;
	wire [16-1:0] node1874;
	wire [16-1:0] node1875;
	wire [16-1:0] node1876;
	wire [16-1:0] node1879;
	wire [16-1:0] node1882;
	wire [16-1:0] node1883;
	wire [16-1:0] node1886;
	wire [16-1:0] node1889;
	wire [16-1:0] node1890;
	wire [16-1:0] node1891;
	wire [16-1:0] node1892;
	wire [16-1:0] node1895;
	wire [16-1:0] node1898;
	wire [16-1:0] node1899;
	wire [16-1:0] node1902;
	wire [16-1:0] node1905;
	wire [16-1:0] node1906;
	wire [16-1:0] node1907;
	wire [16-1:0] node1910;
	wire [16-1:0] node1913;
	wire [16-1:0] node1914;
	wire [16-1:0] node1917;
	wire [16-1:0] node1920;
	wire [16-1:0] node1921;
	wire [16-1:0] node1922;
	wire [16-1:0] node1923;
	wire [16-1:0] node1924;
	wire [16-1:0] node1925;
	wire [16-1:0] node1928;
	wire [16-1:0] node1931;
	wire [16-1:0] node1932;
	wire [16-1:0] node1935;
	wire [16-1:0] node1938;
	wire [16-1:0] node1939;
	wire [16-1:0] node1940;
	wire [16-1:0] node1943;
	wire [16-1:0] node1946;
	wire [16-1:0] node1947;
	wire [16-1:0] node1950;
	wire [16-1:0] node1953;
	wire [16-1:0] node1954;
	wire [16-1:0] node1955;
	wire [16-1:0] node1956;
	wire [16-1:0] node1959;
	wire [16-1:0] node1962;
	wire [16-1:0] node1963;
	wire [16-1:0] node1966;
	wire [16-1:0] node1969;
	wire [16-1:0] node1970;
	wire [16-1:0] node1971;
	wire [16-1:0] node1974;
	wire [16-1:0] node1977;
	wire [16-1:0] node1978;
	wire [16-1:0] node1981;
	wire [16-1:0] node1984;
	wire [16-1:0] node1985;
	wire [16-1:0] node1986;
	wire [16-1:0] node1987;
	wire [16-1:0] node1988;
	wire [16-1:0] node1991;
	wire [16-1:0] node1994;
	wire [16-1:0] node1995;
	wire [16-1:0] node1998;
	wire [16-1:0] node2001;
	wire [16-1:0] node2002;
	wire [16-1:0] node2003;
	wire [16-1:0] node2006;
	wire [16-1:0] node2009;
	wire [16-1:0] node2010;
	wire [16-1:0] node2013;
	wire [16-1:0] node2016;
	wire [16-1:0] node2017;
	wire [16-1:0] node2018;
	wire [16-1:0] node2019;
	wire [16-1:0] node2022;
	wire [16-1:0] node2025;
	wire [16-1:0] node2026;
	wire [16-1:0] node2029;
	wire [16-1:0] node2032;
	wire [16-1:0] node2033;
	wire [16-1:0] node2034;
	wire [16-1:0] node2037;
	wire [16-1:0] node2040;
	wire [16-1:0] node2041;
	wire [16-1:0] node2044;

	assign outp = (inp[15]) ? node1024 : node1;
		assign node1 = (inp[4]) ? node513 : node2;
			assign node2 = (inp[6]) ? node258 : node3;
				assign node3 = (inp[12]) ? node131 : node4;
					assign node4 = (inp[10]) ? node68 : node5;
						assign node5 = (inp[5]) ? node37 : node6;
							assign node6 = (inp[2]) ? node22 : node7;
								assign node7 = (inp[9]) ? node15 : node8;
									assign node8 = (inp[0]) ? node12 : node9;
										assign node9 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
										assign node12 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
									assign node15 = (inp[14]) ? node19 : node16;
										assign node16 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node19 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
								assign node22 = (inp[3]) ? node30 : node23;
									assign node23 = (inp[11]) ? node27 : node24;
										assign node24 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node27 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node30 = (inp[0]) ? node34 : node31;
										assign node31 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node34 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
							assign node37 = (inp[14]) ? node53 : node38;
								assign node38 = (inp[2]) ? node46 : node39;
									assign node39 = (inp[11]) ? node43 : node40;
										assign node40 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node43 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node46 = (inp[8]) ? node50 : node47;
										assign node47 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node50 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node53 = (inp[13]) ? node61 : node54;
									assign node54 = (inp[7]) ? node58 : node55;
										assign node55 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node58 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node61 = (inp[3]) ? node65 : node62;
										assign node62 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node65 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
						assign node68 = (inp[11]) ? node100 : node69;
							assign node69 = (inp[3]) ? node85 : node70;
								assign node70 = (inp[5]) ? node78 : node71;
									assign node71 = (inp[0]) ? node75 : node72;
										assign node72 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node75 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node78 = (inp[0]) ? node82 : node79;
										assign node79 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node82 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node85 = (inp[2]) ? node93 : node86;
									assign node86 = (inp[13]) ? node90 : node87;
										assign node87 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node90 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node93 = (inp[13]) ? node97 : node94;
										assign node94 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node97 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node100 = (inp[0]) ? node116 : node101;
								assign node101 = (inp[14]) ? node109 : node102;
									assign node102 = (inp[9]) ? node106 : node103;
										assign node103 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node106 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node109 = (inp[5]) ? node113 : node110;
										assign node110 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node113 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node116 = (inp[2]) ? node124 : node117;
									assign node117 = (inp[9]) ? node121 : node118;
										assign node118 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node121 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node124 = (inp[13]) ? node128 : node125;
										assign node125 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node128 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
					assign node131 = (inp[9]) ? node195 : node132;
						assign node132 = (inp[5]) ? node164 : node133;
							assign node133 = (inp[0]) ? node149 : node134;
								assign node134 = (inp[11]) ? node142 : node135;
									assign node135 = (inp[1]) ? node139 : node136;
										assign node136 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node139 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node142 = (inp[13]) ? node146 : node143;
										assign node143 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node146 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node149 = (inp[2]) ? node157 : node150;
									assign node150 = (inp[11]) ? node154 : node151;
										assign node151 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node154 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node157 = (inp[1]) ? node161 : node158;
										assign node158 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node161 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node164 = (inp[2]) ? node180 : node165;
								assign node165 = (inp[11]) ? node173 : node166;
									assign node166 = (inp[10]) ? node170 : node167;
										assign node167 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node170 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node173 = (inp[10]) ? node177 : node174;
										assign node174 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node177 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node180 = (inp[7]) ? node188 : node181;
									assign node181 = (inp[3]) ? node185 : node182;
										assign node182 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node185 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node188 = (inp[0]) ? node192 : node189;
										assign node189 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node192 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node195 = (inp[10]) ? node227 : node196;
							assign node196 = (inp[3]) ? node212 : node197;
								assign node197 = (inp[14]) ? node205 : node198;
									assign node198 = (inp[13]) ? node202 : node199;
										assign node199 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node202 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node205 = (inp[2]) ? node209 : node206;
										assign node206 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node209 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node212 = (inp[13]) ? node220 : node213;
									assign node213 = (inp[7]) ? node217 : node214;
										assign node214 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node217 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node220 = (inp[8]) ? node224 : node221;
										assign node221 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node224 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node227 = (inp[13]) ? node243 : node228;
								assign node228 = (inp[0]) ? node236 : node229;
									assign node229 = (inp[5]) ? node233 : node230;
										assign node230 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node233 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node236 = (inp[8]) ? node240 : node237;
										assign node237 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node240 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node243 = (inp[5]) ? node251 : node244;
									assign node244 = (inp[8]) ? node248 : node245;
										assign node245 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node248 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node251 = (inp[2]) ? node255 : node252;
										assign node252 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node255 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
				assign node258 = (inp[5]) ? node386 : node259;
					assign node259 = (inp[1]) ? node323 : node260;
						assign node260 = (inp[0]) ? node292 : node261;
							assign node261 = (inp[2]) ? node277 : node262;
								assign node262 = (inp[3]) ? node270 : node263;
									assign node263 = (inp[7]) ? node267 : node264;
										assign node264 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node267 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node270 = (inp[8]) ? node274 : node271;
										assign node271 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node274 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node277 = (inp[10]) ? node285 : node278;
									assign node278 = (inp[14]) ? node282 : node279;
										assign node279 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node282 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node285 = (inp[9]) ? node289 : node286;
										assign node286 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node289 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node292 = (inp[13]) ? node308 : node293;
								assign node293 = (inp[3]) ? node301 : node294;
									assign node294 = (inp[11]) ? node298 : node295;
										assign node295 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node298 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node301 = (inp[12]) ? node305 : node302;
										assign node302 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node305 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node308 = (inp[3]) ? node316 : node309;
									assign node309 = (inp[14]) ? node313 : node310;
										assign node310 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node313 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node316 = (inp[14]) ? node320 : node317;
										assign node317 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node320 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node323 = (inp[8]) ? node355 : node324;
							assign node324 = (inp[14]) ? node340 : node325;
								assign node325 = (inp[11]) ? node333 : node326;
									assign node326 = (inp[9]) ? node330 : node327;
										assign node327 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node330 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node333 = (inp[7]) ? node337 : node334;
										assign node334 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node337 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node340 = (inp[12]) ? node348 : node341;
									assign node341 = (inp[7]) ? node345 : node342;
										assign node342 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node345 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node348 = (inp[11]) ? node352 : node349;
										assign node349 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node352 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node355 = (inp[9]) ? node371 : node356;
								assign node356 = (inp[14]) ? node364 : node357;
									assign node357 = (inp[7]) ? node361 : node358;
										assign node358 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node361 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node364 = (inp[0]) ? node368 : node365;
										assign node365 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node368 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node371 = (inp[11]) ? node379 : node372;
									assign node372 = (inp[12]) ? node376 : node373;
										assign node373 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node376 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node379 = (inp[10]) ? node383 : node380;
										assign node380 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node383 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node386 = (inp[3]) ? node450 : node387;
						assign node387 = (inp[13]) ? node419 : node388;
							assign node388 = (inp[9]) ? node404 : node389;
								assign node389 = (inp[12]) ? node397 : node390;
									assign node390 = (inp[2]) ? node394 : node391;
										assign node391 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node394 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node397 = (inp[8]) ? node401 : node398;
										assign node398 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node401 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node404 = (inp[0]) ? node412 : node405;
									assign node405 = (inp[7]) ? node409 : node406;
										assign node406 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node409 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node412 = (inp[14]) ? node416 : node413;
										assign node413 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node416 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node419 = (inp[0]) ? node435 : node420;
								assign node420 = (inp[10]) ? node428 : node421;
									assign node421 = (inp[8]) ? node425 : node422;
										assign node422 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node425 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node428 = (inp[9]) ? node432 : node429;
										assign node429 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node432 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node435 = (inp[12]) ? node443 : node436;
									assign node436 = (inp[2]) ? node440 : node437;
										assign node437 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node440 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node443 = (inp[8]) ? node447 : node444;
										assign node444 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node447 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node450 = (inp[7]) ? node482 : node451;
							assign node451 = (inp[14]) ? node467 : node452;
								assign node452 = (inp[13]) ? node460 : node453;
									assign node453 = (inp[8]) ? node457 : node454;
										assign node454 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node457 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node460 = (inp[1]) ? node464 : node461;
										assign node461 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node464 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node467 = (inp[12]) ? node475 : node468;
									assign node468 = (inp[1]) ? node472 : node469;
										assign node469 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node472 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node475 = (inp[2]) ? node479 : node476;
										assign node476 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node479 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node482 = (inp[10]) ? node498 : node483;
								assign node483 = (inp[2]) ? node491 : node484;
									assign node484 = (inp[1]) ? node488 : node485;
										assign node485 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node488 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node491 = (inp[13]) ? node495 : node492;
										assign node492 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node495 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node498 = (inp[9]) ? node506 : node499;
									assign node499 = (inp[2]) ? node503 : node500;
										assign node500 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node503 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node506 = (inp[12]) ? node510 : node507;
										assign node507 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node510 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
			assign node513 = (inp[11]) ? node769 : node514;
				assign node514 = (inp[2]) ? node642 : node515;
					assign node515 = (inp[9]) ? node579 : node516;
						assign node516 = (inp[1]) ? node548 : node517;
							assign node517 = (inp[0]) ? node533 : node518;
								assign node518 = (inp[6]) ? node526 : node519;
									assign node519 = (inp[14]) ? node523 : node520;
										assign node520 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node523 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node526 = (inp[13]) ? node530 : node527;
										assign node527 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node530 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node533 = (inp[14]) ? node541 : node534;
									assign node534 = (inp[7]) ? node538 : node535;
										assign node535 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node538 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node541 = (inp[8]) ? node545 : node542;
										assign node542 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node545 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node548 = (inp[8]) ? node564 : node549;
								assign node549 = (inp[5]) ? node557 : node550;
									assign node550 = (inp[6]) ? node554 : node551;
										assign node551 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node554 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node557 = (inp[0]) ? node561 : node558;
										assign node558 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node561 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node564 = (inp[10]) ? node572 : node565;
									assign node565 = (inp[13]) ? node569 : node566;
										assign node566 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node569 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node572 = (inp[7]) ? node576 : node573;
										assign node573 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node576 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node579 = (inp[10]) ? node611 : node580;
							assign node580 = (inp[1]) ? node596 : node581;
								assign node581 = (inp[6]) ? node589 : node582;
									assign node582 = (inp[12]) ? node586 : node583;
										assign node583 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node586 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node589 = (inp[8]) ? node593 : node590;
										assign node590 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node593 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node596 = (inp[5]) ? node604 : node597;
									assign node597 = (inp[8]) ? node601 : node598;
										assign node598 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node601 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node604 = (inp[8]) ? node608 : node605;
										assign node605 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node608 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node611 = (inp[7]) ? node627 : node612;
								assign node612 = (inp[14]) ? node620 : node613;
									assign node613 = (inp[13]) ? node617 : node614;
										assign node614 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node617 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node620 = (inp[12]) ? node624 : node621;
										assign node621 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node624 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node627 = (inp[6]) ? node635 : node628;
									assign node628 = (inp[3]) ? node632 : node629;
										assign node629 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node632 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node635 = (inp[13]) ? node639 : node636;
										assign node636 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node639 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node642 = (inp[3]) ? node706 : node643;
						assign node643 = (inp[6]) ? node675 : node644;
							assign node644 = (inp[5]) ? node660 : node645;
								assign node645 = (inp[12]) ? node653 : node646;
									assign node646 = (inp[7]) ? node650 : node647;
										assign node647 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node650 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node653 = (inp[8]) ? node657 : node654;
										assign node654 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node657 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node660 = (inp[9]) ? node668 : node661;
									assign node661 = (inp[0]) ? node665 : node662;
										assign node662 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node665 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node668 = (inp[14]) ? node672 : node669;
										assign node669 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node672 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node675 = (inp[9]) ? node691 : node676;
								assign node676 = (inp[7]) ? node684 : node677;
									assign node677 = (inp[14]) ? node681 : node678;
										assign node678 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node681 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node684 = (inp[10]) ? node688 : node685;
										assign node685 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node688 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node691 = (inp[7]) ? node699 : node692;
									assign node692 = (inp[12]) ? node696 : node693;
										assign node693 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node696 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node699 = (inp[13]) ? node703 : node700;
										assign node700 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node703 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node706 = (inp[0]) ? node738 : node707;
							assign node707 = (inp[8]) ? node723 : node708;
								assign node708 = (inp[5]) ? node716 : node709;
									assign node709 = (inp[7]) ? node713 : node710;
										assign node710 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node713 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node716 = (inp[14]) ? node720 : node717;
										assign node717 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node720 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node723 = (inp[10]) ? node731 : node724;
									assign node724 = (inp[14]) ? node728 : node725;
										assign node725 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node728 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node731 = (inp[6]) ? node735 : node732;
										assign node732 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node735 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node738 = (inp[12]) ? node754 : node739;
								assign node739 = (inp[14]) ? node747 : node740;
									assign node740 = (inp[1]) ? node744 : node741;
										assign node741 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node744 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node747 = (inp[6]) ? node751 : node748;
										assign node748 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node751 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node754 = (inp[5]) ? node762 : node755;
									assign node755 = (inp[6]) ? node759 : node756;
										assign node756 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node759 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node762 = (inp[14]) ? node766 : node763;
										assign node763 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node766 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
				assign node769 = (inp[7]) ? node897 : node770;
					assign node770 = (inp[5]) ? node834 : node771;
						assign node771 = (inp[13]) ? node803 : node772;
							assign node772 = (inp[14]) ? node788 : node773;
								assign node773 = (inp[10]) ? node781 : node774;
									assign node774 = (inp[1]) ? node778 : node775;
										assign node775 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node778 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node781 = (inp[3]) ? node785 : node782;
										assign node782 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node785 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node788 = (inp[12]) ? node796 : node789;
									assign node789 = (inp[2]) ? node793 : node790;
										assign node790 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node793 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node796 = (inp[8]) ? node800 : node797;
										assign node797 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node800 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node803 = (inp[0]) ? node819 : node804;
								assign node804 = (inp[9]) ? node812 : node805;
									assign node805 = (inp[8]) ? node809 : node806;
										assign node806 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node809 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node812 = (inp[1]) ? node816 : node813;
										assign node813 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node816 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node819 = (inp[9]) ? node827 : node820;
									assign node820 = (inp[3]) ? node824 : node821;
										assign node821 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node824 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node827 = (inp[10]) ? node831 : node828;
										assign node828 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node831 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node834 = (inp[3]) ? node866 : node835;
							assign node835 = (inp[14]) ? node851 : node836;
								assign node836 = (inp[10]) ? node844 : node837;
									assign node837 = (inp[9]) ? node841 : node838;
										assign node838 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node841 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node844 = (inp[12]) ? node848 : node845;
										assign node845 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node848 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node851 = (inp[10]) ? node859 : node852;
									assign node852 = (inp[8]) ? node856 : node853;
										assign node853 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node856 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node859 = (inp[2]) ? node863 : node860;
										assign node860 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node863 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node866 = (inp[0]) ? node882 : node867;
								assign node867 = (inp[12]) ? node875 : node868;
									assign node868 = (inp[1]) ? node872 : node869;
										assign node869 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node872 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node875 = (inp[6]) ? node879 : node876;
										assign node876 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node879 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node882 = (inp[8]) ? node890 : node883;
									assign node883 = (inp[14]) ? node887 : node884;
										assign node884 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node887 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node890 = (inp[9]) ? node894 : node891;
										assign node891 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node894 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node897 = (inp[14]) ? node961 : node898;
						assign node898 = (inp[0]) ? node930 : node899;
							assign node899 = (inp[9]) ? node915 : node900;
								assign node900 = (inp[2]) ? node908 : node901;
									assign node901 = (inp[3]) ? node905 : node902;
										assign node902 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node905 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node908 = (inp[8]) ? node912 : node909;
										assign node909 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node912 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node915 = (inp[2]) ? node923 : node916;
									assign node916 = (inp[13]) ? node920 : node917;
										assign node917 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node920 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node923 = (inp[8]) ? node927 : node924;
										assign node924 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node927 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node930 = (inp[10]) ? node946 : node931;
								assign node931 = (inp[13]) ? node939 : node932;
									assign node932 = (inp[12]) ? node936 : node933;
										assign node933 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node936 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node939 = (inp[9]) ? node943 : node940;
										assign node940 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node943 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node946 = (inp[5]) ? node954 : node947;
									assign node947 = (inp[13]) ? node951 : node948;
										assign node948 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node951 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node954 = (inp[8]) ? node958 : node955;
										assign node955 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node958 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node961 = (inp[9]) ? node993 : node962;
							assign node962 = (inp[6]) ? node978 : node963;
								assign node963 = (inp[13]) ? node971 : node964;
									assign node964 = (inp[3]) ? node968 : node965;
										assign node965 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node968 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node971 = (inp[12]) ? node975 : node972;
										assign node972 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node975 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node978 = (inp[1]) ? node986 : node979;
									assign node979 = (inp[8]) ? node983 : node980;
										assign node980 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node983 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node986 = (inp[10]) ? node990 : node987;
										assign node987 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node990 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node993 = (inp[5]) ? node1009 : node994;
								assign node994 = (inp[2]) ? node1002 : node995;
									assign node995 = (inp[10]) ? node999 : node996;
										assign node996 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node999 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1002 = (inp[1]) ? node1006 : node1003;
										assign node1003 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1006 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1009 = (inp[3]) ? node1017 : node1010;
									assign node1010 = (inp[0]) ? node1014 : node1011;
										assign node1011 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1014 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1017 = (inp[13]) ? node1021 : node1018;
										assign node1018 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node1021 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
		assign node1024 = (inp[4]) ? node1536 : node1025;
			assign node1025 = (inp[13]) ? node1281 : node1026;
				assign node1026 = (inp[8]) ? node1154 : node1027;
					assign node1027 = (inp[10]) ? node1091 : node1028;
						assign node1028 = (inp[7]) ? node1060 : node1029;
							assign node1029 = (inp[2]) ? node1045 : node1030;
								assign node1030 = (inp[11]) ? node1038 : node1031;
									assign node1031 = (inp[6]) ? node1035 : node1032;
										assign node1032 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node1035 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node1038 = (inp[9]) ? node1042 : node1039;
										assign node1039 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1042 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node1045 = (inp[1]) ? node1053 : node1046;
									assign node1046 = (inp[3]) ? node1050 : node1047;
										assign node1047 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1050 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1053 = (inp[12]) ? node1057 : node1054;
										assign node1054 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1057 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node1060 = (inp[11]) ? node1076 : node1061;
								assign node1061 = (inp[14]) ? node1069 : node1062;
									assign node1062 = (inp[1]) ? node1066 : node1063;
										assign node1063 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1066 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1069 = (inp[5]) ? node1073 : node1070;
										assign node1070 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1073 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1076 = (inp[5]) ? node1084 : node1077;
									assign node1077 = (inp[14]) ? node1081 : node1078;
										assign node1078 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1081 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1084 = (inp[9]) ? node1088 : node1085;
										assign node1085 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1088 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node1091 = (inp[0]) ? node1123 : node1092;
							assign node1092 = (inp[14]) ? node1108 : node1093;
								assign node1093 = (inp[11]) ? node1101 : node1094;
									assign node1094 = (inp[3]) ? node1098 : node1095;
										assign node1095 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1098 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1101 = (inp[7]) ? node1105 : node1102;
										assign node1102 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1105 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1108 = (inp[1]) ? node1116 : node1109;
									assign node1109 = (inp[9]) ? node1113 : node1110;
										assign node1110 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1113 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1116 = (inp[5]) ? node1120 : node1117;
										assign node1117 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1120 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1123 = (inp[14]) ? node1139 : node1124;
								assign node1124 = (inp[9]) ? node1132 : node1125;
									assign node1125 = (inp[3]) ? node1129 : node1126;
										assign node1126 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1129 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1132 = (inp[5]) ? node1136 : node1133;
										assign node1133 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1136 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1139 = (inp[11]) ? node1147 : node1140;
									assign node1140 = (inp[9]) ? node1144 : node1141;
										assign node1141 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1144 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1147 = (inp[2]) ? node1151 : node1148;
										assign node1148 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1151 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node1154 = (inp[12]) ? node1218 : node1155;
						assign node1155 = (inp[11]) ? node1187 : node1156;
							assign node1156 = (inp[10]) ? node1172 : node1157;
								assign node1157 = (inp[14]) ? node1165 : node1158;
									assign node1158 = (inp[5]) ? node1162 : node1159;
										assign node1159 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1162 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1165 = (inp[6]) ? node1169 : node1166;
										assign node1166 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1169 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1172 = (inp[7]) ? node1180 : node1173;
									assign node1173 = (inp[5]) ? node1177 : node1174;
										assign node1174 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1177 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1180 = (inp[5]) ? node1184 : node1181;
										assign node1181 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1184 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1187 = (inp[9]) ? node1203 : node1188;
								assign node1188 = (inp[1]) ? node1196 : node1189;
									assign node1189 = (inp[6]) ? node1193 : node1190;
										assign node1190 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1193 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1196 = (inp[14]) ? node1200 : node1197;
										assign node1197 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1200 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1203 = (inp[7]) ? node1211 : node1204;
									assign node1204 = (inp[6]) ? node1208 : node1205;
										assign node1205 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1208 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1211 = (inp[1]) ? node1215 : node1212;
										assign node1212 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1215 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node1218 = (inp[7]) ? node1250 : node1219;
							assign node1219 = (inp[9]) ? node1235 : node1220;
								assign node1220 = (inp[10]) ? node1228 : node1221;
									assign node1221 = (inp[3]) ? node1225 : node1222;
										assign node1222 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1225 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1228 = (inp[0]) ? node1232 : node1229;
										assign node1229 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1232 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1235 = (inp[5]) ? node1243 : node1236;
									assign node1236 = (inp[14]) ? node1240 : node1237;
										assign node1237 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1240 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1243 = (inp[10]) ? node1247 : node1244;
										assign node1244 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1247 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1250 = (inp[3]) ? node1266 : node1251;
								assign node1251 = (inp[2]) ? node1259 : node1252;
									assign node1252 = (inp[9]) ? node1256 : node1253;
										assign node1253 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1256 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1259 = (inp[0]) ? node1263 : node1260;
										assign node1260 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1263 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1266 = (inp[2]) ? node1274 : node1267;
									assign node1267 = (inp[11]) ? node1271 : node1268;
										assign node1268 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1271 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1274 = (inp[1]) ? node1278 : node1275;
										assign node1275 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1278 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
				assign node1281 = (inp[2]) ? node1409 : node1282;
					assign node1282 = (inp[0]) ? node1346 : node1283;
						assign node1283 = (inp[9]) ? node1315 : node1284;
							assign node1284 = (inp[10]) ? node1300 : node1285;
								assign node1285 = (inp[11]) ? node1293 : node1286;
									assign node1286 = (inp[7]) ? node1290 : node1287;
										assign node1287 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1290 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1293 = (inp[7]) ? node1297 : node1294;
										assign node1294 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1297 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1300 = (inp[7]) ? node1308 : node1301;
									assign node1301 = (inp[14]) ? node1305 : node1302;
										assign node1302 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1305 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1308 = (inp[12]) ? node1312 : node1309;
										assign node1309 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1312 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1315 = (inp[14]) ? node1331 : node1316;
								assign node1316 = (inp[8]) ? node1324 : node1317;
									assign node1317 = (inp[6]) ? node1321 : node1318;
										assign node1318 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1321 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1324 = (inp[7]) ? node1328 : node1325;
										assign node1325 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1328 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1331 = (inp[6]) ? node1339 : node1332;
									assign node1332 = (inp[1]) ? node1336 : node1333;
										assign node1333 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1336 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1339 = (inp[12]) ? node1343 : node1340;
										assign node1340 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1343 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node1346 = (inp[14]) ? node1378 : node1347;
							assign node1347 = (inp[1]) ? node1363 : node1348;
								assign node1348 = (inp[7]) ? node1356 : node1349;
									assign node1349 = (inp[11]) ? node1353 : node1350;
										assign node1350 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1353 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1356 = (inp[6]) ? node1360 : node1357;
										assign node1357 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1360 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1363 = (inp[11]) ? node1371 : node1364;
									assign node1364 = (inp[10]) ? node1368 : node1365;
										assign node1365 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1368 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1371 = (inp[10]) ? node1375 : node1372;
										assign node1372 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1375 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1378 = (inp[3]) ? node1394 : node1379;
								assign node1379 = (inp[5]) ? node1387 : node1380;
									assign node1380 = (inp[6]) ? node1384 : node1381;
										assign node1381 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1384 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1387 = (inp[11]) ? node1391 : node1388;
										assign node1388 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1391 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1394 = (inp[10]) ? node1402 : node1395;
									assign node1395 = (inp[7]) ? node1399 : node1396;
										assign node1396 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1399 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1402 = (inp[5]) ? node1406 : node1403;
										assign node1403 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1406 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node1409 = (inp[6]) ? node1473 : node1410;
						assign node1410 = (inp[5]) ? node1442 : node1411;
							assign node1411 = (inp[14]) ? node1427 : node1412;
								assign node1412 = (inp[7]) ? node1420 : node1413;
									assign node1413 = (inp[8]) ? node1417 : node1414;
										assign node1414 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1417 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1420 = (inp[10]) ? node1424 : node1421;
										assign node1421 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1424 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1427 = (inp[12]) ? node1435 : node1428;
									assign node1428 = (inp[0]) ? node1432 : node1429;
										assign node1429 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1432 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1435 = (inp[3]) ? node1439 : node1436;
										assign node1436 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1439 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1442 = (inp[1]) ? node1458 : node1443;
								assign node1443 = (inp[8]) ? node1451 : node1444;
									assign node1444 = (inp[3]) ? node1448 : node1445;
										assign node1445 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1448 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1451 = (inp[9]) ? node1455 : node1452;
										assign node1452 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1455 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1458 = (inp[8]) ? node1466 : node1459;
									assign node1459 = (inp[11]) ? node1463 : node1460;
										assign node1460 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1463 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1466 = (inp[0]) ? node1470 : node1467;
										assign node1467 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1470 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1473 = (inp[5]) ? node1505 : node1474;
							assign node1474 = (inp[0]) ? node1490 : node1475;
								assign node1475 = (inp[9]) ? node1483 : node1476;
									assign node1476 = (inp[12]) ? node1480 : node1477;
										assign node1477 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1480 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1483 = (inp[10]) ? node1487 : node1484;
										assign node1484 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1487 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1490 = (inp[12]) ? node1498 : node1491;
									assign node1491 = (inp[10]) ? node1495 : node1492;
										assign node1492 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1495 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1498 = (inp[1]) ? node1502 : node1499;
										assign node1499 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1502 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1505 = (inp[3]) ? node1521 : node1506;
								assign node1506 = (inp[0]) ? node1514 : node1507;
									assign node1507 = (inp[12]) ? node1511 : node1508;
										assign node1508 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1511 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1514 = (inp[8]) ? node1518 : node1515;
										assign node1515 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1518 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1521 = (inp[1]) ? node1529 : node1522;
									assign node1522 = (inp[10]) ? node1526 : node1523;
										assign node1523 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1526 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1529 = (inp[9]) ? node1533 : node1530;
										assign node1530 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node1533 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
			assign node1536 = (inp[3]) ? node1792 : node1537;
				assign node1537 = (inp[6]) ? node1665 : node1538;
					assign node1538 = (inp[0]) ? node1602 : node1539;
						assign node1539 = (inp[8]) ? node1571 : node1540;
							assign node1540 = (inp[5]) ? node1556 : node1541;
								assign node1541 = (inp[7]) ? node1549 : node1542;
									assign node1542 = (inp[12]) ? node1546 : node1543;
										assign node1543 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1546 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1549 = (inp[14]) ? node1553 : node1550;
										assign node1550 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1553 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1556 = (inp[11]) ? node1564 : node1557;
									assign node1557 = (inp[9]) ? node1561 : node1558;
										assign node1558 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1561 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1564 = (inp[12]) ? node1568 : node1565;
										assign node1565 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1568 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1571 = (inp[2]) ? node1587 : node1572;
								assign node1572 = (inp[7]) ? node1580 : node1573;
									assign node1573 = (inp[11]) ? node1577 : node1574;
										assign node1574 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1577 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1580 = (inp[11]) ? node1584 : node1581;
										assign node1581 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1584 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1587 = (inp[10]) ? node1595 : node1588;
									assign node1588 = (inp[14]) ? node1592 : node1589;
										assign node1589 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1592 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1595 = (inp[13]) ? node1599 : node1596;
										assign node1596 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1599 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node1602 = (inp[13]) ? node1634 : node1603;
							assign node1603 = (inp[7]) ? node1619 : node1604;
								assign node1604 = (inp[14]) ? node1612 : node1605;
									assign node1605 = (inp[1]) ? node1609 : node1606;
										assign node1606 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1609 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1612 = (inp[10]) ? node1616 : node1613;
										assign node1613 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1616 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1619 = (inp[5]) ? node1627 : node1620;
									assign node1620 = (inp[10]) ? node1624 : node1621;
										assign node1621 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1624 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1627 = (inp[10]) ? node1631 : node1628;
										assign node1628 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1631 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1634 = (inp[5]) ? node1650 : node1635;
								assign node1635 = (inp[2]) ? node1643 : node1636;
									assign node1636 = (inp[11]) ? node1640 : node1637;
										assign node1637 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1640 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1643 = (inp[1]) ? node1647 : node1644;
										assign node1644 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1647 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1650 = (inp[8]) ? node1658 : node1651;
									assign node1651 = (inp[9]) ? node1655 : node1652;
										assign node1652 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1655 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1658 = (inp[10]) ? node1662 : node1659;
										assign node1659 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1662 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node1665 = (inp[7]) ? node1729 : node1666;
						assign node1666 = (inp[5]) ? node1698 : node1667;
							assign node1667 = (inp[1]) ? node1683 : node1668;
								assign node1668 = (inp[11]) ? node1676 : node1669;
									assign node1669 = (inp[13]) ? node1673 : node1670;
										assign node1670 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1673 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1676 = (inp[9]) ? node1680 : node1677;
										assign node1677 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1680 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1683 = (inp[2]) ? node1691 : node1684;
									assign node1684 = (inp[13]) ? node1688 : node1685;
										assign node1685 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1688 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1691 = (inp[14]) ? node1695 : node1692;
										assign node1692 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1695 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1698 = (inp[9]) ? node1714 : node1699;
								assign node1699 = (inp[11]) ? node1707 : node1700;
									assign node1700 = (inp[0]) ? node1704 : node1701;
										assign node1701 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1704 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1707 = (inp[10]) ? node1711 : node1708;
										assign node1708 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1711 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1714 = (inp[2]) ? node1722 : node1715;
									assign node1715 = (inp[13]) ? node1719 : node1716;
										assign node1716 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1719 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1722 = (inp[1]) ? node1726 : node1723;
										assign node1723 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1726 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1729 = (inp[12]) ? node1761 : node1730;
							assign node1730 = (inp[0]) ? node1746 : node1731;
								assign node1731 = (inp[14]) ? node1739 : node1732;
									assign node1732 = (inp[11]) ? node1736 : node1733;
										assign node1733 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1736 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1739 = (inp[8]) ? node1743 : node1740;
										assign node1740 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1743 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1746 = (inp[10]) ? node1754 : node1747;
									assign node1747 = (inp[8]) ? node1751 : node1748;
										assign node1748 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1751 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1754 = (inp[9]) ? node1758 : node1755;
										assign node1755 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1758 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1761 = (inp[1]) ? node1777 : node1762;
								assign node1762 = (inp[10]) ? node1770 : node1763;
									assign node1763 = (inp[2]) ? node1767 : node1764;
										assign node1764 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1767 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1770 = (inp[8]) ? node1774 : node1771;
										assign node1771 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1774 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1777 = (inp[11]) ? node1785 : node1778;
									assign node1778 = (inp[9]) ? node1782 : node1779;
										assign node1779 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1782 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1785 = (inp[8]) ? node1789 : node1786;
										assign node1786 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node1789 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
				assign node1792 = (inp[10]) ? node1920 : node1793;
					assign node1793 = (inp[0]) ? node1857 : node1794;
						assign node1794 = (inp[12]) ? node1826 : node1795;
							assign node1795 = (inp[14]) ? node1811 : node1796;
								assign node1796 = (inp[5]) ? node1804 : node1797;
									assign node1797 = (inp[8]) ? node1801 : node1798;
										assign node1798 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1801 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1804 = (inp[7]) ? node1808 : node1805;
										assign node1805 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1808 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1811 = (inp[11]) ? node1819 : node1812;
									assign node1812 = (inp[9]) ? node1816 : node1813;
										assign node1813 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1816 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1819 = (inp[8]) ? node1823 : node1820;
										assign node1820 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1823 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1826 = (inp[7]) ? node1842 : node1827;
								assign node1827 = (inp[5]) ? node1835 : node1828;
									assign node1828 = (inp[6]) ? node1832 : node1829;
										assign node1829 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1832 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1835 = (inp[13]) ? node1839 : node1836;
										assign node1836 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1839 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1842 = (inp[11]) ? node1850 : node1843;
									assign node1843 = (inp[13]) ? node1847 : node1844;
										assign node1844 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1847 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1850 = (inp[9]) ? node1854 : node1851;
										assign node1851 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1854 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1857 = (inp[6]) ? node1889 : node1858;
							assign node1858 = (inp[5]) ? node1874 : node1859;
								assign node1859 = (inp[2]) ? node1867 : node1860;
									assign node1860 = (inp[8]) ? node1864 : node1861;
										assign node1861 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1864 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1867 = (inp[9]) ? node1871 : node1868;
										assign node1868 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1871 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1874 = (inp[1]) ? node1882 : node1875;
									assign node1875 = (inp[9]) ? node1879 : node1876;
										assign node1876 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1879 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1882 = (inp[13]) ? node1886 : node1883;
										assign node1883 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1886 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1889 = (inp[13]) ? node1905 : node1890;
								assign node1890 = (inp[5]) ? node1898 : node1891;
									assign node1891 = (inp[1]) ? node1895 : node1892;
										assign node1892 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1895 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1898 = (inp[1]) ? node1902 : node1899;
										assign node1899 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1902 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1905 = (inp[9]) ? node1913 : node1906;
									assign node1906 = (inp[8]) ? node1910 : node1907;
										assign node1907 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1910 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1913 = (inp[12]) ? node1917 : node1914;
										assign node1914 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node1917 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node1920 = (inp[1]) ? node1984 : node1921;
						assign node1921 = (inp[14]) ? node1953 : node1922;
							assign node1922 = (inp[0]) ? node1938 : node1923;
								assign node1923 = (inp[7]) ? node1931 : node1924;
									assign node1924 = (inp[12]) ? node1928 : node1925;
										assign node1925 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1928 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1931 = (inp[5]) ? node1935 : node1932;
										assign node1932 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1935 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1938 = (inp[8]) ? node1946 : node1939;
									assign node1939 = (inp[7]) ? node1943 : node1940;
										assign node1940 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1943 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1946 = (inp[12]) ? node1950 : node1947;
										assign node1947 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1950 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1953 = (inp[12]) ? node1969 : node1954;
								assign node1954 = (inp[6]) ? node1962 : node1955;
									assign node1955 = (inp[8]) ? node1959 : node1956;
										assign node1956 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1959 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1962 = (inp[13]) ? node1966 : node1963;
										assign node1963 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1966 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1969 = (inp[7]) ? node1977 : node1970;
									assign node1970 = (inp[13]) ? node1974 : node1971;
										assign node1971 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1974 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1977 = (inp[2]) ? node1981 : node1978;
										assign node1978 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node1981 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node1984 = (inp[5]) ? node2016 : node1985;
							assign node1985 = (inp[6]) ? node2001 : node1986;
								assign node1986 = (inp[14]) ? node1994 : node1987;
									assign node1987 = (inp[12]) ? node1991 : node1988;
										assign node1988 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1991 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1994 = (inp[7]) ? node1998 : node1995;
										assign node1995 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1998 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node2001 = (inp[7]) ? node2009 : node2002;
									assign node2002 = (inp[0]) ? node2006 : node2003;
										assign node2003 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2006 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2009 = (inp[13]) ? node2013 : node2010;
										assign node2010 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2013 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node2016 = (inp[12]) ? node2032 : node2017;
								assign node2017 = (inp[13]) ? node2025 : node2018;
									assign node2018 = (inp[7]) ? node2022 : node2019;
										assign node2019 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2022 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2025 = (inp[11]) ? node2029 : node2026;
										assign node2026 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2029 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node2032 = (inp[2]) ? node2040 : node2033;
									assign node2033 = (inp[9]) ? node2037 : node2034;
										assign node2034 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2037 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node2040 = (inp[14]) ? node2044 : node2041;
										assign node2041 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node2044 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;

endmodule