module dtc_split875_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node12;
	wire [14-1:0] node14;
	wire [14-1:0] node17;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node30;
	wire [14-1:0] node32;
	wire [14-1:0] node34;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node47;
	wire [14-1:0] node49;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node64;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node71;
	wire [14-1:0] node78;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node84;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node92;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node101;
	wire [14-1:0] node106;
	wire [14-1:0] node108;
	wire [14-1:0] node109;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node117;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node123;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node132;
	wire [14-1:0] node134;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node137;
	wire [14-1:0] node143;
	wire [14-1:0] node145;
	wire [14-1:0] node146;
	wire [14-1:0] node148;
	wire [14-1:0] node149;
	wire [14-1:0] node150;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node165;
	wire [14-1:0] node166;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node176;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node180;
	wire [14-1:0] node182;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node198;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node209;
	wire [14-1:0] node215;
	wire [14-1:0] node216;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node220;
	wire [14-1:0] node221;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node232;
	wire [14-1:0] node233;
	wire [14-1:0] node234;
	wire [14-1:0] node236;
	wire [14-1:0] node238;
	wire [14-1:0] node243;
	wire [14-1:0] node244;
	wire [14-1:0] node245;
	wire [14-1:0] node246;
	wire [14-1:0] node248;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node259;
	wire [14-1:0] node261;
	wire [14-1:0] node262;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node272;
	wire [14-1:0] node274;
	wire [14-1:0] node276;
	wire [14-1:0] node277;
	wire [14-1:0] node278;
	wire [14-1:0] node284;
	wire [14-1:0] node286;
	wire [14-1:0] node287;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node295;
	wire [14-1:0] node297;
	wire [14-1:0] node301;
	wire [14-1:0] node302;
	wire [14-1:0] node303;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node311;
	wire [14-1:0] node315;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node319;
	wire [14-1:0] node321;
	wire [14-1:0] node322;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node326;
	wire [14-1:0] node328;
	wire [14-1:0] node334;
	wire [14-1:0] node335;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node341;
	wire [14-1:0] node344;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node348;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node362;
	wire [14-1:0] node364;
	wire [14-1:0] node366;
	wire [14-1:0] node368;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node372;
	wire [14-1:0] node377;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node390;
	wire [14-1:0] node392;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node397;
	wire [14-1:0] node402;
	wire [14-1:0] node403;
	wire [14-1:0] node404;
	wire [14-1:0] node405;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node413;
	wire [14-1:0] node415;
	wire [14-1:0] node416;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node425;
	wire [14-1:0] node428;
	wire [14-1:0] node434;
	wire [14-1:0] node436;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node447;
	wire [14-1:0] node449;
	wire [14-1:0] node452;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node457;
	wire [14-1:0] node463;
	wire [14-1:0] node464;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node470;
	wire [14-1:0] node471;
	wire [14-1:0] node474;
	wire [14-1:0] node475;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node484;
	wire [14-1:0] node487;
	wire [14-1:0] node488;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node504;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node508;
	wire [14-1:0] node511;
	wire [14-1:0] node512;
	wire [14-1:0] node513;
	wire [14-1:0] node515;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node524;
	wire [14-1:0] node525;
	wire [14-1:0] node526;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node531;
	wire [14-1:0] node532;
	wire [14-1:0] node533;
	wire [14-1:0] node537;
	wire [14-1:0] node538;
	wire [14-1:0] node541;
	wire [14-1:0] node544;
	wire [14-1:0] node548;
	wire [14-1:0] node550;
	wire [14-1:0] node552;
	wire [14-1:0] node554;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node559;
	wire [14-1:0] node561;
	wire [14-1:0] node563;
	wire [14-1:0] node566;
	wire [14-1:0] node567;
	wire [14-1:0] node568;
	wire [14-1:0] node572;
	wire [14-1:0] node574;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node579;
	wire [14-1:0] node580;
	wire [14-1:0] node586;
	wire [14-1:0] node590;
	wire [14-1:0] node591;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node595;
	wire [14-1:0] node596;
	wire [14-1:0] node601;
	wire [14-1:0] node603;
	wire [14-1:0] node605;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node611;
	wire [14-1:0] node612;
	wire [14-1:0] node613;
	wire [14-1:0] node618;
	wire [14-1:0] node620;
	wire [14-1:0] node622;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node628;
	wire [14-1:0] node633;
	wire [14-1:0] node635;
	wire [14-1:0] node637;
	wire [14-1:0] node640;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node649;
	wire [14-1:0] node651;
	wire [14-1:0] node653;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node660;
	wire [14-1:0] node665;
	wire [14-1:0] node667;
	wire [14-1:0] node669;
	wire [14-1:0] node672;
	wire [14-1:0] node673;
	wire [14-1:0] node674;
	wire [14-1:0] node675;
	wire [14-1:0] node680;
	wire [14-1:0] node682;
	wire [14-1:0] node684;
	wire [14-1:0] node687;
	wire [14-1:0] node688;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node692;
	wire [14-1:0] node693;
	wire [14-1:0] node698;
	wire [14-1:0] node700;
	wire [14-1:0] node702;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node708;
	wire [14-1:0] node709;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node718;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node725;
	wire [14-1:0] node726;
	wire [14-1:0] node731;
	wire [14-1:0] node733;
	wire [14-1:0] node735;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node741;
	wire [14-1:0] node746;
	wire [14-1:0] node748;
	wire [14-1:0] node750;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node756;
	wire [14-1:0] node757;
	wire [14-1:0] node762;
	wire [14-1:0] node764;
	wire [14-1:0] node766;
	wire [14-1:0] node769;
	wire [14-1:0] node770;
	wire [14-1:0] node771;
	wire [14-1:0] node772;
	wire [14-1:0] node778;
	wire [14-1:0] node779;
	wire [14-1:0] node780;
	wire [14-1:0] node781;
	wire [14-1:0] node786;
	wire [14-1:0] node788;
	wire [14-1:0] node790;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node800;
	wire [14-1:0] node801;
	wire [14-1:0] node802;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node815;
	wire [14-1:0] node816;
	wire [14-1:0] node817;
	wire [14-1:0] node818;
	wire [14-1:0] node819;
	wire [14-1:0] node820;
	wire [14-1:0] node821;
	wire [14-1:0] node822;
	wire [14-1:0] node829;
	wire [14-1:0] node832;
	wire [14-1:0] node833;
	wire [14-1:0] node837;
	wire [14-1:0] node838;
	wire [14-1:0] node839;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node857;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node863;
	wire [14-1:0] node864;
	wire [14-1:0] node865;
	wire [14-1:0] node866;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node872;
	wire [14-1:0] node876;
	wire [14-1:0] node878;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node882;
	wire [14-1:0] node884;
	wire [14-1:0] node888;
	wire [14-1:0] node889;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node895;
	wire [14-1:0] node896;
	wire [14-1:0] node900;
	wire [14-1:0] node903;
	wire [14-1:0] node904;
	wire [14-1:0] node909;
	wire [14-1:0] node910;
	wire [14-1:0] node911;
	wire [14-1:0] node912;
	wire [14-1:0] node913;
	wire [14-1:0] node914;
	wire [14-1:0] node918;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node922;
	wire [14-1:0] node926;
	wire [14-1:0] node928;
	wire [14-1:0] node931;
	wire [14-1:0] node933;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node940;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node946;
	wire [14-1:0] node947;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node959;
	wire [14-1:0] node960;
	wire [14-1:0] node961;
	wire [14-1:0] node962;
	wire [14-1:0] node963;
	wire [14-1:0] node965;
	wire [14-1:0] node967;
	wire [14-1:0] node970;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node977;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node985;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node997;
	wire [14-1:0] node998;
	wire [14-1:0] node999;
	wire [14-1:0] node1000;
	wire [14-1:0] node1001;
	wire [14-1:0] node1003;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1012;
	wire [14-1:0] node1013;
	wire [14-1:0] node1014;
	wire [14-1:0] node1020;
	wire [14-1:0] node1022;
	wire [14-1:0] node1023;
	wire [14-1:0] node1025;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1029;
	wire [14-1:0] node1034;
	wire [14-1:0] node1037;
	wire [14-1:0] node1038;
	wire [14-1:0] node1039;
	wire [14-1:0] node1040;
	wire [14-1:0] node1041;
	wire [14-1:0] node1042;
	wire [14-1:0] node1043;
	wire [14-1:0] node1046;
	wire [14-1:0] node1047;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1055;
	wire [14-1:0] node1056;
	wire [14-1:0] node1057;
	wire [14-1:0] node1060;
	wire [14-1:0] node1061;
	wire [14-1:0] node1065;
	wire [14-1:0] node1066;
	wire [14-1:0] node1070;
	wire [14-1:0] node1071;
	wire [14-1:0] node1072;
	wire [14-1:0] node1073;
	wire [14-1:0] node1077;
	wire [14-1:0] node1078;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1084;
	wire [14-1:0] node1088;
	wire [14-1:0] node1089;
	wire [14-1:0] node1090;
	wire [14-1:0] node1094;
	wire [14-1:0] node1097;
	wire [14-1:0] node1098;
	wire [14-1:0] node1099;
	wire [14-1:0] node1100;
	wire [14-1:0] node1105;
	wire [14-1:0] node1107;
	wire [14-1:0] node1109;
	wire [14-1:0] node1112;
	wire [14-1:0] node1113;
	wire [14-1:0] node1114;
	wire [14-1:0] node1115;
	wire [14-1:0] node1116;
	wire [14-1:0] node1121;
	wire [14-1:0] node1123;
	wire [14-1:0] node1125;
	wire [14-1:0] node1128;
	wire [14-1:0] node1129;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1136;
	wire [14-1:0] node1138;
	wire [14-1:0] node1140;
	wire [14-1:0] node1143;
	wire [14-1:0] node1144;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1147;
	wire [14-1:0] node1152;
	wire [14-1:0] node1154;
	wire [14-1:0] node1156;
	wire [14-1:0] node1159;
	wire [14-1:0] node1160;
	wire [14-1:0] node1161;
	wire [14-1:0] node1162;
	wire [14-1:0] node1167;
	wire [14-1:0] node1169;
	wire [14-1:0] node1171;
	wire [14-1:0] node1174;
	wire [14-1:0] node1175;
	wire [14-1:0] node1176;
	wire [14-1:0] node1177;
	wire [14-1:0] node1178;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1185;
	wire [14-1:0] node1187;
	wire [14-1:0] node1189;
	wire [14-1:0] node1192;
	wire [14-1:0] node1193;
	wire [14-1:0] node1194;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1197;
	wire [14-1:0] node1202;
	wire [14-1:0] node1204;
	wire [14-1:0] node1206;
	wire [14-1:0] node1209;
	wire [14-1:0] node1210;
	wire [14-1:0] node1211;
	wire [14-1:0] node1212;
	wire [14-1:0] node1217;
	wire [14-1:0] node1219;
	wire [14-1:0] node1221;
	wire [14-1:0] node1224;
	wire [14-1:0] node1225;
	wire [14-1:0] node1226;
	wire [14-1:0] node1227;
	wire [14-1:0] node1228;
	wire [14-1:0] node1229;
	wire [14-1:0] node1234;
	wire [14-1:0] node1236;
	wire [14-1:0] node1238;
	wire [14-1:0] node1241;
	wire [14-1:0] node1242;
	wire [14-1:0] node1243;
	wire [14-1:0] node1244;
	wire [14-1:0] node1245;
	wire [14-1:0] node1250;
	wire [14-1:0] node1252;
	wire [14-1:0] node1254;
	wire [14-1:0] node1257;
	wire [14-1:0] node1258;
	wire [14-1:0] node1259;
	wire [14-1:0] node1260;
	wire [14-1:0] node1265;
	wire [14-1:0] node1267;
	wire [14-1:0] node1269;
	wire [14-1:0] node1272;
	wire [14-1:0] node1273;
	wire [14-1:0] node1274;
	wire [14-1:0] node1275;
	wire [14-1:0] node1276;
	wire [14-1:0] node1281;
	wire [14-1:0] node1283;
	wire [14-1:0] node1285;
	wire [14-1:0] node1288;
	wire [14-1:0] node1289;
	wire [14-1:0] node1290;
	wire [14-1:0] node1291;
	wire [14-1:0] node1292;
	wire [14-1:0] node1297;
	wire [14-1:0] node1299;
	wire [14-1:0] node1301;
	wire [14-1:0] node1304;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1310;
	wire [14-1:0] node1312;
	wire [14-1:0] node1314;
	wire [14-1:0] node1317;
	wire [14-1:0] node1318;
	wire [14-1:0] node1319;
	wire [14-1:0] node1320;
	wire [14-1:0] node1323;
	wire [14-1:0] node1324;
	wire [14-1:0] node1325;
	wire [14-1:0] node1326;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1334;
	wire [14-1:0] node1335;
	wire [14-1:0] node1336;
	wire [14-1:0] node1343;
	wire [14-1:0] node1345;
	wire [14-1:0] node1347;
	wire [14-1:0] node1350;
	wire [14-1:0] node1351;
	wire [14-1:0] node1352;
	wire [14-1:0] node1353;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1356;
	wire [14-1:0] node1359;
	wire [14-1:0] node1360;
	wire [14-1:0] node1363;
	wire [14-1:0] node1366;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1371;
	wire [14-1:0] node1373;
	wire [14-1:0] node1377;
	wire [14-1:0] node1378;
	wire [14-1:0] node1379;
	wire [14-1:0] node1380;
	wire [14-1:0] node1383;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1391;
	wire [14-1:0] node1392;
	wire [14-1:0] node1393;
	wire [14-1:0] node1397;
	wire [14-1:0] node1398;
	wire [14-1:0] node1399;
	wire [14-1:0] node1403;
	wire [14-1:0] node1406;
	wire [14-1:0] node1407;
	wire [14-1:0] node1408;
	wire [14-1:0] node1409;
	wire [14-1:0] node1410;
	wire [14-1:0] node1415;
	wire [14-1:0] node1417;
	wire [14-1:0] node1419;
	wire [14-1:0] node1422;
	wire [14-1:0] node1423;
	wire [14-1:0] node1424;
	wire [14-1:0] node1425;
	wire [14-1:0] node1426;
	wire [14-1:0] node1431;
	wire [14-1:0] node1433;
	wire [14-1:0] node1435;
	wire [14-1:0] node1438;
	wire [14-1:0] node1439;
	wire [14-1:0] node1440;
	wire [14-1:0] node1441;
	wire [14-1:0] node1446;
	wire [14-1:0] node1448;
	wire [14-1:0] node1450;
	wire [14-1:0] node1453;
	wire [14-1:0] node1454;
	wire [14-1:0] node1455;
	wire [14-1:0] node1456;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1463;
	wire [14-1:0] node1465;
	wire [14-1:0] node1467;
	wire [14-1:0] node1470;
	wire [14-1:0] node1471;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1474;
	wire [14-1:0] node1479;
	wire [14-1:0] node1481;
	wire [14-1:0] node1483;
	wire [14-1:0] node1486;
	wire [14-1:0] node1487;
	wire [14-1:0] node1488;
	wire [14-1:0] node1489;
	wire [14-1:0] node1494;
	wire [14-1:0] node1496;
	wire [14-1:0] node1498;
	wire [14-1:0] node1501;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1504;
	wire [14-1:0] node1505;
	wire [14-1:0] node1510;
	wire [14-1:0] node1512;
	wire [14-1:0] node1514;
	wire [14-1:0] node1517;
	wire [14-1:0] node1518;
	wire [14-1:0] node1519;
	wire [14-1:0] node1520;
	wire [14-1:0] node1525;
	wire [14-1:0] node1527;
	wire [14-1:0] node1529;
	wire [14-1:0] node1532;
	wire [14-1:0] node1533;
	wire [14-1:0] node1534;
	wire [14-1:0] node1535;
	wire [14-1:0] node1536;
	wire [14-1:0] node1541;
	wire [14-1:0] node1542;
	wire [14-1:0] node1544;
	wire [14-1:0] node1546;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1551;
	wire [14-1:0] node1554;
	wire [14-1:0] node1557;
	wire [14-1:0] node1559;
	wire [14-1:0] node1562;
	wire [14-1:0] node1563;
	wire [14-1:0] node1564;
	wire [14-1:0] node1565;
	wire [14-1:0] node1567;
	wire [14-1:0] node1568;
	wire [14-1:0] node1569;
	wire [14-1:0] node1571;
	wire [14-1:0] node1576;
	wire [14-1:0] node1577;
	wire [14-1:0] node1578;
	wire [14-1:0] node1579;
	wire [14-1:0] node1581;
	wire [14-1:0] node1584;
	wire [14-1:0] node1586;
	wire [14-1:0] node1591;
	wire [14-1:0] node1592;
	wire [14-1:0] node1593;
	wire [14-1:0] node1594;
	wire [14-1:0] node1595;
	wire [14-1:0] node1599;
	wire [14-1:0] node1600;
	wire [14-1:0] node1602;
	wire [14-1:0] node1606;
	wire [14-1:0] node1609;
	wire [14-1:0] node1610;
	wire [14-1:0] node1611;
	wire [14-1:0] node1613;
	wire [14-1:0] node1618;
	wire [14-1:0] node1620;
	wire [14-1:0] node1621;
	wire [14-1:0] node1623;
	wire [14-1:0] node1626;
	wire [14-1:0] node1627;

	assign outp = (inp[10]) ? node590 : node1;
		assign node1 = (inp[8]) ? node315 : node2;
			assign node2 = (inp[13]) ? node176 : node3;
				assign node3 = (inp[11]) ? node61 : node4;
					assign node4 = (inp[12]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[9]) ? 14'b00000000000000 : node7;
							assign node7 = (inp[2]) ? node47 : node8;
								assign node8 = (inp[7]) ? node28 : node9;
									assign node9 = (inp[1]) ? node17 : node10;
										assign node10 = (inp[3]) ? node12 : 14'b00000000000000;
											assign node12 = (inp[6]) ? node14 : 14'b00000000000000;
												assign node14 = (inp[0]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node17 = (inp[6]) ? 14'b00000000000000 : node18;
											assign node18 = (inp[5]) ? 14'b00000000000000 : node19;
												assign node19 = (inp[0]) ? node21 : 14'b00000000000000;
													assign node21 = (inp[4]) ? 14'b00000000000000 : node22;
														assign node22 = (inp[3]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node28 = (inp[3]) ? 14'b00000000000000 : node29;
										assign node29 = (inp[0]) ? node37 : node30;
											assign node30 = (inp[6]) ? node32 : 14'b00000000000000;
												assign node32 = (inp[5]) ? node34 : 14'b00000000000000;
													assign node34 = (inp[1]) ? 14'b00001000000101 : 14'b00000000000000;
											assign node37 = (inp[4]) ? 14'b00000000000000 : node38;
												assign node38 = (inp[6]) ? 14'b00000000000000 : node39;
													assign node39 = (inp[5]) ? 14'b00000000000000 : node40;
														assign node40 = (inp[1]) ? 14'b00100000000011 : 14'b00000000000000;
								assign node47 = (inp[1]) ? node49 : 14'b00000000000000;
									assign node49 = (inp[0]) ? node51 : 14'b00000000000000;
										assign node51 = (inp[3]) ? 14'b00000000000000 : node52;
											assign node52 = (inp[4]) ? 14'b00000000000000 : node53;
												assign node53 = (inp[6]) ? 14'b00000000000000 : node54;
													assign node54 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node61 = (inp[12]) ? node113 : node62;
						assign node62 = (inp[1]) ? node64 : 14'b00000000000000;
							assign node64 = (inp[7]) ? node78 : node65;
								assign node65 = (inp[9]) ? 14'b00000000000000 : node66;
									assign node66 = (inp[2]) ? node68 : 14'b00000000000000;
										assign node68 = (inp[3]) ? 14'b00000000000000 : node69;
											assign node69 = (inp[4]) ? 14'b00000000000000 : node70;
												assign node70 = (inp[6]) ? 14'b00000000000000 : node71;
													assign node71 = (inp[0]) ? 14'b00100000000011 : 14'b00000000000000;
								assign node78 = (inp[2]) ? node96 : node79;
									assign node79 = (inp[6]) ? node89 : node80;
										assign node80 = (inp[0]) ? 14'b00000000000000 : node81;
											assign node81 = (inp[9]) ? 14'b10010000001101 : node82;
												assign node82 = (inp[3]) ? node84 : 14'b00000000000000;
													assign node84 = (inp[5]) ? 14'b10010000001101 : 14'b00000000000000;
										assign node89 = (inp[5]) ? 14'b00000000000000 : node90;
											assign node90 = (inp[9]) ? node92 : 14'b00000000000000;
												assign node92 = (inp[3]) ? 14'b01001000000100 : 14'b00000000000000;
									assign node96 = (inp[3]) ? node106 : node97;
										assign node97 = (inp[0]) ? node99 : 14'b00000000000000;
											assign node99 = (inp[9]) ? 14'b00000000000000 : node100;
												assign node100 = (inp[6]) ? 14'b00000000000000 : node101;
													assign node101 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node106 = (inp[6]) ? node108 : 14'b00000000000000;
											assign node108 = (inp[5]) ? 14'b00000000000000 : node109;
												assign node109 = (inp[9]) ? 14'b01001000000100 : 14'b00000000000000;
						assign node113 = (inp[9]) ? node143 : node114;
							assign node114 = (inp[3]) ? node128 : node115;
								assign node115 = (inp[1]) ? node117 : 14'b00000000000000;
									assign node117 = (inp[6]) ? node119 : 14'b10000100011000;
										assign node119 = (inp[0]) ? 14'b00000000000000 : node120;
											assign node120 = (inp[2]) ? 14'b00000000000000 : node121;
												assign node121 = (inp[7]) ? node123 : 14'b00000000000000;
													assign node123 = (inp[5]) ? 14'b10100000001000 : 14'b00000000000000;
								assign node128 = (inp[1]) ? node132 : node129;
									assign node129 = (inp[6]) ? 14'b01100000001010 : 14'b00000000000000;
									assign node132 = (inp[7]) ? node134 : 14'b00000000000000;
										assign node134 = (inp[2]) ? 14'b00000000000000 : node135;
											assign node135 = (inp[0]) ? 14'b00000000000000 : node136;
												assign node136 = (inp[6]) ? 14'b00000000000000 : node137;
													assign node137 = (inp[5]) ? 14'b01001000000100 : 14'b01001000000101;
							assign node143 = (inp[1]) ? node145 : 14'b00000000000000;
								assign node145 = (inp[5]) ? node155 : node146;
									assign node146 = (inp[7]) ? node148 : 14'b00000000000000;
										assign node148 = (inp[0]) ? 14'b00000000000000 : node149;
											assign node149 = (inp[2]) ? 14'b00000000000000 : node150;
												assign node150 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000100;
									assign node155 = (inp[3]) ? node165 : node156;
										assign node156 = (inp[2]) ? 14'b00000000000000 : node157;
											assign node157 = (inp[7]) ? node159 : 14'b00000000000000;
												assign node159 = (inp[6]) ? 14'b00000000000000 : node160;
													assign node160 = (inp[0]) ? 14'b00000000000000 : 14'b01001000000100;
										assign node165 = (inp[7]) ? node169 : node166;
											assign node166 = (inp[6]) ? 14'b01001000001100 : 14'b00000000000000;
											assign node169 = (inp[0]) ? 14'b00000000000000 : node170;
												assign node170 = (inp[6]) ? 14'b00000000000000 : node171;
													assign node171 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000100;
				assign node176 = (inp[1]) ? node198 : node177;
					assign node177 = (inp[9]) ? 14'b00000000000000 : node178;
						assign node178 = (inp[3]) ? node180 : 14'b00000000000000;
							assign node180 = (inp[6]) ? node182 : 14'b00000000000000;
								assign node182 = (inp[12]) ? node188 : node183;
									assign node183 = (inp[11]) ? 14'b00000000000000 : node184;
										assign node184 = (inp[7]) ? 14'b00000000000000 : 14'b11000000000100;
									assign node188 = (inp[11]) ? 14'b00100100001101 : node189;
										assign node189 = (inp[2]) ? 14'b00000000000000 : node190;
											assign node190 = (inp[7]) ? 14'b00000000000000 : node191;
												assign node191 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
					assign node198 = (inp[6]) ? node268 : node199;
						assign node199 = (inp[3]) ? node243 : node200;
							assign node200 = (inp[9]) ? node232 : node201;
								assign node201 = (inp[11]) ? node215 : node202;
									assign node202 = (inp[12]) ? node204 : 14'b11000000000100;
										assign node204 = (inp[4]) ? 14'b00000000000000 : node205;
											assign node205 = (inp[0]) ? node207 : 14'b00000000000000;
												assign node207 = (inp[2]) ? 14'b10000000101100 : node208;
													assign node208 = (inp[5]) ? 14'b00000000000000 : node209;
														assign node209 = (inp[7]) ? 14'b10000100001100 : 14'b10010000001100;
									assign node215 = (inp[4]) ? 14'b00000000000000 : node216;
										assign node216 = (inp[0]) ? node218 : 14'b00000000000000;
											assign node218 = (inp[12]) ? node226 : node219;
												assign node219 = (inp[2]) ? 14'b10110101111111 : node220;
													assign node220 = (inp[5]) ? 14'b00000000000000 : node221;
														assign node221 = (inp[7]) ? 14'b01001000000100 : 14'b00000000000000;
												assign node226 = (inp[5]) ? 14'b00000000000000 : node227;
													assign node227 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000101;
								assign node232 = (inp[0]) ? 14'b00000000000000 : node233;
									assign node233 = (inp[2]) ? 14'b00000000000000 : node234;
										assign node234 = (inp[7]) ? node236 : 14'b00000000000000;
											assign node236 = (inp[12]) ? node238 : 14'b00000000000000;
												assign node238 = (inp[11]) ? 14'b10100010001100 : 14'b11110111110010;
							assign node243 = (inp[2]) ? 14'b00000000000000 : node244;
								assign node244 = (inp[0]) ? 14'b00000000000000 : node245;
									assign node245 = (inp[11]) ? node255 : node246;
										assign node246 = (inp[7]) ? node248 : 14'b00000000000000;
											assign node248 = (inp[12]) ? node250 : 14'b00000000000000;
												assign node250 = (inp[5]) ? 14'b11110111110010 : node251;
													assign node251 = (inp[9]) ? 14'b11110111110010 : 14'b00000000000000;
										assign node255 = (inp[12]) ? node259 : node256;
											assign node256 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
											assign node259 = (inp[7]) ? node261 : 14'b00000000000000;
												assign node261 = (inp[5]) ? 14'b10100010001100 : node262;
													assign node262 = (inp[9]) ? 14'b10100010001100 : 14'b10010101111110;
						assign node268 = (inp[3]) ? node284 : node269;
							assign node269 = (inp[9]) ? 14'b00000000000000 : node270;
								assign node270 = (inp[7]) ? node272 : 14'b00000000000000;
									assign node272 = (inp[5]) ? node274 : 14'b00000000000000;
										assign node274 = (inp[12]) ? node276 : 14'b00000000000000;
											assign node276 = (inp[0]) ? 14'b00000000000000 : node277;
												assign node277 = (inp[2]) ? 14'b00000000000000 : node278;
													assign node278 = (inp[11]) ? 14'b00001000000001 : 14'b01001000000101;
							assign node284 = (inp[9]) ? node286 : 14'b00000000000000;
								assign node286 = (inp[12]) ? node308 : node287;
									assign node287 = (inp[7]) ? node289 : 14'b00000000000000;
										assign node289 = (inp[11]) ? node301 : node290;
											assign node290 = (inp[5]) ? 14'b00000000000000 : node291;
												assign node291 = (inp[2]) ? node295 : node292;
													assign node292 = (inp[0]) ? 14'b01100000000110 : 14'b00001000000101;
													assign node295 = (inp[4]) ? node297 : 14'b01100000000110;
														assign node297 = (inp[0]) ? 14'b00000000000000 : 14'b01100000000110;
											assign node301 = (inp[5]) ? 14'b01001000000101 : node302;
												assign node302 = (inp[0]) ? 14'b10000010001100 : node303;
													assign node303 = (inp[2]) ? 14'b10000010001100 : 14'b10000100101000;
									assign node308 = (inp[7]) ? 14'b00000000000000 : node309;
										assign node309 = (inp[5]) ? node311 : 14'b00000000000000;
											assign node311 = (inp[11]) ? 14'b00000000011100 : 14'b00000000011101;
			assign node315 = (inp[12]) ? node463 : node316;
				assign node316 = (inp[1]) ? node334 : node317;
					assign node317 = (inp[3]) ? node319 : 14'b00000000000000;
						assign node319 = (inp[6]) ? node321 : 14'b00000000000000;
							assign node321 = (inp[0]) ? 14'b00000000000000 : node322;
								assign node322 = (inp[11]) ? node324 : 14'b00000000000000;
									assign node324 = (inp[9]) ? 14'b00000000000000 : node325;
										assign node325 = (inp[7]) ? 14'b00000000000000 : node326;
											assign node326 = (inp[13]) ? node328 : 14'b00000000000000;
												assign node328 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node334 = (inp[11]) ? node402 : node335;
						assign node335 = (inp[13]) ? node377 : node336;
							assign node336 = (inp[6]) ? node362 : node337;
								assign node337 = (inp[2]) ? node353 : node338;
									assign node338 = (inp[0]) ? node344 : node339;
										assign node339 = (inp[3]) ? node341 : 14'b00000000000000;
											assign node341 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
										assign node344 = (inp[7]) ? node346 : 14'b00000000000000;
											assign node346 = (inp[4]) ? 14'b00000000000000 : node347;
												assign node347 = (inp[5]) ? 14'b00000000000000 : node348;
													assign node348 = (inp[3]) ? 14'b00000000000000 : 14'b00100100001100;
									assign node353 = (inp[9]) ? 14'b00000000000000 : node354;
										assign node354 = (inp[0]) ? node356 : 14'b00000000000000;
											assign node356 = (inp[4]) ? 14'b00000000000000 : node357;
												assign node357 = (inp[3]) ? 14'b00000000000000 : 14'b10000000011010;
								assign node362 = (inp[7]) ? node364 : 14'b00000000000000;
									assign node364 = (inp[9]) ? node366 : 14'b00000000000000;
										assign node366 = (inp[3]) ? node368 : 14'b00000000000000;
											assign node368 = (inp[5]) ? 14'b00000000011100 : node369;
												assign node369 = (inp[0]) ? 14'b00000000000000 : node370;
													assign node370 = (inp[2]) ? node372 : 14'b01000000010000;
														assign node372 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node377 = (inp[7]) ? node379 : 14'b00000000000000;
								assign node379 = (inp[5]) ? 14'b00000000000000 : node380;
									assign node380 = (inp[3]) ? node390 : node381;
										assign node381 = (inp[6]) ? 14'b00000000000000 : node382;
											assign node382 = (inp[0]) ? node384 : 14'b00000000000000;
												assign node384 = (inp[4]) ? 14'b00000000000000 : node385;
													assign node385 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000101;
										assign node390 = (inp[9]) ? node392 : 14'b00000000000000;
											assign node392 = (inp[6]) ? node394 : 14'b00000000000000;
												assign node394 = (inp[0]) ? 14'b00000000000000 : node395;
													assign node395 = (inp[4]) ? node397 : 14'b00000000011100;
														assign node397 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
						assign node402 = (inp[9]) ? node434 : node403;
							assign node403 = (inp[3]) ? node421 : node404;
								assign node404 = (inp[6]) ? node408 : node405;
									assign node405 = (inp[13]) ? 14'b00000000011100 : 14'b01001000000100;
									assign node408 = (inp[13]) ? 14'b00000000000000 : node409;
										assign node409 = (inp[7]) ? node413 : node410;
											assign node410 = (inp[5]) ? 14'b00000000000000 : 14'b11000000000100;
											assign node413 = (inp[5]) ? node415 : 14'b00000000000000;
												assign node415 = (inp[2]) ? 14'b00000000000000 : node416;
													assign node416 = (inp[0]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node421 = (inp[2]) ? 14'b00000000000000 : node422;
									assign node422 = (inp[6]) ? 14'b00000000000000 : node423;
										assign node423 = (inp[7]) ? 14'b00000000000000 : node424;
											assign node424 = (inp[13]) ? node428 : node425;
												assign node425 = (inp[0]) ? 14'b00000000000000 : 14'b00000100000001;
												assign node428 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node434 = (inp[3]) ? node436 : 14'b00000000000000;
								assign node436 = (inp[5]) ? node452 : node437;
									assign node437 = (inp[7]) ? node447 : node438;
										assign node438 = (inp[2]) ? 14'b00000000000000 : node439;
											assign node439 = (inp[6]) ? 14'b00000000000000 : node440;
												assign node440 = (inp[13]) ? 14'b00000000011100 : node441;
													assign node441 = (inp[0]) ? 14'b00000000000000 : 14'b00000100000001;
										assign node447 = (inp[6]) ? node449 : 14'b00000000000000;
											assign node449 = (inp[13]) ? 14'b10100010001100 : 14'b01100000001010;
									assign node452 = (inp[6]) ? 14'b00000000000000 : node453;
										assign node453 = (inp[7]) ? 14'b00000000000000 : node454;
											assign node454 = (inp[0]) ? 14'b00000000000000 : node455;
												assign node455 = (inp[13]) ? node457 : 14'b00000100000001;
													assign node457 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
				assign node463 = (inp[11]) ? node557 : node464;
					assign node464 = (inp[6]) ? node504 : node465;
						assign node465 = (inp[2]) ? 14'b00000000000000 : node466;
							assign node466 = (inp[1]) ? node468 : 14'b00000000000000;
								assign node468 = (inp[0]) ? node492 : node469;
									assign node469 = (inp[13]) ? node479 : node470;
										assign node470 = (inp[3]) ? node474 : node471;
											assign node471 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node474 = (inp[7]) ? 14'b00000000000000 : node475;
												assign node475 = (inp[9]) ? 14'b00001000000101 : 14'b00001000000000;
										assign node479 = (inp[7]) ? node487 : node480;
											assign node480 = (inp[3]) ? node484 : node481;
												assign node481 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
												assign node484 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
											assign node487 = (inp[3]) ? 14'b00000000000000 : node488;
												assign node488 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
									assign node492 = (inp[13]) ? 14'b00000000000000 : node493;
										assign node493 = (inp[9]) ? 14'b00000000000000 : node494;
											assign node494 = (inp[4]) ? 14'b00000000000000 : node495;
												assign node495 = (inp[3]) ? 14'b00000000000000 : node496;
													assign node496 = (inp[5]) ? 14'b00000000000000 : 14'b00000000011100;
						assign node504 = (inp[13]) ? node524 : node505;
							assign node505 = (inp[1]) ? node511 : node506;
								assign node506 = (inp[9]) ? node508 : 14'b00000000000000;
									assign node508 = (inp[3]) ? 14'b11110111110010 : 14'b00000000000000;
								assign node511 = (inp[0]) ? 14'b00000000000000 : node512;
									assign node512 = (inp[9]) ? 14'b00000000000000 : node513;
										assign node513 = (inp[7]) ? node515 : 14'b00000000000000;
											assign node515 = (inp[2]) ? 14'b00000000000000 : node516;
												assign node516 = (inp[3]) ? 14'b00000000000000 : node517;
													assign node517 = (inp[5]) ? 14'b10100100111111 : 14'b00000000000000;
							assign node524 = (inp[9]) ? node548 : node525;
								assign node525 = (inp[3]) ? 14'b00000000000000 : node526;
									assign node526 = (inp[1]) ? node528 : 14'b00000000000000;
										assign node528 = (inp[5]) ? node544 : node529;
											assign node529 = (inp[7]) ? node531 : 14'b10010100011100;
												assign node531 = (inp[4]) ? node537 : node532;
													assign node532 = (inp[0]) ? 14'b00000000000000 : node533;
														assign node533 = (inp[2]) ? 14'b00000000000000 : 14'b10010010001100;
													assign node537 = (inp[2]) ? node541 : node538;
														assign node538 = (inp[0]) ? 14'b00000000000000 : 14'b10010010001100;
														assign node541 = (inp[0]) ? 14'b10010010001100 : 14'b00000000000000;
											assign node544 = (inp[7]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node548 = (inp[3]) ? node550 : 14'b00000000000000;
									assign node550 = (inp[1]) ? node552 : 14'b01001000000100;
										assign node552 = (inp[5]) ? node554 : 14'b00000000000000;
											assign node554 = (inp[7]) ? 14'b01001000001001 : 14'b00000000000000;
					assign node557 = (inp[13]) ? 14'b01000000010100 : node558;
						assign node558 = (inp[1]) ? node566 : node559;
							assign node559 = (inp[6]) ? node561 : 14'b00000000000000;
								assign node561 = (inp[3]) ? node563 : 14'b00000000000000;
									assign node563 = (inp[9]) ? 14'b10100010001100 : 14'b00000000000000;
							assign node566 = (inp[9]) ? node572 : node567;
								assign node567 = (inp[3]) ? 14'b00000000000000 : node568;
									assign node568 = (inp[6]) ? 14'b01000100000100 : 14'b00100100011111;
								assign node572 = (inp[3]) ? node574 : 14'b00000000000000;
									assign node574 = (inp[5]) ? node576 : 14'b00000000000000;
										assign node576 = (inp[7]) ? node586 : node577;
											assign node577 = (inp[0]) ? 14'b00000000000000 : node578;
												assign node578 = (inp[6]) ? 14'b00000000000000 : node579;
													assign node579 = (inp[2]) ? 14'b00000000000000 : node580;
														assign node580 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
											assign node586 = (inp[6]) ? 14'b10000000011010 : 14'b00000000000000;
		assign node590 = (inp[1]) ? node860 : node591;
			assign node591 = (inp[6]) ? node687 : node592;
				assign node592 = (inp[5]) ? node608 : node593;
					assign node593 = (inp[8]) ? node601 : node594;
						assign node594 = (inp[13]) ? 14'b00000000000000 : node595;
							assign node595 = (inp[12]) ? 14'b00000000000000 : node596;
								assign node596 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
						assign node601 = (inp[13]) ? node603 : 14'b00000000000000;
							assign node603 = (inp[11]) ? node605 : 14'b00000000000000;
								assign node605 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node608 = (inp[7]) ? node640 : node609;
						assign node609 = (inp[3]) ? node625 : node610;
							assign node610 = (inp[11]) ? node618 : node611;
								assign node611 = (inp[12]) ? 14'b00000000000000 : node612;
									assign node612 = (inp[8]) ? 14'b00000000000000 : node613;
										assign node613 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node618 = (inp[12]) ? node620 : 14'b00000000000000;
									assign node620 = (inp[8]) ? node622 : 14'b00000000000000;
										assign node622 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node625 = (inp[13]) ? node633 : node626;
								assign node626 = (inp[12]) ? 14'b00000000000000 : node627;
									assign node627 = (inp[8]) ? 14'b00000000000000 : node628;
										assign node628 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node633 = (inp[11]) ? node635 : 14'b00000000000000;
									assign node635 = (inp[8]) ? node637 : 14'b00000000000000;
										assign node637 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node640 = (inp[4]) ? node656 : node641;
							assign node641 = (inp[8]) ? node649 : node642;
								assign node642 = (inp[11]) ? 14'b00000000000000 : node643;
									assign node643 = (inp[12]) ? 14'b00000000000000 : node644;
										assign node644 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node649 = (inp[11]) ? node651 : 14'b00000000000000;
									assign node651 = (inp[13]) ? node653 : 14'b00000000000000;
										assign node653 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node656 = (inp[9]) ? node672 : node657;
								assign node657 = (inp[8]) ? node665 : node658;
									assign node658 = (inp[13]) ? 14'b00000000000000 : node659;
										assign node659 = (inp[12]) ? 14'b00000000000000 : node660;
											assign node660 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node665 = (inp[13]) ? node667 : 14'b00000000000000;
										assign node667 = (inp[12]) ? node669 : 14'b00000000000000;
											assign node669 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node672 = (inp[11]) ? node680 : node673;
									assign node673 = (inp[8]) ? 14'b00000000000000 : node674;
										assign node674 = (inp[13]) ? 14'b00000000000000 : node675;
											assign node675 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node680 = (inp[13]) ? node682 : 14'b00000000000000;
										assign node682 = (inp[12]) ? node684 : 14'b00000000000000;
											assign node684 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node687 = (inp[3]) ? node793 : node688;
					assign node688 = (inp[5]) ? node778 : node689;
						assign node689 = (inp[7]) ? node705 : node690;
							assign node690 = (inp[13]) ? node698 : node691;
								assign node691 = (inp[12]) ? 14'b00000000000000 : node692;
									assign node692 = (inp[11]) ? 14'b00000000000000 : node693;
										assign node693 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node698 = (inp[12]) ? node700 : 14'b00000000000000;
									assign node700 = (inp[11]) ? node702 : 14'b00000000000000;
										assign node702 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node705 = (inp[4]) ? node721 : node706;
								assign node706 = (inp[11]) ? node714 : node707;
									assign node707 = (inp[8]) ? 14'b00000000000000 : node708;
										assign node708 = (inp[12]) ? 14'b00000000000000 : node709;
											assign node709 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node714 = (inp[8]) ? node716 : 14'b00000000000000;
										assign node716 = (inp[13]) ? node718 : 14'b00000000000000;
											assign node718 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node721 = (inp[0]) ? node753 : node722;
									assign node722 = (inp[2]) ? node738 : node723;
										assign node723 = (inp[8]) ? node731 : node724;
											assign node724 = (inp[11]) ? 14'b00000000000000 : node725;
												assign node725 = (inp[12]) ? 14'b00000000000000 : node726;
													assign node726 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node731 = (inp[11]) ? node733 : 14'b00000000000000;
												assign node733 = (inp[13]) ? node735 : 14'b00000000000000;
													assign node735 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node738 = (inp[13]) ? node746 : node739;
											assign node739 = (inp[12]) ? 14'b00000000000000 : node740;
												assign node740 = (inp[8]) ? 14'b00000000000000 : node741;
													assign node741 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node746 = (inp[12]) ? node748 : 14'b00000000000000;
												assign node748 = (inp[11]) ? node750 : 14'b00000000000000;
													assign node750 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node753 = (inp[2]) ? node769 : node754;
										assign node754 = (inp[12]) ? node762 : node755;
											assign node755 = (inp[8]) ? 14'b00000000000000 : node756;
												assign node756 = (inp[13]) ? 14'b00000000000000 : node757;
													assign node757 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node762 = (inp[11]) ? node764 : 14'b00000000000000;
												assign node764 = (inp[13]) ? node766 : 14'b00000000000000;
													assign node766 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node769 = (inp[8]) ? 14'b00000000000000 : node770;
											assign node770 = (inp[12]) ? 14'b00000000000000 : node771;
												assign node771 = (inp[11]) ? 14'b00000000000000 : node772;
													assign node772 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
						assign node778 = (inp[11]) ? node786 : node779;
							assign node779 = (inp[8]) ? 14'b00000000000000 : node780;
								assign node780 = (inp[13]) ? 14'b00000000000000 : node781;
									assign node781 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node786 = (inp[8]) ? node788 : 14'b00000000000000;
								assign node788 = (inp[13]) ? node790 : 14'b00000000000000;
									assign node790 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node793 = (inp[12]) ? node815 : node794;
						assign node794 = (inp[11]) ? node800 : node795;
							assign node795 = (inp[8]) ? 14'b00000000000000 : node796;
								assign node796 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node800 = (inp[7]) ? 14'b00000000000000 : node801;
								assign node801 = (inp[0]) ? 14'b00000000000000 : node802;
									assign node802 = (inp[13]) ? node804 : 14'b00000000000000;
										assign node804 = (inp[2]) ? 14'b00000000000000 : node805;
											assign node805 = (inp[8]) ? node807 : 14'b00000000000000;
												assign node807 = (inp[9]) ? 14'b00000000000000 : node808;
													assign node808 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
						assign node815 = (inp[13]) ? node837 : node816;
							assign node816 = (inp[11]) ? node832 : node817;
								assign node817 = (inp[8]) ? node829 : node818;
									assign node818 = (inp[2]) ? 14'b00000000000000 : node819;
										assign node819 = (inp[0]) ? 14'b00000000000000 : node820;
											assign node820 = (inp[9]) ? 14'b00000000000000 : node821;
												assign node821 = (inp[7]) ? 14'b00000000000000 : node822;
													assign node822 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
									assign node829 = (inp[9]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node832 = (inp[9]) ? 14'b00000000000000 : node833;
									assign node833 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000101;
							assign node837 = (inp[11]) ? node853 : node838;
								assign node838 = (inp[9]) ? node850 : node839;
									assign node839 = (inp[8]) ? 14'b00000000000000 : node840;
										assign node840 = (inp[0]) ? 14'b00000000000000 : node841;
											assign node841 = (inp[7]) ? 14'b00000000000000 : node842;
												assign node842 = (inp[2]) ? 14'b00000000000000 : node843;
													assign node843 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
									assign node850 = (inp[8]) ? 14'b00100100001101 : 14'b00000000000000;
								assign node853 = (inp[9]) ? node857 : node854;
									assign node854 = (inp[8]) ? 14'b10000100001000 : 14'b10010101111110;
									assign node857 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
			assign node860 = (inp[9]) ? node1174 : node861;
				assign node861 = (inp[3]) ? node1037 : node862;
					assign node862 = (inp[6]) ? node990 : node863;
						assign node863 = (inp[8]) ? node909 : node864;
							assign node864 = (inp[11]) ? node876 : node865;
								assign node865 = (inp[12]) ? node869 : node866;
									assign node866 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node869 = (inp[13]) ? 14'b00000000011101 : node870;
										assign node870 = (inp[0]) ? node872 : 14'b00000000000000;
											assign node872 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node876 = (inp[0]) ? node878 : 14'b00000000000000;
									assign node878 = (inp[4]) ? 14'b00000000000000 : node879;
										assign node879 = (inp[13]) ? node893 : node880;
											assign node880 = (inp[12]) ? node888 : node881;
												assign node881 = (inp[2]) ? 14'b01001000000101 : node882;
													assign node882 = (inp[7]) ? node884 : 14'b00000000000000;
														assign node884 = (inp[5]) ? 14'b00000000000000 : 14'b01100000001010;
												assign node888 = (inp[5]) ? 14'b00000000000000 : node889;
													assign node889 = (inp[2]) ? 14'b00000000000000 : 14'b00001000000101;
											assign node893 = (inp[5]) ? node903 : node894;
												assign node894 = (inp[2]) ? node900 : node895;
													assign node895 = (inp[12]) ? 14'b10000000001111 : node896;
														assign node896 = (inp[7]) ? 14'b10000100001101 : 14'b00000000000000;
													assign node900 = (inp[12]) ? 14'b00000000000000 : 14'b00000000011100;
												assign node903 = (inp[12]) ? 14'b00000000000000 : node904;
													assign node904 = (inp[2]) ? 14'b00000000011100 : 14'b00000000000000;
							assign node909 = (inp[11]) ? node959 : node910;
								assign node910 = (inp[12]) ? node940 : node911;
									assign node911 = (inp[13]) ? node931 : node912;
										assign node912 = (inp[0]) ? node918 : node913;
											assign node913 = (inp[4]) ? 14'b00100000000011 : node914;
												assign node914 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node918 = (inp[4]) ? node926 : node919;
												assign node919 = (inp[2]) ? 14'b00100000000011 : node920;
													assign node920 = (inp[7]) ? node922 : 14'b00000000000000;
														assign node922 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
												assign node926 = (inp[5]) ? node928 : 14'b00000000000000;
													assign node928 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node931 = (inp[0]) ? node933 : 14'b00000000000000;
											assign node933 = (inp[2]) ? 14'b00000000000000 : node934;
												assign node934 = (inp[5]) ? 14'b00000000000000 : node935;
													assign node935 = (inp[4]) ? 14'b00000000000000 : 14'b10110111101111;
									assign node940 = (inp[13]) ? node952 : node941;
										assign node941 = (inp[2]) ? 14'b00000000000000 : node942;
											assign node942 = (inp[0]) ? node946 : node943;
												assign node943 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
												assign node946 = (inp[5]) ? 14'b00000000000000 : node947;
													assign node947 = (inp[4]) ? 14'b00000000000000 : 14'b10000100011000;
										assign node952 = (inp[0]) ? 14'b00001000000100 : node953;
											assign node953 = (inp[2]) ? 14'b00001000000100 : node954;
												assign node954 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
								assign node959 = (inp[13]) ? node981 : node960;
									assign node960 = (inp[12]) ? 14'b00000000000000 : node961;
										assign node961 = (inp[4]) ? node973 : node962;
											assign node962 = (inp[2]) ? node970 : node963;
												assign node963 = (inp[0]) ? node965 : 14'b10000001001101;
													assign node965 = (inp[7]) ? node967 : 14'b00000000000000;
														assign node967 = (inp[5]) ? 14'b00000000000000 : 14'b10100000001101;
												assign node970 = (inp[0]) ? 14'b10010000001101 : 14'b00000000000000;
											assign node973 = (inp[0]) ? node977 : node974;
												assign node974 = (inp[2]) ? 14'b10000100001101 : 14'b10000010001101;
												assign node977 = (inp[5]) ? 14'b10000000011101 : 14'b00000000000000;
									assign node981 = (inp[12]) ? 14'b10000100001000 : node982;
										assign node982 = (inp[0]) ? 14'b10100100011000 : node983;
											assign node983 = (inp[2]) ? node985 : 14'b10000000001010;
												assign node985 = (inp[4]) ? 14'b10100100011000 : 14'b00000000000000;
						assign node990 = (inp[11]) ? node1020 : node991;
							assign node991 = (inp[12]) ? node997 : node992;
								assign node992 = (inp[13]) ? 14'b00000000000000 : node993;
									assign node993 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node997 = (inp[13]) ? node1009 : node998;
									assign node998 = (inp[8]) ? 14'b00000000000000 : node999;
										assign node999 = (inp[0]) ? 14'b00000000000000 : node1000;
											assign node1000 = (inp[2]) ? 14'b00000000000000 : node1001;
												assign node1001 = (inp[5]) ? node1003 : 14'b00000000000000;
													assign node1003 = (inp[7]) ? 14'b00000100001101 : 14'b00000000000000;
									assign node1009 = (inp[8]) ? 14'b00000100001110 : node1010;
										assign node1010 = (inp[5]) ? node1012 : 14'b00000000000000;
											assign node1012 = (inp[0]) ? 14'b00000000000000 : node1013;
												assign node1013 = (inp[2]) ? 14'b00000000000000 : node1014;
													assign node1014 = (inp[7]) ? 14'b00000000011100 : 14'b00000000000000;
							assign node1020 = (inp[12]) ? node1022 : 14'b00000000000000;
								assign node1022 = (inp[8]) ? node1034 : node1023;
									assign node1023 = (inp[5]) ? node1025 : 14'b00000000000000;
										assign node1025 = (inp[7]) ? node1027 : 14'b00000000000000;
											assign node1027 = (inp[0]) ? 14'b00000000000000 : node1028;
												assign node1028 = (inp[2]) ? 14'b00000000000000 : node1029;
													assign node1029 = (inp[13]) ? 14'b01001000000101 : 14'b01100000000010;
									assign node1034 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node1037 = (inp[0]) ? node1143 : node1038;
						assign node1038 = (inp[2]) ? node1112 : node1039;
							assign node1039 = (inp[6]) ? node1097 : node1040;
								assign node1040 = (inp[11]) ? node1070 : node1041;
									assign node1041 = (inp[13]) ? node1055 : node1042;
										assign node1042 = (inp[8]) ? node1046 : node1043;
											assign node1043 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1046 = (inp[7]) ? node1050 : node1047;
												assign node1047 = (inp[12]) ? 14'b00000000011100 : 14'b00000000000000;
												assign node1050 = (inp[12]) ? 14'b00000000000000 : node1051;
													assign node1051 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
										assign node1055 = (inp[12]) ? node1065 : node1056;
											assign node1056 = (inp[7]) ? node1060 : node1057;
												assign node1057 = (inp[8]) ? 14'b00001000001001 : 14'b00000000000000;
												assign node1060 = (inp[8]) ? 14'b00000000000000 : node1061;
													assign node1061 = (inp[5]) ? 14'b00001000000100 : 14'b00000000000000;
											assign node1065 = (inp[8]) ? 14'b00000000000000 : node1066;
												assign node1066 = (inp[7]) ? 14'b01100000001010 : 14'b00000000000000;
									assign node1070 = (inp[8]) ? node1082 : node1071;
										assign node1071 = (inp[12]) ? node1077 : node1072;
											assign node1072 = (inp[5]) ? 14'b00100000000011 : node1073;
												assign node1073 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node1077 = (inp[13]) ? 14'b00000000000000 : node1078;
												assign node1078 = (inp[7]) ? 14'b00100100001101 : 14'b00000000000000;
										assign node1082 = (inp[13]) ? node1088 : node1083;
											assign node1083 = (inp[12]) ? 14'b00000000000000 : node1084;
												assign node1084 = (inp[7]) ? 14'b00000000000000 : 14'b00100000001010;
											assign node1088 = (inp[7]) ? node1094 : node1089;
												assign node1089 = (inp[12]) ? 14'b10000100001000 : node1090;
													assign node1090 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
												assign node1094 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1097 = (inp[12]) ? node1105 : node1098;
									assign node1098 = (inp[8]) ? 14'b00000000000000 : node1099;
										assign node1099 = (inp[13]) ? 14'b00000000000000 : node1100;
											assign node1100 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node1105 = (inp[8]) ? node1107 : 14'b00000000000000;
										assign node1107 = (inp[13]) ? node1109 : 14'b00000000000000;
											assign node1109 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1112 = (inp[6]) ? node1128 : node1113;
								assign node1113 = (inp[12]) ? node1121 : node1114;
									assign node1114 = (inp[11]) ? 14'b00000000000000 : node1115;
										assign node1115 = (inp[13]) ? 14'b00000000000000 : node1116;
											assign node1116 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node1121 = (inp[11]) ? node1123 : 14'b00000000000000;
										assign node1123 = (inp[13]) ? node1125 : 14'b00000000000000;
											assign node1125 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1128 = (inp[12]) ? node1136 : node1129;
									assign node1129 = (inp[13]) ? 14'b00000000000000 : node1130;
										assign node1130 = (inp[8]) ? 14'b00000000000000 : node1131;
											assign node1131 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node1136 = (inp[11]) ? node1138 : 14'b00000000000000;
										assign node1138 = (inp[8]) ? node1140 : 14'b00000000000000;
											assign node1140 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node1143 = (inp[5]) ? node1159 : node1144;
							assign node1144 = (inp[8]) ? node1152 : node1145;
								assign node1145 = (inp[13]) ? 14'b00000000000000 : node1146;
									assign node1146 = (inp[12]) ? 14'b00000000000000 : node1147;
										assign node1147 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node1152 = (inp[13]) ? node1154 : 14'b00000000000000;
									assign node1154 = (inp[12]) ? node1156 : 14'b00000000000000;
										assign node1156 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1159 = (inp[13]) ? node1167 : node1160;
								assign node1160 = (inp[12]) ? 14'b00000000000000 : node1161;
									assign node1161 = (inp[11]) ? 14'b00000000000000 : node1162;
										assign node1162 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node1167 = (inp[11]) ? node1169 : 14'b00000000000000;
									assign node1169 = (inp[12]) ? node1171 : 14'b00000000000000;
										assign node1171 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node1174 = (inp[3]) ? node1350 : node1175;
					assign node1175 = (inp[7]) ? node1317 : node1176;
						assign node1176 = (inp[4]) ? node1192 : node1177;
							assign node1177 = (inp[13]) ? node1185 : node1178;
								assign node1178 = (inp[12]) ? 14'b00000000000000 : node1179;
									assign node1179 = (inp[11]) ? 14'b00000000000000 : node1180;
										assign node1180 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node1185 = (inp[8]) ? node1187 : 14'b00000000000000;
									assign node1187 = (inp[12]) ? node1189 : 14'b00000000000000;
										assign node1189 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1192 = (inp[2]) ? node1224 : node1193;
								assign node1193 = (inp[5]) ? node1209 : node1194;
									assign node1194 = (inp[12]) ? node1202 : node1195;
										assign node1195 = (inp[8]) ? 14'b00000000000000 : node1196;
											assign node1196 = (inp[11]) ? 14'b00000000000000 : node1197;
												assign node1197 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1202 = (inp[11]) ? node1204 : 14'b00000000000000;
											assign node1204 = (inp[13]) ? node1206 : 14'b00000000000000;
												assign node1206 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1209 = (inp[8]) ? node1217 : node1210;
										assign node1210 = (inp[13]) ? 14'b00000000000000 : node1211;
											assign node1211 = (inp[11]) ? 14'b00000000000000 : node1212;
												assign node1212 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1217 = (inp[12]) ? node1219 : 14'b00000000000000;
											assign node1219 = (inp[13]) ? node1221 : 14'b00000000000000;
												assign node1221 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1224 = (inp[5]) ? node1272 : node1225;
									assign node1225 = (inp[6]) ? node1241 : node1226;
										assign node1226 = (inp[12]) ? node1234 : node1227;
											assign node1227 = (inp[11]) ? 14'b00000000000000 : node1228;
												assign node1228 = (inp[13]) ? 14'b00000000000000 : node1229;
													assign node1229 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1234 = (inp[11]) ? node1236 : 14'b00000000000000;
												assign node1236 = (inp[8]) ? node1238 : 14'b00000000000000;
													assign node1238 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node1241 = (inp[0]) ? node1257 : node1242;
											assign node1242 = (inp[12]) ? node1250 : node1243;
												assign node1243 = (inp[8]) ? 14'b00000000000000 : node1244;
													assign node1244 = (inp[13]) ? 14'b00000000000000 : node1245;
														assign node1245 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
												assign node1250 = (inp[11]) ? node1252 : 14'b00000000000000;
													assign node1252 = (inp[8]) ? node1254 : 14'b00000000000000;
														assign node1254 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
											assign node1257 = (inp[11]) ? node1265 : node1258;
												assign node1258 = (inp[13]) ? 14'b00000000000000 : node1259;
													assign node1259 = (inp[12]) ? 14'b00000000000000 : node1260;
														assign node1260 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
												assign node1265 = (inp[8]) ? node1267 : 14'b00000000000000;
													assign node1267 = (inp[12]) ? node1269 : 14'b00000000000000;
														assign node1269 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1272 = (inp[6]) ? node1288 : node1273;
										assign node1273 = (inp[12]) ? node1281 : node1274;
											assign node1274 = (inp[8]) ? 14'b00000000000000 : node1275;
												assign node1275 = (inp[11]) ? 14'b00000000000000 : node1276;
													assign node1276 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1281 = (inp[13]) ? node1283 : 14'b00000000000000;
												assign node1283 = (inp[11]) ? node1285 : 14'b00000000000000;
													assign node1285 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node1288 = (inp[0]) ? node1304 : node1289;
											assign node1289 = (inp[13]) ? node1297 : node1290;
												assign node1290 = (inp[12]) ? 14'b00000000000000 : node1291;
													assign node1291 = (inp[8]) ? 14'b00000000000000 : node1292;
														assign node1292 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
												assign node1297 = (inp[11]) ? node1299 : 14'b00000000000000;
													assign node1299 = (inp[8]) ? node1301 : 14'b00000000000000;
														assign node1301 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
											assign node1304 = (inp[13]) ? node1310 : node1305;
												assign node1305 = (inp[11]) ? 14'b00000000000000 : node1306;
													assign node1306 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
												assign node1310 = (inp[12]) ? node1312 : 14'b00000000000000;
													assign node1312 = (inp[11]) ? node1314 : 14'b00000000000000;
														assign node1314 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node1317 = (inp[8]) ? node1343 : node1318;
							assign node1318 = (inp[13]) ? node1332 : node1319;
								assign node1319 = (inp[11]) ? node1323 : node1320;
									assign node1320 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node1323 = (inp[0]) ? 14'b00000000000000 : node1324;
										assign node1324 = (inp[6]) ? 14'b00000000000000 : node1325;
											assign node1325 = (inp[2]) ? 14'b00000000000000 : node1326;
												assign node1326 = (inp[12]) ? 14'b00100100001101 : 14'b00000000000000;
								assign node1332 = (inp[2]) ? 14'b00000000000000 : node1333;
									assign node1333 = (inp[6]) ? 14'b00000000000000 : node1334;
										assign node1334 = (inp[11]) ? 14'b00000000000000 : node1335;
											assign node1335 = (inp[0]) ? 14'b00000000000000 : node1336;
												assign node1336 = (inp[12]) ? 14'b01100000001010 : 14'b00001000000100;
							assign node1343 = (inp[11]) ? node1345 : 14'b00000000000000;
								assign node1345 = (inp[13]) ? node1347 : 14'b00000000000000;
									assign node1347 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node1350 = (inp[6]) ? node1532 : node1351;
						assign node1351 = (inp[0]) ? node1453 : node1352;
							assign node1352 = (inp[2]) ? node1406 : node1353;
								assign node1353 = (inp[11]) ? node1377 : node1354;
									assign node1354 = (inp[8]) ? node1366 : node1355;
										assign node1355 = (inp[13]) ? node1359 : node1356;
											assign node1356 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1359 = (inp[12]) ? node1363 : node1360;
												assign node1360 = (inp[7]) ? 14'b00001000000100 : 14'b00000000000000;
												assign node1363 = (inp[7]) ? 14'b01100000001010 : 14'b00000000000000;
										assign node1366 = (inp[7]) ? 14'b00000000000000 : node1367;
											assign node1367 = (inp[12]) ? node1371 : node1368;
												assign node1368 = (inp[13]) ? 14'b00001000001001 : 14'b00000000000000;
												assign node1371 = (inp[13]) ? node1373 : 14'b00000000011100;
													assign node1373 = (inp[5]) ? 14'b00000000011101 : 14'b00000000000000;
									assign node1377 = (inp[8]) ? node1391 : node1378;
										assign node1378 = (inp[13]) ? node1386 : node1379;
											assign node1379 = (inp[12]) ? node1383 : node1380;
												assign node1380 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
												assign node1383 = (inp[7]) ? 14'b00100100001101 : 14'b00000000000000;
											assign node1386 = (inp[7]) ? 14'b00000000000000 : node1387;
												assign node1387 = (inp[12]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node1391 = (inp[13]) ? node1397 : node1392;
											assign node1392 = (inp[7]) ? 14'b00000000000000 : node1393;
												assign node1393 = (inp[12]) ? 14'b00000000000000 : 14'b00100000001010;
											assign node1397 = (inp[7]) ? node1403 : node1398;
												assign node1398 = (inp[12]) ? 14'b10000100001000 : node1399;
													assign node1399 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
												assign node1403 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1406 = (inp[5]) ? node1422 : node1407;
									assign node1407 = (inp[11]) ? node1415 : node1408;
										assign node1408 = (inp[13]) ? 14'b00000000000000 : node1409;
											assign node1409 = (inp[12]) ? 14'b00000000000000 : node1410;
												assign node1410 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1415 = (inp[12]) ? node1417 : 14'b00000000000000;
											assign node1417 = (inp[13]) ? node1419 : 14'b00000000000000;
												assign node1419 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1422 = (inp[4]) ? node1438 : node1423;
										assign node1423 = (inp[11]) ? node1431 : node1424;
											assign node1424 = (inp[12]) ? 14'b00000000000000 : node1425;
												assign node1425 = (inp[8]) ? 14'b00000000000000 : node1426;
													assign node1426 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1431 = (inp[13]) ? node1433 : 14'b00000000000000;
												assign node1433 = (inp[12]) ? node1435 : 14'b00000000000000;
													assign node1435 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node1438 = (inp[12]) ? node1446 : node1439;
											assign node1439 = (inp[11]) ? 14'b00000000000000 : node1440;
												assign node1440 = (inp[13]) ? 14'b00000000000000 : node1441;
													assign node1441 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1446 = (inp[8]) ? node1448 : 14'b00000000000000;
												assign node1448 = (inp[13]) ? node1450 : 14'b00000000000000;
													assign node1450 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1453 = (inp[4]) ? node1501 : node1454;
								assign node1454 = (inp[2]) ? node1470 : node1455;
									assign node1455 = (inp[8]) ? node1463 : node1456;
										assign node1456 = (inp[13]) ? 14'b00000000000000 : node1457;
											assign node1457 = (inp[11]) ? 14'b00000000000000 : node1458;
												assign node1458 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1463 = (inp[11]) ? node1465 : 14'b00000000000000;
											assign node1465 = (inp[12]) ? node1467 : 14'b00000000000000;
												assign node1467 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1470 = (inp[5]) ? node1486 : node1471;
										assign node1471 = (inp[12]) ? node1479 : node1472;
											assign node1472 = (inp[11]) ? 14'b00000000000000 : node1473;
												assign node1473 = (inp[13]) ? 14'b00000000000000 : node1474;
													assign node1474 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1479 = (inp[11]) ? node1481 : 14'b00000000000000;
												assign node1481 = (inp[13]) ? node1483 : 14'b00000000000000;
													assign node1483 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node1486 = (inp[12]) ? node1494 : node1487;
											assign node1487 = (inp[11]) ? 14'b00000000000000 : node1488;
												assign node1488 = (inp[13]) ? 14'b00000000000000 : node1489;
													assign node1489 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1494 = (inp[13]) ? node1496 : 14'b00000000000000;
												assign node1496 = (inp[8]) ? node1498 : 14'b00000000000000;
													assign node1498 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1501 = (inp[5]) ? node1517 : node1502;
									assign node1502 = (inp[12]) ? node1510 : node1503;
										assign node1503 = (inp[13]) ? 14'b00000000000000 : node1504;
											assign node1504 = (inp[11]) ? 14'b00000000000000 : node1505;
												assign node1505 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1510 = (inp[13]) ? node1512 : 14'b00000000000000;
											assign node1512 = (inp[11]) ? node1514 : 14'b00000000000000;
												assign node1514 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1517 = (inp[8]) ? node1525 : node1518;
										assign node1518 = (inp[11]) ? 14'b00000000000000 : node1519;
											assign node1519 = (inp[12]) ? 14'b00000000000000 : node1520;
												assign node1520 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1525 = (inp[11]) ? node1527 : 14'b00000000000000;
											assign node1527 = (inp[13]) ? node1529 : 14'b00000000000000;
												assign node1529 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node1532 = (inp[7]) ? node1562 : node1533;
							assign node1533 = (inp[12]) ? node1541 : node1534;
								assign node1534 = (inp[8]) ? 14'b00000000000000 : node1535;
									assign node1535 = (inp[11]) ? 14'b00000000000000 : node1536;
										assign node1536 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node1541 = (inp[5]) ? node1549 : node1542;
									assign node1542 = (inp[8]) ? node1544 : 14'b00000000000000;
										assign node1544 = (inp[11]) ? node1546 : 14'b00000000000000;
											assign node1546 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1549 = (inp[8]) ? node1557 : node1550;
										assign node1550 = (inp[13]) ? node1554 : node1551;
											assign node1551 = (inp[11]) ? 14'b00000100001111 : 14'b00001000001100;
											assign node1554 = (inp[11]) ? 14'b10100100001000 : 14'b10100000001000;
										assign node1557 = (inp[11]) ? node1559 : 14'b00000000000000;
											assign node1559 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1562 = (inp[12]) ? node1618 : node1563;
								assign node1563 = (inp[11]) ? node1591 : node1564;
									assign node1564 = (inp[13]) ? node1576 : node1565;
										assign node1565 = (inp[8]) ? node1567 : 14'b10000100001000;
											assign node1567 = (inp[5]) ? 14'b10100000001000 : node1568;
												assign node1568 = (inp[0]) ? 14'b00000000000000 : node1569;
													assign node1569 = (inp[4]) ? node1571 : 14'b10010010001101;
														assign node1571 = (inp[2]) ? 14'b00000000000000 : 14'b00100000001010;
										assign node1576 = (inp[0]) ? 14'b00000000000000 : node1577;
											assign node1577 = (inp[5]) ? 14'b00000000000000 : node1578;
												assign node1578 = (inp[2]) ? node1584 : node1579;
													assign node1579 = (inp[8]) ? node1581 : 14'b00000000011101;
														assign node1581 = (inp[4]) ? 14'b10000100101000 : 14'b10000100111000;
													assign node1584 = (inp[8]) ? node1586 : 14'b00000000000000;
														assign node1586 = (inp[4]) ? 14'b00000000000000 : 14'b10100000001000;
									assign node1591 = (inp[5]) ? node1609 : node1592;
										assign node1592 = (inp[8]) ? node1606 : node1593;
											assign node1593 = (inp[13]) ? node1599 : node1594;
												assign node1594 = (inp[0]) ? 14'b00000100001111 : node1595;
													assign node1595 = (inp[2]) ? 14'b00000100001111 : 14'b00100000000011;
												assign node1599 = (inp[0]) ? 14'b01000100000010 : node1600;
													assign node1600 = (inp[2]) ? node1602 : 14'b00001000001001;
														assign node1602 = (inp[4]) ? 14'b01000100000010 : 14'b01100000000010;
											assign node1606 = (inp[13]) ? 14'b00100100001101 : 14'b01001000000100;
										assign node1609 = (inp[8]) ? 14'b00000000000000 : node1610;
											assign node1610 = (inp[13]) ? 14'b10100101111111 : node1611;
												assign node1611 = (inp[0]) ? node1613 : 14'b00000000000000;
													assign node1613 = (inp[4]) ? 14'b00100000000011 : 14'b00000000000000;
								assign node1618 = (inp[8]) ? node1620 : 14'b00000000000000;
									assign node1620 = (inp[13]) ? node1626 : node1621;
										assign node1621 = (inp[5]) ? node1623 : 14'b00000000000000;
											assign node1623 = (inp[11]) ? 14'b00000000000000 : 14'b01100000000110;
										assign node1626 = (inp[11]) ? 14'b10000100001000 : node1627;
											assign node1627 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;

endmodule