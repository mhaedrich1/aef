module dtc_split05_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node14;
	wire [16-1:0] node16;
	wire [16-1:0] node19;
	wire [16-1:0] node20;
	wire [16-1:0] node21;
	wire [16-1:0] node22;
	wire [16-1:0] node25;
	wire [16-1:0] node26;
	wire [16-1:0] node27;
	wire [16-1:0] node31;
	wire [16-1:0] node34;
	wire [16-1:0] node36;
	wire [16-1:0] node39;
	wire [16-1:0] node41;
	wire [16-1:0] node42;
	wire [16-1:0] node46;
	wire [16-1:0] node47;
	wire [16-1:0] node48;
	wire [16-1:0] node49;
	wire [16-1:0] node50;
	wire [16-1:0] node51;
	wire [16-1:0] node55;
	wire [16-1:0] node57;
	wire [16-1:0] node61;
	wire [16-1:0] node62;
	wire [16-1:0] node63;
	wire [16-1:0] node66;
	wire [16-1:0] node70;
	wire [16-1:0] node71;
	wire [16-1:0] node72;
	wire [16-1:0] node73;
	wire [16-1:0] node74;
	wire [16-1:0] node75;
	wire [16-1:0] node80;
	wire [16-1:0] node84;
	wire [16-1:0] node85;
	wire [16-1:0] node87;
	wire [16-1:0] node90;
	wire [16-1:0] node92;
	wire [16-1:0] node93;
	wire [16-1:0] node95;
	wire [16-1:0] node99;
	wire [16-1:0] node100;
	wire [16-1:0] node101;
	wire [16-1:0] node102;
	wire [16-1:0] node103;
	wire [16-1:0] node106;
	wire [16-1:0] node107;
	wire [16-1:0] node111;
	wire [16-1:0] node112;
	wire [16-1:0] node113;
	wire [16-1:0] node116;
	wire [16-1:0] node120;
	wire [16-1:0] node121;
	wire [16-1:0] node123;
	wire [16-1:0] node126;
	wire [16-1:0] node129;
	wire [16-1:0] node130;
	wire [16-1:0] node131;
	wire [16-1:0] node132;
	wire [16-1:0] node134;
	wire [16-1:0] node137;
	wire [16-1:0] node138;
	wire [16-1:0] node140;
	wire [16-1:0] node144;
	wire [16-1:0] node145;
	wire [16-1:0] node146;
	wire [16-1:0] node149;
	wire [16-1:0] node152;
	wire [16-1:0] node155;
	wire [16-1:0] node156;
	wire [16-1:0] node157;
	wire [16-1:0] node159;
	wire [16-1:0] node162;
	wire [16-1:0] node163;
	wire [16-1:0] node167;
	wire [16-1:0] node168;
	wire [16-1:0] node169;
	wire [16-1:0] node171;
	wire [16-1:0] node175;
	wire [16-1:0] node176;
	wire [16-1:0] node179;
	wire [16-1:0] node182;
	wire [16-1:0] node183;
	wire [16-1:0] node184;
	wire [16-1:0] node185;
	wire [16-1:0] node186;
	wire [16-1:0] node187;
	wire [16-1:0] node191;
	wire [16-1:0] node193;
	wire [16-1:0] node194;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node200;
	wire [16-1:0] node202;
	wire [16-1:0] node205;
	wire [16-1:0] node208;
	wire [16-1:0] node211;
	wire [16-1:0] node212;
	wire [16-1:0] node213;
	wire [16-1:0] node215;
	wire [16-1:0] node218;
	wire [16-1:0] node219;
	wire [16-1:0] node222;
	wire [16-1:0] node224;
	wire [16-1:0] node226;
	wire [16-1:0] node229;
	wire [16-1:0] node230;
	wire [16-1:0] node231;
	wire [16-1:0] node234;
	wire [16-1:0] node237;
	wire [16-1:0] node238;
	wire [16-1:0] node240;
	wire [16-1:0] node244;
	wire [16-1:0] node245;
	wire [16-1:0] node246;
	wire [16-1:0] node247;
	wire [16-1:0] node248;
	wire [16-1:0] node249;
	wire [16-1:0] node254;
	wire [16-1:0] node256;
	wire [16-1:0] node259;
	wire [16-1:0] node260;
	wire [16-1:0] node261;
	wire [16-1:0] node262;
	wire [16-1:0] node264;
	wire [16-1:0] node269;
	wire [16-1:0] node270;
	wire [16-1:0] node271;
	wire [16-1:0] node273;
	wire [16-1:0] node276;
	wire [16-1:0] node278;
	wire [16-1:0] node280;
	wire [16-1:0] node281;
	wire [16-1:0] node285;
	wire [16-1:0] node287;
	wire [16-1:0] node288;
	wire [16-1:0] node289;
	wire [16-1:0] node294;
	wire [16-1:0] node295;
	wire [16-1:0] node298;
	wire [16-1:0] node299;
	wire [16-1:0] node300;
	wire [16-1:0] node301;
	wire [16-1:0] node305;
	wire [16-1:0] node306;
	wire [16-1:0] node309;
	wire [16-1:0] node312;
	wire [16-1:0] node313;
	wire [16-1:0] node316;
	wire [16-1:0] node317;
	wire [16-1:0] node319;
	wire [16-1:0] node323;
	wire [16-1:0] node324;
	wire [16-1:0] node325;
	wire [16-1:0] node326;
	wire [16-1:0] node327;
	wire [16-1:0] node328;
	wire [16-1:0] node329;
	wire [16-1:0] node331;
	wire [16-1:0] node334;
	wire [16-1:0] node337;
	wire [16-1:0] node338;
	wire [16-1:0] node340;
	wire [16-1:0] node344;
	wire [16-1:0] node345;
	wire [16-1:0] node346;
	wire [16-1:0] node347;
	wire [16-1:0] node349;
	wire [16-1:0] node353;
	wire [16-1:0] node355;
	wire [16-1:0] node358;
	wire [16-1:0] node361;
	wire [16-1:0] node362;
	wire [16-1:0] node363;
	wire [16-1:0] node366;
	wire [16-1:0] node367;
	wire [16-1:0] node368;
	wire [16-1:0] node372;
	wire [16-1:0] node375;
	wire [16-1:0] node376;
	wire [16-1:0] node377;
	wire [16-1:0] node378;
	wire [16-1:0] node382;
	wire [16-1:0] node385;
	wire [16-1:0] node386;
	wire [16-1:0] node389;
	wire [16-1:0] node391;
	wire [16-1:0] node394;
	wire [16-1:0] node395;
	wire [16-1:0] node396;
	wire [16-1:0] node397;
	wire [16-1:0] node398;
	wire [16-1:0] node400;
	wire [16-1:0] node403;
	wire [16-1:0] node404;
	wire [16-1:0] node408;
	wire [16-1:0] node410;
	wire [16-1:0] node413;
	wire [16-1:0] node414;
	wire [16-1:0] node415;
	wire [16-1:0] node417;
	wire [16-1:0] node420;
	wire [16-1:0] node421;
	wire [16-1:0] node425;
	wire [16-1:0] node427;
	wire [16-1:0] node428;
	wire [16-1:0] node429;
	wire [16-1:0] node434;
	wire [16-1:0] node435;
	wire [16-1:0] node436;
	wire [16-1:0] node437;
	wire [16-1:0] node440;
	wire [16-1:0] node441;
	wire [16-1:0] node442;
	wire [16-1:0] node447;
	wire [16-1:0] node449;
	wire [16-1:0] node450;
	wire [16-1:0] node453;
	wire [16-1:0] node456;
	wire [16-1:0] node457;
	wire [16-1:0] node458;
	wire [16-1:0] node461;
	wire [16-1:0] node464;
	wire [16-1:0] node465;
	wire [16-1:0] node466;
	wire [16-1:0] node468;
	wire [16-1:0] node472;
	wire [16-1:0] node474;
	wire [16-1:0] node477;
	wire [16-1:0] node478;
	wire [16-1:0] node479;
	wire [16-1:0] node480;
	wire [16-1:0] node481;
	wire [16-1:0] node482;
	wire [16-1:0] node484;
	wire [16-1:0] node488;
	wire [16-1:0] node489;
	wire [16-1:0] node493;
	wire [16-1:0] node494;
	wire [16-1:0] node495;
	wire [16-1:0] node496;
	wire [16-1:0] node501;
	wire [16-1:0] node502;
	wire [16-1:0] node505;
	wire [16-1:0] node508;
	wire [16-1:0] node509;
	wire [16-1:0] node510;
	wire [16-1:0] node511;
	wire [16-1:0] node513;
	wire [16-1:0] node516;
	wire [16-1:0] node518;
	wire [16-1:0] node521;
	wire [16-1:0] node524;
	wire [16-1:0] node525;
	wire [16-1:0] node526;
	wire [16-1:0] node527;
	wire [16-1:0] node531;
	wire [16-1:0] node534;
	wire [16-1:0] node535;
	wire [16-1:0] node539;
	wire [16-1:0] node540;
	wire [16-1:0] node541;
	wire [16-1:0] node542;
	wire [16-1:0] node543;
	wire [16-1:0] node545;
	wire [16-1:0] node549;
	wire [16-1:0] node550;
	wire [16-1:0] node553;
	wire [16-1:0] node554;
	wire [16-1:0] node558;
	wire [16-1:0] node559;
	wire [16-1:0] node560;
	wire [16-1:0] node563;
	wire [16-1:0] node566;
	wire [16-1:0] node567;
	wire [16-1:0] node568;
	wire [16-1:0] node571;
	wire [16-1:0] node574;
	wire [16-1:0] node577;
	wire [16-1:0] node578;
	wire [16-1:0] node579;
	wire [16-1:0] node580;
	wire [16-1:0] node582;
	wire [16-1:0] node585;
	wire [16-1:0] node586;
	wire [16-1:0] node590;
	wire [16-1:0] node591;
	wire [16-1:0] node594;
	wire [16-1:0] node597;
	wire [16-1:0] node598;
	wire [16-1:0] node600;
	wire [16-1:0] node602;
	wire [16-1:0] node605;
	wire [16-1:0] node606;
	wire [16-1:0] node609;
	wire [16-1:0] node611;
	wire [16-1:0] node614;
	wire [16-1:0] node615;
	wire [16-1:0] node616;
	wire [16-1:0] node617;
	wire [16-1:0] node618;
	wire [16-1:0] node619;
	wire [16-1:0] node620;
	wire [16-1:0] node622;
	wire [16-1:0] node623;
	wire [16-1:0] node625;
	wire [16-1:0] node629;
	wire [16-1:0] node630;
	wire [16-1:0] node631;
	wire [16-1:0] node635;
	wire [16-1:0] node638;
	wire [16-1:0] node639;
	wire [16-1:0] node640;
	wire [16-1:0] node644;
	wire [16-1:0] node646;
	wire [16-1:0] node647;
	wire [16-1:0] node651;
	wire [16-1:0] node652;
	wire [16-1:0] node653;
	wire [16-1:0] node654;
	wire [16-1:0] node656;
	wire [16-1:0] node659;
	wire [16-1:0] node660;
	wire [16-1:0] node663;
	wire [16-1:0] node667;
	wire [16-1:0] node668;
	wire [16-1:0] node669;
	wire [16-1:0] node672;
	wire [16-1:0] node675;
	wire [16-1:0] node676;
	wire [16-1:0] node680;
	wire [16-1:0] node681;
	wire [16-1:0] node682;
	wire [16-1:0] node683;
	wire [16-1:0] node684;
	wire [16-1:0] node686;
	wire [16-1:0] node688;
	wire [16-1:0] node691;
	wire [16-1:0] node693;
	wire [16-1:0] node696;
	wire [16-1:0] node697;
	wire [16-1:0] node698;
	wire [16-1:0] node701;
	wire [16-1:0] node703;
	wire [16-1:0] node704;
	wire [16-1:0] node708;
	wire [16-1:0] node710;
	wire [16-1:0] node713;
	wire [16-1:0] node714;
	wire [16-1:0] node715;
	wire [16-1:0] node719;
	wire [16-1:0] node720;
	wire [16-1:0] node723;
	wire [16-1:0] node724;
	wire [16-1:0] node727;
	wire [16-1:0] node730;
	wire [16-1:0] node731;
	wire [16-1:0] node732;
	wire [16-1:0] node733;
	wire [16-1:0] node734;
	wire [16-1:0] node739;
	wire [16-1:0] node741;
	wire [16-1:0] node742;
	wire [16-1:0] node744;
	wire [16-1:0] node748;
	wire [16-1:0] node749;
	wire [16-1:0] node750;
	wire [16-1:0] node752;
	wire [16-1:0] node756;
	wire [16-1:0] node757;
	wire [16-1:0] node758;
	wire [16-1:0] node760;
	wire [16-1:0] node764;
	wire [16-1:0] node767;
	wire [16-1:0] node768;
	wire [16-1:0] node769;
	wire [16-1:0] node770;
	wire [16-1:0] node771;
	wire [16-1:0] node772;
	wire [16-1:0] node773;
	wire [16-1:0] node776;
	wire [16-1:0] node780;
	wire [16-1:0] node781;
	wire [16-1:0] node783;
	wire [16-1:0] node784;
	wire [16-1:0] node788;
	wire [16-1:0] node791;
	wire [16-1:0] node792;
	wire [16-1:0] node793;
	wire [16-1:0] node796;
	wire [16-1:0] node798;
	wire [16-1:0] node801;
	wire [16-1:0] node804;
	wire [16-1:0] node805;
	wire [16-1:0] node806;
	wire [16-1:0] node809;
	wire [16-1:0] node811;
	wire [16-1:0] node812;
	wire [16-1:0] node814;
	wire [16-1:0] node818;
	wire [16-1:0] node819;
	wire [16-1:0] node820;
	wire [16-1:0] node821;
	wire [16-1:0] node824;
	wire [16-1:0] node825;
	wire [16-1:0] node829;
	wire [16-1:0] node832;
	wire [16-1:0] node833;
	wire [16-1:0] node834;
	wire [16-1:0] node838;
	wire [16-1:0] node840;
	wire [16-1:0] node843;
	wire [16-1:0] node844;
	wire [16-1:0] node845;
	wire [16-1:0] node846;
	wire [16-1:0] node848;
	wire [16-1:0] node851;
	wire [16-1:0] node853;
	wire [16-1:0] node856;
	wire [16-1:0] node857;
	wire [16-1:0] node858;
	wire [16-1:0] node859;
	wire [16-1:0] node863;
	wire [16-1:0] node865;
	wire [16-1:0] node866;
	wire [16-1:0] node868;
	wire [16-1:0] node872;
	wire [16-1:0] node873;
	wire [16-1:0] node875;
	wire [16-1:0] node878;
	wire [16-1:0] node879;
	wire [16-1:0] node880;
	wire [16-1:0] node882;
	wire [16-1:0] node885;
	wire [16-1:0] node889;
	wire [16-1:0] node890;
	wire [16-1:0] node891;
	wire [16-1:0] node892;
	wire [16-1:0] node896;
	wire [16-1:0] node898;
	wire [16-1:0] node899;
	wire [16-1:0] node903;
	wire [16-1:0] node904;
	wire [16-1:0] node905;
	wire [16-1:0] node908;
	wire [16-1:0] node911;
	wire [16-1:0] node913;
	wire [16-1:0] node915;
	wire [16-1:0] node917;
	wire [16-1:0] node920;
	wire [16-1:0] node921;
	wire [16-1:0] node922;
	wire [16-1:0] node923;
	wire [16-1:0] node924;
	wire [16-1:0] node925;
	wire [16-1:0] node926;
	wire [16-1:0] node928;
	wire [16-1:0] node932;
	wire [16-1:0] node935;
	wire [16-1:0] node936;
	wire [16-1:0] node937;
	wire [16-1:0] node939;
	wire [16-1:0] node943;
	wire [16-1:0] node945;
	wire [16-1:0] node948;
	wire [16-1:0] node949;
	wire [16-1:0] node950;
	wire [16-1:0] node951;
	wire [16-1:0] node952;
	wire [16-1:0] node956;
	wire [16-1:0] node959;
	wire [16-1:0] node961;
	wire [16-1:0] node964;
	wire [16-1:0] node965;
	wire [16-1:0] node966;
	wire [16-1:0] node969;
	wire [16-1:0] node972;
	wire [16-1:0] node973;
	wire [16-1:0] node977;
	wire [16-1:0] node978;
	wire [16-1:0] node979;
	wire [16-1:0] node980;
	wire [16-1:0] node981;
	wire [16-1:0] node983;
	wire [16-1:0] node987;
	wire [16-1:0] node988;
	wire [16-1:0] node991;
	wire [16-1:0] node993;
	wire [16-1:0] node995;
	wire [16-1:0] node998;
	wire [16-1:0] node999;
	wire [16-1:0] node1000;
	wire [16-1:0] node1001;
	wire [16-1:0] node1004;
	wire [16-1:0] node1008;
	wire [16-1:0] node1009;
	wire [16-1:0] node1012;
	wire [16-1:0] node1015;
	wire [16-1:0] node1016;
	wire [16-1:0] node1017;
	wire [16-1:0] node1019;
	wire [16-1:0] node1021;
	wire [16-1:0] node1024;
	wire [16-1:0] node1025;
	wire [16-1:0] node1026;
	wire [16-1:0] node1030;
	wire [16-1:0] node1031;
	wire [16-1:0] node1033;
	wire [16-1:0] node1037;
	wire [16-1:0] node1038;
	wire [16-1:0] node1039;
	wire [16-1:0] node1043;
	wire [16-1:0] node1045;
	wire [16-1:0] node1047;
	wire [16-1:0] node1050;
	wire [16-1:0] node1051;
	wire [16-1:0] node1052;
	wire [16-1:0] node1053;
	wire [16-1:0] node1055;
	wire [16-1:0] node1056;
	wire [16-1:0] node1057;
	wire [16-1:0] node1061;
	wire [16-1:0] node1064;
	wire [16-1:0] node1065;
	wire [16-1:0] node1067;
	wire [16-1:0] node1068;
	wire [16-1:0] node1069;
	wire [16-1:0] node1075;
	wire [16-1:0] node1076;
	wire [16-1:0] node1077;
	wire [16-1:0] node1078;
	wire [16-1:0] node1080;
	wire [16-1:0] node1083;
	wire [16-1:0] node1085;
	wire [16-1:0] node1088;
	wire [16-1:0] node1090;
	wire [16-1:0] node1093;
	wire [16-1:0] node1094;
	wire [16-1:0] node1095;
	wire [16-1:0] node1098;
	wire [16-1:0] node1100;
	wire [16-1:0] node1103;
	wire [16-1:0] node1104;
	wire [16-1:0] node1106;
	wire [16-1:0] node1108;
	wire [16-1:0] node1111;
	wire [16-1:0] node1114;
	wire [16-1:0] node1115;
	wire [16-1:0] node1116;
	wire [16-1:0] node1117;
	wire [16-1:0] node1119;
	wire [16-1:0] node1122;
	wire [16-1:0] node1123;
	wire [16-1:0] node1125;
	wire [16-1:0] node1127;
	wire [16-1:0] node1131;
	wire [16-1:0] node1132;
	wire [16-1:0] node1133;
	wire [16-1:0] node1134;
	wire [16-1:0] node1139;
	wire [16-1:0] node1140;
	wire [16-1:0] node1141;
	wire [16-1:0] node1146;
	wire [16-1:0] node1147;
	wire [16-1:0] node1148;
	wire [16-1:0] node1150;
	wire [16-1:0] node1152;
	wire [16-1:0] node1155;
	wire [16-1:0] node1156;
	wire [16-1:0] node1157;
	wire [16-1:0] node1159;
	wire [16-1:0] node1164;
	wire [16-1:0] node1165;
	wire [16-1:0] node1166;
	wire [16-1:0] node1169;
	wire [16-1:0] node1170;
	wire [16-1:0] node1174;
	wire [16-1:0] node1175;
	wire [16-1:0] node1176;
	wire [16-1:0] node1179;
	wire [16-1:0] node1182;
	wire [16-1:0] node1184;
	wire [16-1:0] node1187;
	wire [16-1:0] node1188;
	wire [16-1:0] node1189;
	wire [16-1:0] node1190;
	wire [16-1:0] node1191;
	wire [16-1:0] node1192;
	wire [16-1:0] node1193;
	wire [16-1:0] node1194;
	wire [16-1:0] node1196;
	wire [16-1:0] node1198;
	wire [16-1:0] node1200;
	wire [16-1:0] node1203;
	wire [16-1:0] node1204;
	wire [16-1:0] node1207;
	wire [16-1:0] node1209;
	wire [16-1:0] node1212;
	wire [16-1:0] node1213;
	wire [16-1:0] node1216;
	wire [16-1:0] node1217;
	wire [16-1:0] node1218;
	wire [16-1:0] node1223;
	wire [16-1:0] node1224;
	wire [16-1:0] node1225;
	wire [16-1:0] node1226;
	wire [16-1:0] node1227;
	wire [16-1:0] node1232;
	wire [16-1:0] node1233;
	wire [16-1:0] node1234;
	wire [16-1:0] node1236;
	wire [16-1:0] node1239;
	wire [16-1:0] node1240;
	wire [16-1:0] node1245;
	wire [16-1:0] node1246;
	wire [16-1:0] node1248;
	wire [16-1:0] node1249;
	wire [16-1:0] node1252;
	wire [16-1:0] node1254;
	wire [16-1:0] node1257;
	wire [16-1:0] node1258;
	wire [16-1:0] node1261;
	wire [16-1:0] node1264;
	wire [16-1:0] node1265;
	wire [16-1:0] node1266;
	wire [16-1:0] node1267;
	wire [16-1:0] node1268;
	wire [16-1:0] node1269;
	wire [16-1:0] node1275;
	wire [16-1:0] node1276;
	wire [16-1:0] node1277;
	wire [16-1:0] node1278;
	wire [16-1:0] node1282;
	wire [16-1:0] node1283;
	wire [16-1:0] node1287;
	wire [16-1:0] node1288;
	wire [16-1:0] node1290;
	wire [16-1:0] node1294;
	wire [16-1:0] node1295;
	wire [16-1:0] node1296;
	wire [16-1:0] node1298;
	wire [16-1:0] node1300;
	wire [16-1:0] node1303;
	wire [16-1:0] node1304;
	wire [16-1:0] node1307;
	wire [16-1:0] node1309;
	wire [16-1:0] node1312;
	wire [16-1:0] node1313;
	wire [16-1:0] node1315;
	wire [16-1:0] node1316;
	wire [16-1:0] node1318;
	wire [16-1:0] node1322;
	wire [16-1:0] node1325;
	wire [16-1:0] node1326;
	wire [16-1:0] node1327;
	wire [16-1:0] node1328;
	wire [16-1:0] node1329;
	wire [16-1:0] node1330;
	wire [16-1:0] node1333;
	wire [16-1:0] node1334;
	wire [16-1:0] node1336;
	wire [16-1:0] node1340;
	wire [16-1:0] node1341;
	wire [16-1:0] node1343;
	wire [16-1:0] node1346;
	wire [16-1:0] node1349;
	wire [16-1:0] node1350;
	wire [16-1:0] node1351;
	wire [16-1:0] node1353;
	wire [16-1:0] node1356;
	wire [16-1:0] node1357;
	wire [16-1:0] node1361;
	wire [16-1:0] node1362;
	wire [16-1:0] node1366;
	wire [16-1:0] node1367;
	wire [16-1:0] node1368;
	wire [16-1:0] node1369;
	wire [16-1:0] node1372;
	wire [16-1:0] node1374;
	wire [16-1:0] node1377;
	wire [16-1:0] node1380;
	wire [16-1:0] node1381;
	wire [16-1:0] node1382;
	wire [16-1:0] node1385;
	wire [16-1:0] node1387;
	wire [16-1:0] node1390;
	wire [16-1:0] node1391;
	wire [16-1:0] node1394;
	wire [16-1:0] node1397;
	wire [16-1:0] node1398;
	wire [16-1:0] node1399;
	wire [16-1:0] node1400;
	wire [16-1:0] node1401;
	wire [16-1:0] node1404;
	wire [16-1:0] node1408;
	wire [16-1:0] node1409;
	wire [16-1:0] node1410;
	wire [16-1:0] node1412;
	wire [16-1:0] node1415;
	wire [16-1:0] node1416;
	wire [16-1:0] node1420;
	wire [16-1:0] node1422;
	wire [16-1:0] node1424;
	wire [16-1:0] node1427;
	wire [16-1:0] node1428;
	wire [16-1:0] node1429;
	wire [16-1:0] node1430;
	wire [16-1:0] node1431;
	wire [16-1:0] node1432;
	wire [16-1:0] node1437;
	wire [16-1:0] node1439;
	wire [16-1:0] node1442;
	wire [16-1:0] node1444;
	wire [16-1:0] node1446;
	wire [16-1:0] node1449;
	wire [16-1:0] node1450;
	wire [16-1:0] node1451;
	wire [16-1:0] node1453;
	wire [16-1:0] node1456;
	wire [16-1:0] node1458;
	wire [16-1:0] node1461;
	wire [16-1:0] node1462;
	wire [16-1:0] node1463;
	wire [16-1:0] node1466;
	wire [16-1:0] node1467;
	wire [16-1:0] node1471;
	wire [16-1:0] node1472;
	wire [16-1:0] node1476;
	wire [16-1:0] node1477;
	wire [16-1:0] node1478;
	wire [16-1:0] node1479;
	wire [16-1:0] node1480;
	wire [16-1:0] node1481;
	wire [16-1:0] node1482;
	wire [16-1:0] node1485;
	wire [16-1:0] node1486;
	wire [16-1:0] node1488;
	wire [16-1:0] node1492;
	wire [16-1:0] node1493;
	wire [16-1:0] node1497;
	wire [16-1:0] node1498;
	wire [16-1:0] node1499;
	wire [16-1:0] node1502;
	wire [16-1:0] node1503;
	wire [16-1:0] node1504;
	wire [16-1:0] node1508;
	wire [16-1:0] node1511;
	wire [16-1:0] node1512;
	wire [16-1:0] node1513;
	wire [16-1:0] node1515;
	wire [16-1:0] node1520;
	wire [16-1:0] node1521;
	wire [16-1:0] node1522;
	wire [16-1:0] node1524;
	wire [16-1:0] node1525;
	wire [16-1:0] node1528;
	wire [16-1:0] node1529;
	wire [16-1:0] node1533;
	wire [16-1:0] node1534;
	wire [16-1:0] node1536;
	wire [16-1:0] node1538;
	wire [16-1:0] node1540;
	wire [16-1:0] node1544;
	wire [16-1:0] node1545;
	wire [16-1:0] node1546;
	wire [16-1:0] node1549;
	wire [16-1:0] node1552;
	wire [16-1:0] node1553;
	wire [16-1:0] node1554;
	wire [16-1:0] node1559;
	wire [16-1:0] node1560;
	wire [16-1:0] node1561;
	wire [16-1:0] node1562;
	wire [16-1:0] node1563;
	wire [16-1:0] node1566;
	wire [16-1:0] node1567;
	wire [16-1:0] node1568;
	wire [16-1:0] node1573;
	wire [16-1:0] node1574;
	wire [16-1:0] node1577;
	wire [16-1:0] node1580;
	wire [16-1:0] node1581;
	wire [16-1:0] node1584;
	wire [16-1:0] node1585;
	wire [16-1:0] node1587;
	wire [16-1:0] node1589;
	wire [16-1:0] node1592;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1597;
	wire [16-1:0] node1599;
	wire [16-1:0] node1602;
	wire [16-1:0] node1603;
	wire [16-1:0] node1604;
	wire [16-1:0] node1608;
	wire [16-1:0] node1609;
	wire [16-1:0] node1612;
	wire [16-1:0] node1615;
	wire [16-1:0] node1616;
	wire [16-1:0] node1618;
	wire [16-1:0] node1621;
	wire [16-1:0] node1622;
	wire [16-1:0] node1623;
	wire [16-1:0] node1627;
	wire [16-1:0] node1629;
	wire [16-1:0] node1630;
	wire [16-1:0] node1634;
	wire [16-1:0] node1635;
	wire [16-1:0] node1636;
	wire [16-1:0] node1637;
	wire [16-1:0] node1639;
	wire [16-1:0] node1642;
	wire [16-1:0] node1643;
	wire [16-1:0] node1645;
	wire [16-1:0] node1647;
	wire [16-1:0] node1651;
	wire [16-1:0] node1652;
	wire [16-1:0] node1653;
	wire [16-1:0] node1655;
	wire [16-1:0] node1656;
	wire [16-1:0] node1660;
	wire [16-1:0] node1661;
	wire [16-1:0] node1663;
	wire [16-1:0] node1667;
	wire [16-1:0] node1668;
	wire [16-1:0] node1669;
	wire [16-1:0] node1673;
	wire [16-1:0] node1676;
	wire [16-1:0] node1677;
	wire [16-1:0] node1678;
	wire [16-1:0] node1679;
	wire [16-1:0] node1680;
	wire [16-1:0] node1681;
	wire [16-1:0] node1686;
	wire [16-1:0] node1688;
	wire [16-1:0] node1691;
	wire [16-1:0] node1692;
	wire [16-1:0] node1693;
	wire [16-1:0] node1694;
	wire [16-1:0] node1695;
	wire [16-1:0] node1700;
	wire [16-1:0] node1702;
	wire [16-1:0] node1705;
	wire [16-1:0] node1707;
	wire [16-1:0] node1708;
	wire [16-1:0] node1712;
	wire [16-1:0] node1713;
	wire [16-1:0] node1714;
	wire [16-1:0] node1715;
	wire [16-1:0] node1719;
	wire [16-1:0] node1722;
	wire [16-1:0] node1723;
	wire [16-1:0] node1724;
	wire [16-1:0] node1728;
	wire [16-1:0] node1729;
	wire [16-1:0] node1733;
	wire [16-1:0] node1734;
	wire [16-1:0] node1735;
	wire [16-1:0] node1736;
	wire [16-1:0] node1737;
	wire [16-1:0] node1738;
	wire [16-1:0] node1739;
	wire [16-1:0] node1740;
	wire [16-1:0] node1743;
	wire [16-1:0] node1744;
	wire [16-1:0] node1746;
	wire [16-1:0] node1750;
	wire [16-1:0] node1751;
	wire [16-1:0] node1752;
	wire [16-1:0] node1756;
	wire [16-1:0] node1759;
	wire [16-1:0] node1760;
	wire [16-1:0] node1763;
	wire [16-1:0] node1764;
	wire [16-1:0] node1765;
	wire [16-1:0] node1769;
	wire [16-1:0] node1772;
	wire [16-1:0] node1773;
	wire [16-1:0] node1774;
	wire [16-1:0] node1775;
	wire [16-1:0] node1778;
	wire [16-1:0] node1780;
	wire [16-1:0] node1783;
	wire [16-1:0] node1784;
	wire [16-1:0] node1788;
	wire [16-1:0] node1789;
	wire [16-1:0] node1790;
	wire [16-1:0] node1791;
	wire [16-1:0] node1796;
	wire [16-1:0] node1797;
	wire [16-1:0] node1799;
	wire [16-1:0] node1800;
	wire [16-1:0] node1804;
	wire [16-1:0] node1807;
	wire [16-1:0] node1808;
	wire [16-1:0] node1809;
	wire [16-1:0] node1810;
	wire [16-1:0] node1811;
	wire [16-1:0] node1813;
	wire [16-1:0] node1817;
	wire [16-1:0] node1818;
	wire [16-1:0] node1820;
	wire [16-1:0] node1822;
	wire [16-1:0] node1823;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1831;
	wire [16-1:0] node1833;
	wire [16-1:0] node1836;
	wire [16-1:0] node1837;
	wire [16-1:0] node1841;
	wire [16-1:0] node1842;
	wire [16-1:0] node1844;
	wire [16-1:0] node1845;
	wire [16-1:0] node1847;
	wire [16-1:0] node1848;
	wire [16-1:0] node1853;
	wire [16-1:0] node1854;
	wire [16-1:0] node1856;
	wire [16-1:0] node1857;
	wire [16-1:0] node1861;
	wire [16-1:0] node1864;
	wire [16-1:0] node1865;
	wire [16-1:0] node1866;
	wire [16-1:0] node1867;
	wire [16-1:0] node1868;
	wire [16-1:0] node1869;
	wire [16-1:0] node1870;
	wire [16-1:0] node1874;
	wire [16-1:0] node1875;
	wire [16-1:0] node1877;
	wire [16-1:0] node1880;
	wire [16-1:0] node1883;
	wire [16-1:0] node1886;
	wire [16-1:0] node1887;
	wire [16-1:0] node1889;
	wire [16-1:0] node1890;
	wire [16-1:0] node1894;
	wire [16-1:0] node1897;
	wire [16-1:0] node1898;
	wire [16-1:0] node1899;
	wire [16-1:0] node1900;
	wire [16-1:0] node1903;
	wire [16-1:0] node1905;
	wire [16-1:0] node1908;
	wire [16-1:0] node1909;
	wire [16-1:0] node1911;
	wire [16-1:0] node1912;
	wire [16-1:0] node1916;
	wire [16-1:0] node1918;
	wire [16-1:0] node1921;
	wire [16-1:0] node1922;
	wire [16-1:0] node1925;
	wire [16-1:0] node1927;
	wire [16-1:0] node1929;
	wire [16-1:0] node1930;
	wire [16-1:0] node1932;
	wire [16-1:0] node1936;
	wire [16-1:0] node1937;
	wire [16-1:0] node1938;
	wire [16-1:0] node1939;
	wire [16-1:0] node1940;
	wire [16-1:0] node1942;
	wire [16-1:0] node1946;
	wire [16-1:0] node1947;
	wire [16-1:0] node1950;
	wire [16-1:0] node1952;
	wire [16-1:0] node1954;
	wire [16-1:0] node1957;
	wire [16-1:0] node1958;
	wire [16-1:0] node1960;
	wire [16-1:0] node1963;
	wire [16-1:0] node1965;
	wire [16-1:0] node1966;
	wire [16-1:0] node1969;
	wire [16-1:0] node1972;
	wire [16-1:0] node1973;
	wire [16-1:0] node1974;
	wire [16-1:0] node1975;
	wire [16-1:0] node1978;
	wire [16-1:0] node1981;
	wire [16-1:0] node1982;
	wire [16-1:0] node1986;
	wire [16-1:0] node1987;
	wire [16-1:0] node1988;
	wire [16-1:0] node1989;
	wire [16-1:0] node1994;
	wire [16-1:0] node1995;
	wire [16-1:0] node1998;
	wire [16-1:0] node2000;
	wire [16-1:0] node2003;
	wire [16-1:0] node2004;
	wire [16-1:0] node2005;
	wire [16-1:0] node2006;
	wire [16-1:0] node2007;
	wire [16-1:0] node2008;
	wire [16-1:0] node2009;
	wire [16-1:0] node2010;
	wire [16-1:0] node2014;
	wire [16-1:0] node2016;
	wire [16-1:0] node2019;
	wire [16-1:0] node2022;
	wire [16-1:0] node2023;
	wire [16-1:0] node2024;
	wire [16-1:0] node2026;
	wire [16-1:0] node2029;
	wire [16-1:0] node2031;
	wire [16-1:0] node2034;
	wire [16-1:0] node2036;
	wire [16-1:0] node2037;
	wire [16-1:0] node2041;
	wire [16-1:0] node2042;
	wire [16-1:0] node2044;
	wire [16-1:0] node2045;
	wire [16-1:0] node2048;
	wire [16-1:0] node2049;
	wire [16-1:0] node2053;
	wire [16-1:0] node2054;
	wire [16-1:0] node2055;
	wire [16-1:0] node2057;
	wire [16-1:0] node2060;
	wire [16-1:0] node2063;
	wire [16-1:0] node2065;
	wire [16-1:0] node2068;
	wire [16-1:0] node2069;
	wire [16-1:0] node2070;
	wire [16-1:0] node2071;
	wire [16-1:0] node2073;
	wire [16-1:0] node2075;
	wire [16-1:0] node2078;
	wire [16-1:0] node2080;
	wire [16-1:0] node2081;
	wire [16-1:0] node2084;
	wire [16-1:0] node2087;
	wire [16-1:0] node2088;
	wire [16-1:0] node2091;
	wire [16-1:0] node2093;
	wire [16-1:0] node2094;
	wire [16-1:0] node2096;
	wire [16-1:0] node2097;
	wire [16-1:0] node2101;
	wire [16-1:0] node2104;
	wire [16-1:0] node2105;
	wire [16-1:0] node2106;
	wire [16-1:0] node2108;
	wire [16-1:0] node2109;
	wire [16-1:0] node2113;
	wire [16-1:0] node2114;
	wire [16-1:0] node2115;
	wire [16-1:0] node2116;
	wire [16-1:0] node2119;
	wire [16-1:0] node2121;
	wire [16-1:0] node2124;
	wire [16-1:0] node2125;
	wire [16-1:0] node2130;
	wire [16-1:0] node2131;
	wire [16-1:0] node2132;
	wire [16-1:0] node2134;
	wire [16-1:0] node2137;
	wire [16-1:0] node2140;
	wire [16-1:0] node2142;
	wire [16-1:0] node2143;
	wire [16-1:0] node2144;
	wire [16-1:0] node2149;
	wire [16-1:0] node2150;
	wire [16-1:0] node2151;
	wire [16-1:0] node2152;
	wire [16-1:0] node2153;
	wire [16-1:0] node2155;
	wire [16-1:0] node2157;
	wire [16-1:0] node2160;
	wire [16-1:0] node2162;
	wire [16-1:0] node2163;
	wire [16-1:0] node2167;
	wire [16-1:0] node2168;
	wire [16-1:0] node2170;
	wire [16-1:0] node2172;
	wire [16-1:0] node2175;
	wire [16-1:0] node2177;
	wire [16-1:0] node2178;
	wire [16-1:0] node2179;
	wire [16-1:0] node2182;
	wire [16-1:0] node2183;
	wire [16-1:0] node2184;
	wire [16-1:0] node2189;
	wire [16-1:0] node2191;
	wire [16-1:0] node2194;
	wire [16-1:0] node2195;
	wire [16-1:0] node2196;
	wire [16-1:0] node2197;
	wire [16-1:0] node2200;
	wire [16-1:0] node2201;
	wire [16-1:0] node2205;
	wire [16-1:0] node2206;
	wire [16-1:0] node2209;
	wire [16-1:0] node2212;
	wire [16-1:0] node2213;
	wire [16-1:0] node2215;
	wire [16-1:0] node2216;
	wire [16-1:0] node2217;
	wire [16-1:0] node2222;
	wire [16-1:0] node2225;
	wire [16-1:0] node2226;
	wire [16-1:0] node2227;
	wire [16-1:0] node2228;
	wire [16-1:0] node2231;
	wire [16-1:0] node2232;
	wire [16-1:0] node2234;
	wire [16-1:0] node2238;
	wire [16-1:0] node2239;
	wire [16-1:0] node2240;
	wire [16-1:0] node2243;
	wire [16-1:0] node2246;
	wire [16-1:0] node2249;
	wire [16-1:0] node2250;
	wire [16-1:0] node2251;
	wire [16-1:0] node2254;
	wire [16-1:0] node2255;
	wire [16-1:0] node2257;
	wire [16-1:0] node2258;
	wire [16-1:0] node2263;
	wire [16-1:0] node2264;
	wire [16-1:0] node2266;
	wire [16-1:0] node2269;
	wire [16-1:0] node2270;
	wire [16-1:0] node2273;
	wire [16-1:0] node2274;
	wire [16-1:0] node2277;
	wire [16-1:0] node2279;
	wire [16-1:0] node2282;
	wire [16-1:0] node2283;
	wire [16-1:0] node2284;
	wire [16-1:0] node2285;
	wire [16-1:0] node2286;
	wire [16-1:0] node2287;
	wire [16-1:0] node2288;
	wire [16-1:0] node2289;
	wire [16-1:0] node2290;
	wire [16-1:0] node2291;
	wire [16-1:0] node2292;
	wire [16-1:0] node2297;
	wire [16-1:0] node2298;
	wire [16-1:0] node2301;
	wire [16-1:0] node2303;
	wire [16-1:0] node2306;
	wire [16-1:0] node2307;
	wire [16-1:0] node2308;
	wire [16-1:0] node2309;
	wire [16-1:0] node2312;
	wire [16-1:0] node2315;
	wire [16-1:0] node2316;
	wire [16-1:0] node2318;
	wire [16-1:0] node2319;
	wire [16-1:0] node2324;
	wire [16-1:0] node2325;
	wire [16-1:0] node2326;
	wire [16-1:0] node2329;
	wire [16-1:0] node2332;
	wire [16-1:0] node2335;
	wire [16-1:0] node2336;
	wire [16-1:0] node2337;
	wire [16-1:0] node2338;
	wire [16-1:0] node2340;
	wire [16-1:0] node2343;
	wire [16-1:0] node2346;
	wire [16-1:0] node2347;
	wire [16-1:0] node2348;
	wire [16-1:0] node2352;
	wire [16-1:0] node2353;
	wire [16-1:0] node2357;
	wire [16-1:0] node2358;
	wire [16-1:0] node2360;
	wire [16-1:0] node2362;
	wire [16-1:0] node2365;
	wire [16-1:0] node2366;
	wire [16-1:0] node2369;
	wire [16-1:0] node2371;
	wire [16-1:0] node2374;
	wire [16-1:0] node2375;
	wire [16-1:0] node2376;
	wire [16-1:0] node2377;
	wire [16-1:0] node2378;
	wire [16-1:0] node2381;
	wire [16-1:0] node2383;
	wire [16-1:0] node2386;
	wire [16-1:0] node2387;
	wire [16-1:0] node2388;
	wire [16-1:0] node2391;
	wire [16-1:0] node2394;
	wire [16-1:0] node2397;
	wire [16-1:0] node2398;
	wire [16-1:0] node2399;
	wire [16-1:0] node2400;
	wire [16-1:0] node2404;
	wire [16-1:0] node2405;
	wire [16-1:0] node2408;
	wire [16-1:0] node2411;
	wire [16-1:0] node2412;
	wire [16-1:0] node2414;
	wire [16-1:0] node2417;
	wire [16-1:0] node2419;
	wire [16-1:0] node2422;
	wire [16-1:0] node2423;
	wire [16-1:0] node2424;
	wire [16-1:0] node2427;
	wire [16-1:0] node2430;
	wire [16-1:0] node2431;
	wire [16-1:0] node2434;
	wire [16-1:0] node2435;
	wire [16-1:0] node2437;
	wire [16-1:0] node2440;
	wire [16-1:0] node2443;
	wire [16-1:0] node2444;
	wire [16-1:0] node2445;
	wire [16-1:0] node2446;
	wire [16-1:0] node2447;
	wire [16-1:0] node2448;
	wire [16-1:0] node2451;
	wire [16-1:0] node2452;
	wire [16-1:0] node2456;
	wire [16-1:0] node2457;
	wire [16-1:0] node2459;
	wire [16-1:0] node2462;
	wire [16-1:0] node2464;
	wire [16-1:0] node2467;
	wire [16-1:0] node2468;
	wire [16-1:0] node2469;
	wire [16-1:0] node2470;
	wire [16-1:0] node2471;
	wire [16-1:0] node2476;
	wire [16-1:0] node2478;
	wire [16-1:0] node2481;
	wire [16-1:0] node2484;
	wire [16-1:0] node2485;
	wire [16-1:0] node2486;
	wire [16-1:0] node2489;
	wire [16-1:0] node2490;
	wire [16-1:0] node2494;
	wire [16-1:0] node2495;
	wire [16-1:0] node2496;
	wire [16-1:0] node2498;
	wire [16-1:0] node2501;
	wire [16-1:0] node2504;
	wire [16-1:0] node2507;
	wire [16-1:0] node2508;
	wire [16-1:0] node2509;
	wire [16-1:0] node2510;
	wire [16-1:0] node2511;
	wire [16-1:0] node2514;
	wire [16-1:0] node2516;
	wire [16-1:0] node2519;
	wire [16-1:0] node2520;
	wire [16-1:0] node2521;
	wire [16-1:0] node2525;
	wire [16-1:0] node2526;
	wire [16-1:0] node2529;
	wire [16-1:0] node2532;
	wire [16-1:0] node2533;
	wire [16-1:0] node2535;
	wire [16-1:0] node2536;
	wire [16-1:0] node2538;
	wire [16-1:0] node2539;
	wire [16-1:0] node2540;
	wire [16-1:0] node2542;
	wire [16-1:0] node2547;
	wire [16-1:0] node2550;
	wire [16-1:0] node2551;
	wire [16-1:0] node2555;
	wire [16-1:0] node2556;
	wire [16-1:0] node2557;
	wire [16-1:0] node2558;
	wire [16-1:0] node2562;
	wire [16-1:0] node2564;
	wire [16-1:0] node2565;
	wire [16-1:0] node2569;
	wire [16-1:0] node2570;
	wire [16-1:0] node2571;
	wire [16-1:0] node2575;
	wire [16-1:0] node2576;
	wire [16-1:0] node2577;
	wire [16-1:0] node2582;
	wire [16-1:0] node2583;
	wire [16-1:0] node2584;
	wire [16-1:0] node2585;
	wire [16-1:0] node2586;
	wire [16-1:0] node2587;
	wire [16-1:0] node2588;
	wire [16-1:0] node2589;
	wire [16-1:0] node2593;
	wire [16-1:0] node2596;
	wire [16-1:0] node2597;
	wire [16-1:0] node2601;
	wire [16-1:0] node2602;
	wire [16-1:0] node2603;
	wire [16-1:0] node2604;
	wire [16-1:0] node2607;
	wire [16-1:0] node2611;
	wire [16-1:0] node2613;
	wire [16-1:0] node2616;
	wire [16-1:0] node2617;
	wire [16-1:0] node2618;
	wire [16-1:0] node2620;
	wire [16-1:0] node2622;
	wire [16-1:0] node2625;
	wire [16-1:0] node2626;
	wire [16-1:0] node2629;
	wire [16-1:0] node2630;
	wire [16-1:0] node2631;
	wire [16-1:0] node2635;
	wire [16-1:0] node2638;
	wire [16-1:0] node2639;
	wire [16-1:0] node2640;
	wire [16-1:0] node2644;
	wire [16-1:0] node2646;
	wire [16-1:0] node2649;
	wire [16-1:0] node2650;
	wire [16-1:0] node2651;
	wire [16-1:0] node2652;
	wire [16-1:0] node2653;
	wire [16-1:0] node2655;
	wire [16-1:0] node2659;
	wire [16-1:0] node2661;
	wire [16-1:0] node2662;
	wire [16-1:0] node2664;
	wire [16-1:0] node2668;
	wire [16-1:0] node2669;
	wire [16-1:0] node2670;
	wire [16-1:0] node2671;
	wire [16-1:0] node2672;
	wire [16-1:0] node2677;
	wire [16-1:0] node2678;
	wire [16-1:0] node2681;
	wire [16-1:0] node2682;
	wire [16-1:0] node2686;
	wire [16-1:0] node2687;
	wire [16-1:0] node2691;
	wire [16-1:0] node2692;
	wire [16-1:0] node2693;
	wire [16-1:0] node2694;
	wire [16-1:0] node2697;
	wire [16-1:0] node2698;
	wire [16-1:0] node2702;
	wire [16-1:0] node2703;
	wire [16-1:0] node2704;
	wire [16-1:0] node2705;
	wire [16-1:0] node2706;
	wire [16-1:0] node2711;
	wire [16-1:0] node2713;
	wire [16-1:0] node2716;
	wire [16-1:0] node2717;
	wire [16-1:0] node2718;
	wire [16-1:0] node2723;
	wire [16-1:0] node2724;
	wire [16-1:0] node2725;
	wire [16-1:0] node2727;
	wire [16-1:0] node2731;
	wire [16-1:0] node2732;
	wire [16-1:0] node2735;
	wire [16-1:0] node2736;
	wire [16-1:0] node2740;
	wire [16-1:0] node2741;
	wire [16-1:0] node2742;
	wire [16-1:0] node2743;
	wire [16-1:0] node2744;
	wire [16-1:0] node2745;
	wire [16-1:0] node2746;
	wire [16-1:0] node2750;
	wire [16-1:0] node2753;
	wire [16-1:0] node2756;
	wire [16-1:0] node2757;
	wire [16-1:0] node2758;
	wire [16-1:0] node2759;
	wire [16-1:0] node2762;
	wire [16-1:0] node2766;
	wire [16-1:0] node2769;
	wire [16-1:0] node2770;
	wire [16-1:0] node2771;
	wire [16-1:0] node2772;
	wire [16-1:0] node2773;
	wire [16-1:0] node2777;
	wire [16-1:0] node2778;
	wire [16-1:0] node2782;
	wire [16-1:0] node2783;
	wire [16-1:0] node2785;
	wire [16-1:0] node2787;
	wire [16-1:0] node2791;
	wire [16-1:0] node2793;
	wire [16-1:0] node2795;
	wire [16-1:0] node2796;
	wire [16-1:0] node2800;
	wire [16-1:0] node2801;
	wire [16-1:0] node2802;
	wire [16-1:0] node2803;
	wire [16-1:0] node2804;
	wire [16-1:0] node2807;
	wire [16-1:0] node2810;
	wire [16-1:0] node2811;
	wire [16-1:0] node2812;
	wire [16-1:0] node2814;
	wire [16-1:0] node2819;
	wire [16-1:0] node2820;
	wire [16-1:0] node2821;
	wire [16-1:0] node2825;
	wire [16-1:0] node2827;
	wire [16-1:0] node2830;
	wire [16-1:0] node2831;
	wire [16-1:0] node2832;
	wire [16-1:0] node2833;
	wire [16-1:0] node2836;
	wire [16-1:0] node2837;
	wire [16-1:0] node2840;
	wire [16-1:0] node2843;
	wire [16-1:0] node2844;
	wire [16-1:0] node2845;
	wire [16-1:0] node2849;
	wire [16-1:0] node2850;
	wire [16-1:0] node2851;
	wire [16-1:0] node2854;
	wire [16-1:0] node2858;
	wire [16-1:0] node2860;
	wire [16-1:0] node2862;
	wire [16-1:0] node2863;
	wire [16-1:0] node2867;
	wire [16-1:0] node2868;
	wire [16-1:0] node2869;
	wire [16-1:0] node2870;
	wire [16-1:0] node2871;
	wire [16-1:0] node2872;
	wire [16-1:0] node2873;
	wire [16-1:0] node2874;
	wire [16-1:0] node2875;
	wire [16-1:0] node2879;
	wire [16-1:0] node2881;
	wire [16-1:0] node2884;
	wire [16-1:0] node2885;
	wire [16-1:0] node2886;
	wire [16-1:0] node2890;
	wire [16-1:0] node2892;
	wire [16-1:0] node2895;
	wire [16-1:0] node2896;
	wire [16-1:0] node2898;
	wire [16-1:0] node2900;
	wire [16-1:0] node2903;
	wire [16-1:0] node2904;
	wire [16-1:0] node2905;
	wire [16-1:0] node2910;
	wire [16-1:0] node2911;
	wire [16-1:0] node2912;
	wire [16-1:0] node2913;
	wire [16-1:0] node2915;
	wire [16-1:0] node2917;
	wire [16-1:0] node2920;
	wire [16-1:0] node2921;
	wire [16-1:0] node2923;
	wire [16-1:0] node2924;
	wire [16-1:0] node2929;
	wire [16-1:0] node2932;
	wire [16-1:0] node2933;
	wire [16-1:0] node2934;
	wire [16-1:0] node2937;
	wire [16-1:0] node2938;
	wire [16-1:0] node2942;
	wire [16-1:0] node2944;
	wire [16-1:0] node2947;
	wire [16-1:0] node2948;
	wire [16-1:0] node2949;
	wire [16-1:0] node2950;
	wire [16-1:0] node2951;
	wire [16-1:0] node2952;
	wire [16-1:0] node2956;
	wire [16-1:0] node2958;
	wire [16-1:0] node2959;
	wire [16-1:0] node2963;
	wire [16-1:0] node2965;
	wire [16-1:0] node2968;
	wire [16-1:0] node2969;
	wire [16-1:0] node2970;
	wire [16-1:0] node2972;
	wire [16-1:0] node2976;
	wire [16-1:0] node2977;
	wire [16-1:0] node2978;
	wire [16-1:0] node2979;
	wire [16-1:0] node2983;
	wire [16-1:0] node2986;
	wire [16-1:0] node2987;
	wire [16-1:0] node2991;
	wire [16-1:0] node2992;
	wire [16-1:0] node2993;
	wire [16-1:0] node2994;
	wire [16-1:0] node2996;
	wire [16-1:0] node3000;
	wire [16-1:0] node3001;
	wire [16-1:0] node3004;
	wire [16-1:0] node3006;
	wire [16-1:0] node3009;
	wire [16-1:0] node3010;
	wire [16-1:0] node3011;
	wire [16-1:0] node3014;
	wire [16-1:0] node3016;
	wire [16-1:0] node3019;
	wire [16-1:0] node3020;
	wire [16-1:0] node3022;
	wire [16-1:0] node3025;
	wire [16-1:0] node3026;
	wire [16-1:0] node3029;
	wire [16-1:0] node3031;
	wire [16-1:0] node3034;
	wire [16-1:0] node3035;
	wire [16-1:0] node3036;
	wire [16-1:0] node3037;
	wire [16-1:0] node3038;
	wire [16-1:0] node3040;
	wire [16-1:0] node3041;
	wire [16-1:0] node3045;
	wire [16-1:0] node3046;
	wire [16-1:0] node3049;
	wire [16-1:0] node3052;
	wire [16-1:0] node3053;
	wire [16-1:0] node3054;
	wire [16-1:0] node3055;
	wire [16-1:0] node3059;
	wire [16-1:0] node3061;
	wire [16-1:0] node3064;
	wire [16-1:0] node3066;
	wire [16-1:0] node3069;
	wire [16-1:0] node3070;
	wire [16-1:0] node3071;
	wire [16-1:0] node3073;
	wire [16-1:0] node3074;
	wire [16-1:0] node3078;
	wire [16-1:0] node3080;
	wire [16-1:0] node3083;
	wire [16-1:0] node3084;
	wire [16-1:0] node3085;
	wire [16-1:0] node3089;
	wire [16-1:0] node3090;
	wire [16-1:0] node3092;
	wire [16-1:0] node3095;
	wire [16-1:0] node3098;
	wire [16-1:0] node3099;
	wire [16-1:0] node3100;
	wire [16-1:0] node3101;
	wire [16-1:0] node3103;
	wire [16-1:0] node3106;
	wire [16-1:0] node3107;
	wire [16-1:0] node3109;
	wire [16-1:0] node3113;
	wire [16-1:0] node3114;
	wire [16-1:0] node3117;
	wire [16-1:0] node3119;
	wire [16-1:0] node3121;
	wire [16-1:0] node3124;
	wire [16-1:0] node3125;
	wire [16-1:0] node3126;
	wire [16-1:0] node3128;
	wire [16-1:0] node3132;
	wire [16-1:0] node3133;
	wire [16-1:0] node3134;
	wire [16-1:0] node3136;
	wire [16-1:0] node3140;
	wire [16-1:0] node3142;
	wire [16-1:0] node3145;
	wire [16-1:0] node3146;
	wire [16-1:0] node3147;
	wire [16-1:0] node3148;
	wire [16-1:0] node3149;
	wire [16-1:0] node3150;
	wire [16-1:0] node3151;
	wire [16-1:0] node3153;
	wire [16-1:0] node3157;
	wire [16-1:0] node3159;
	wire [16-1:0] node3162;
	wire [16-1:0] node3163;
	wire [16-1:0] node3164;
	wire [16-1:0] node3167;
	wire [16-1:0] node3168;
	wire [16-1:0] node3172;
	wire [16-1:0] node3173;
	wire [16-1:0] node3174;
	wire [16-1:0] node3177;
	wire [16-1:0] node3180;
	wire [16-1:0] node3183;
	wire [16-1:0] node3184;
	wire [16-1:0] node3185;
	wire [16-1:0] node3186;
	wire [16-1:0] node3187;
	wire [16-1:0] node3191;
	wire [16-1:0] node3192;
	wire [16-1:0] node3196;
	wire [16-1:0] node3198;
	wire [16-1:0] node3201;
	wire [16-1:0] node3202;
	wire [16-1:0] node3203;
	wire [16-1:0] node3207;
	wire [16-1:0] node3208;
	wire [16-1:0] node3211;
	wire [16-1:0] node3214;
	wire [16-1:0] node3215;
	wire [16-1:0] node3216;
	wire [16-1:0] node3217;
	wire [16-1:0] node3218;
	wire [16-1:0] node3221;
	wire [16-1:0] node3223;
	wire [16-1:0] node3226;
	wire [16-1:0] node3228;
	wire [16-1:0] node3229;
	wire [16-1:0] node3233;
	wire [16-1:0] node3234;
	wire [16-1:0] node3235;
	wire [16-1:0] node3238;
	wire [16-1:0] node3239;
	wire [16-1:0] node3243;
	wire [16-1:0] node3245;
	wire [16-1:0] node3248;
	wire [16-1:0] node3249;
	wire [16-1:0] node3250;
	wire [16-1:0] node3251;
	wire [16-1:0] node3253;
	wire [16-1:0] node3257;
	wire [16-1:0] node3259;
	wire [16-1:0] node3262;
	wire [16-1:0] node3263;
	wire [16-1:0] node3264;
	wire [16-1:0] node3266;
	wire [16-1:0] node3267;
	wire [16-1:0] node3269;
	wire [16-1:0] node3273;
	wire [16-1:0] node3274;
	wire [16-1:0] node3276;
	wire [16-1:0] node3280;
	wire [16-1:0] node3281;
	wire [16-1:0] node3282;
	wire [16-1:0] node3287;
	wire [16-1:0] node3288;
	wire [16-1:0] node3289;
	wire [16-1:0] node3290;
	wire [16-1:0] node3292;
	wire [16-1:0] node3293;
	wire [16-1:0] node3295;
	wire [16-1:0] node3297;
	wire [16-1:0] node3300;
	wire [16-1:0] node3303;
	wire [16-1:0] node3304;
	wire [16-1:0] node3305;
	wire [16-1:0] node3309;
	wire [16-1:0] node3312;
	wire [16-1:0] node3313;
	wire [16-1:0] node3314;
	wire [16-1:0] node3316;
	wire [16-1:0] node3318;
	wire [16-1:0] node3321;
	wire [16-1:0] node3322;
	wire [16-1:0] node3324;
	wire [16-1:0] node3327;
	wire [16-1:0] node3328;
	wire [16-1:0] node3329;
	wire [16-1:0] node3333;
	wire [16-1:0] node3336;
	wire [16-1:0] node3337;
	wire [16-1:0] node3339;
	wire [16-1:0] node3341;
	wire [16-1:0] node3342;
	wire [16-1:0] node3346;
	wire [16-1:0] node3348;
	wire [16-1:0] node3349;
	wire [16-1:0] node3352;
	wire [16-1:0] node3354;
	wire [16-1:0] node3355;
	wire [16-1:0] node3358;
	wire [16-1:0] node3361;
	wire [16-1:0] node3362;
	wire [16-1:0] node3363;
	wire [16-1:0] node3364;
	wire [16-1:0] node3367;
	wire [16-1:0] node3368;
	wire [16-1:0] node3369;
	wire [16-1:0] node3373;
	wire [16-1:0] node3374;
	wire [16-1:0] node3378;
	wire [16-1:0] node3379;
	wire [16-1:0] node3380;
	wire [16-1:0] node3381;
	wire [16-1:0] node3386;
	wire [16-1:0] node3387;
	wire [16-1:0] node3389;
	wire [16-1:0] node3390;
	wire [16-1:0] node3393;
	wire [16-1:0] node3397;
	wire [16-1:0] node3398;
	wire [16-1:0] node3399;
	wire [16-1:0] node3400;
	wire [16-1:0] node3402;
	wire [16-1:0] node3405;
	wire [16-1:0] node3408;
	wire [16-1:0] node3409;
	wire [16-1:0] node3411;
	wire [16-1:0] node3412;
	wire [16-1:0] node3416;
	wire [16-1:0] node3419;
	wire [16-1:0] node3420;
	wire [16-1:0] node3421;
	wire [16-1:0] node3423;
	wire [16-1:0] node3426;
	wire [16-1:0] node3429;
	wire [16-1:0] node3430;
	wire [16-1:0] node3432;
	wire [16-1:0] node3434;
	wire [16-1:0] node3437;
	wire [16-1:0] node3439;
	wire [16-1:0] node3441;
	wire [16-1:0] node3443;
	wire [16-1:0] node3446;
	wire [16-1:0] node3447;
	wire [16-1:0] node3448;
	wire [16-1:0] node3449;
	wire [16-1:0] node3450;
	wire [16-1:0] node3451;
	wire [16-1:0] node3452;
	wire [16-1:0] node3453;
	wire [16-1:0] node3454;
	wire [16-1:0] node3455;
	wire [16-1:0] node3460;
	wire [16-1:0] node3461;
	wire [16-1:0] node3464;
	wire [16-1:0] node3467;
	wire [16-1:0] node3468;
	wire [16-1:0] node3469;
	wire [16-1:0] node3472;
	wire [16-1:0] node3475;
	wire [16-1:0] node3476;
	wire [16-1:0] node3477;
	wire [16-1:0] node3481;
	wire [16-1:0] node3482;
	wire [16-1:0] node3486;
	wire [16-1:0] node3487;
	wire [16-1:0] node3488;
	wire [16-1:0] node3489;
	wire [16-1:0] node3490;
	wire [16-1:0] node3494;
	wire [16-1:0] node3495;
	wire [16-1:0] node3499;
	wire [16-1:0] node3500;
	wire [16-1:0] node3502;
	wire [16-1:0] node3506;
	wire [16-1:0] node3507;
	wire [16-1:0] node3509;
	wire [16-1:0] node3512;
	wire [16-1:0] node3514;
	wire [16-1:0] node3517;
	wire [16-1:0] node3518;
	wire [16-1:0] node3519;
	wire [16-1:0] node3520;
	wire [16-1:0] node3523;
	wire [16-1:0] node3524;
	wire [16-1:0] node3526;
	wire [16-1:0] node3527;
	wire [16-1:0] node3532;
	wire [16-1:0] node3533;
	wire [16-1:0] node3536;
	wire [16-1:0] node3537;
	wire [16-1:0] node3538;
	wire [16-1:0] node3540;
	wire [16-1:0] node3545;
	wire [16-1:0] node3546;
	wire [16-1:0] node3547;
	wire [16-1:0] node3550;
	wire [16-1:0] node3551;
	wire [16-1:0] node3553;
	wire [16-1:0] node3557;
	wire [16-1:0] node3558;
	wire [16-1:0] node3560;
	wire [16-1:0] node3561;
	wire [16-1:0] node3565;
	wire [16-1:0] node3567;
	wire [16-1:0] node3570;
	wire [16-1:0] node3571;
	wire [16-1:0] node3572;
	wire [16-1:0] node3573;
	wire [16-1:0] node3574;
	wire [16-1:0] node3575;
	wire [16-1:0] node3578;
	wire [16-1:0] node3579;
	wire [16-1:0] node3583;
	wire [16-1:0] node3586;
	wire [16-1:0] node3587;
	wire [16-1:0] node3588;
	wire [16-1:0] node3590;
	wire [16-1:0] node3593;
	wire [16-1:0] node3596;
	wire [16-1:0] node3597;
	wire [16-1:0] node3601;
	wire [16-1:0] node3602;
	wire [16-1:0] node3603;
	wire [16-1:0] node3605;
	wire [16-1:0] node3606;
	wire [16-1:0] node3610;
	wire [16-1:0] node3611;
	wire [16-1:0] node3614;
	wire [16-1:0] node3617;
	wire [16-1:0] node3618;
	wire [16-1:0] node3619;
	wire [16-1:0] node3620;
	wire [16-1:0] node3624;
	wire [16-1:0] node3625;
	wire [16-1:0] node3627;
	wire [16-1:0] node3631;
	wire [16-1:0] node3634;
	wire [16-1:0] node3635;
	wire [16-1:0] node3636;
	wire [16-1:0] node3637;
	wire [16-1:0] node3639;
	wire [16-1:0] node3642;
	wire [16-1:0] node3643;
	wire [16-1:0] node3646;
	wire [16-1:0] node3647;
	wire [16-1:0] node3651;
	wire [16-1:0] node3652;
	wire [16-1:0] node3653;
	wire [16-1:0] node3656;
	wire [16-1:0] node3658;
	wire [16-1:0] node3661;
	wire [16-1:0] node3662;
	wire [16-1:0] node3666;
	wire [16-1:0] node3667;
	wire [16-1:0] node3668;
	wire [16-1:0] node3670;
	wire [16-1:0] node3673;
	wire [16-1:0] node3674;
	wire [16-1:0] node3676;
	wire [16-1:0] node3679;
	wire [16-1:0] node3682;
	wire [16-1:0] node3683;
	wire [16-1:0] node3684;
	wire [16-1:0] node3686;
	wire [16-1:0] node3689;
	wire [16-1:0] node3691;
	wire [16-1:0] node3694;
	wire [16-1:0] node3696;
	wire [16-1:0] node3697;
	wire [16-1:0] node3701;
	wire [16-1:0] node3702;
	wire [16-1:0] node3703;
	wire [16-1:0] node3704;
	wire [16-1:0] node3705;
	wire [16-1:0] node3706;
	wire [16-1:0] node3707;
	wire [16-1:0] node3709;
	wire [16-1:0] node3712;
	wire [16-1:0] node3716;
	wire [16-1:0] node3717;
	wire [16-1:0] node3718;
	wire [16-1:0] node3719;
	wire [16-1:0] node3724;
	wire [16-1:0] node3726;
	wire [16-1:0] node3729;
	wire [16-1:0] node3730;
	wire [16-1:0] node3731;
	wire [16-1:0] node3732;
	wire [16-1:0] node3736;
	wire [16-1:0] node3737;
	wire [16-1:0] node3738;
	wire [16-1:0] node3743;
	wire [16-1:0] node3744;
	wire [16-1:0] node3745;
	wire [16-1:0] node3747;
	wire [16-1:0] node3751;
	wire [16-1:0] node3752;
	wire [16-1:0] node3756;
	wire [16-1:0] node3757;
	wire [16-1:0] node3758;
	wire [16-1:0] node3759;
	wire [16-1:0] node3761;
	wire [16-1:0] node3764;
	wire [16-1:0] node3766;
	wire [16-1:0] node3769;
	wire [16-1:0] node3770;
	wire [16-1:0] node3774;
	wire [16-1:0] node3775;
	wire [16-1:0] node3776;
	wire [16-1:0] node3777;
	wire [16-1:0] node3781;
	wire [16-1:0] node3782;
	wire [16-1:0] node3783;
	wire [16-1:0] node3787;
	wire [16-1:0] node3788;
	wire [16-1:0] node3790;
	wire [16-1:0] node3794;
	wire [16-1:0] node3795;
	wire [16-1:0] node3796;
	wire [16-1:0] node3797;
	wire [16-1:0] node3799;
	wire [16-1:0] node3803;
	wire [16-1:0] node3804;
	wire [16-1:0] node3807;
	wire [16-1:0] node3810;
	wire [16-1:0] node3811;
	wire [16-1:0] node3813;
	wire [16-1:0] node3816;
	wire [16-1:0] node3818;
	wire [16-1:0] node3820;
	wire [16-1:0] node3823;
	wire [16-1:0] node3824;
	wire [16-1:0] node3825;
	wire [16-1:0] node3826;
	wire [16-1:0] node3827;
	wire [16-1:0] node3828;
	wire [16-1:0] node3830;
	wire [16-1:0] node3831;
	wire [16-1:0] node3835;
	wire [16-1:0] node3836;
	wire [16-1:0] node3840;
	wire [16-1:0] node3841;
	wire [16-1:0] node3844;
	wire [16-1:0] node3845;
	wire [16-1:0] node3846;
	wire [16-1:0] node3851;
	wire [16-1:0] node3852;
	wire [16-1:0] node3853;
	wire [16-1:0] node3856;
	wire [16-1:0] node3857;
	wire [16-1:0] node3858;
	wire [16-1:0] node3863;
	wire [16-1:0] node3864;
	wire [16-1:0] node3867;
	wire [16-1:0] node3870;
	wire [16-1:0] node3871;
	wire [16-1:0] node3872;
	wire [16-1:0] node3873;
	wire [16-1:0] node3877;
	wire [16-1:0] node3880;
	wire [16-1:0] node3881;
	wire [16-1:0] node3882;
	wire [16-1:0] node3884;
	wire [16-1:0] node3887;
	wire [16-1:0] node3888;
	wire [16-1:0] node3891;
	wire [16-1:0] node3893;
	wire [16-1:0] node3894;
	wire [16-1:0] node3898;
	wire [16-1:0] node3899;
	wire [16-1:0] node3900;
	wire [16-1:0] node3904;
	wire [16-1:0] node3905;
	wire [16-1:0] node3908;
	wire [16-1:0] node3911;
	wire [16-1:0] node3912;
	wire [16-1:0] node3913;
	wire [16-1:0] node3914;
	wire [16-1:0] node3916;
	wire [16-1:0] node3917;
	wire [16-1:0] node3921;
	wire [16-1:0] node3923;
	wire [16-1:0] node3925;
	wire [16-1:0] node3927;
	wire [16-1:0] node3929;
	wire [16-1:0] node3932;
	wire [16-1:0] node3933;
	wire [16-1:0] node3934;
	wire [16-1:0] node3938;
	wire [16-1:0] node3940;
	wire [16-1:0] node3941;
	wire [16-1:0] node3944;
	wire [16-1:0] node3947;
	wire [16-1:0] node3948;
	wire [16-1:0] node3949;
	wire [16-1:0] node3951;
	wire [16-1:0] node3954;
	wire [16-1:0] node3956;
	wire [16-1:0] node3959;
	wire [16-1:0] node3960;
	wire [16-1:0] node3962;
	wire [16-1:0] node3964;
	wire [16-1:0] node3967;
	wire [16-1:0] node3968;
	wire [16-1:0] node3970;
	wire [16-1:0] node3971;
	wire [16-1:0] node3975;
	wire [16-1:0] node3976;
	wire [16-1:0] node3979;
	wire [16-1:0] node3982;
	wire [16-1:0] node3983;
	wire [16-1:0] node3984;
	wire [16-1:0] node3985;
	wire [16-1:0] node3986;
	wire [16-1:0] node3987;
	wire [16-1:0] node3988;
	wire [16-1:0] node3990;
	wire [16-1:0] node3991;
	wire [16-1:0] node3995;
	wire [16-1:0] node3996;
	wire [16-1:0] node3998;
	wire [16-1:0] node4001;
	wire [16-1:0] node4003;
	wire [16-1:0] node4006;
	wire [16-1:0] node4007;
	wire [16-1:0] node4009;
	wire [16-1:0] node4010;
	wire [16-1:0] node4014;
	wire [16-1:0] node4015;
	wire [16-1:0] node4018;
	wire [16-1:0] node4021;
	wire [16-1:0] node4022;
	wire [16-1:0] node4023;
	wire [16-1:0] node4024;
	wire [16-1:0] node4028;
	wire [16-1:0] node4029;
	wire [16-1:0] node4031;
	wire [16-1:0] node4035;
	wire [16-1:0] node4036;
	wire [16-1:0] node4038;
	wire [16-1:0] node4039;
	wire [16-1:0] node4043;
	wire [16-1:0] node4044;
	wire [16-1:0] node4046;
	wire [16-1:0] node4050;
	wire [16-1:0] node4051;
	wire [16-1:0] node4052;
	wire [16-1:0] node4053;
	wire [16-1:0] node4054;
	wire [16-1:0] node4057;
	wire [16-1:0] node4061;
	wire [16-1:0] node4062;
	wire [16-1:0] node4063;
	wire [16-1:0] node4064;
	wire [16-1:0] node4069;
	wire [16-1:0] node4072;
	wire [16-1:0] node4073;
	wire [16-1:0] node4074;
	wire [16-1:0] node4075;
	wire [16-1:0] node4079;
	wire [16-1:0] node4080;
	wire [16-1:0] node4083;
	wire [16-1:0] node4085;
	wire [16-1:0] node4088;
	wire [16-1:0] node4089;
	wire [16-1:0] node4091;
	wire [16-1:0] node4092;
	wire [16-1:0] node4095;
	wire [16-1:0] node4096;
	wire [16-1:0] node4098;
	wire [16-1:0] node4102;
	wire [16-1:0] node4103;
	wire [16-1:0] node4104;
	wire [16-1:0] node4108;
	wire [16-1:0] node4111;
	wire [16-1:0] node4112;
	wire [16-1:0] node4113;
	wire [16-1:0] node4114;
	wire [16-1:0] node4115;
	wire [16-1:0] node4116;
	wire [16-1:0] node4117;
	wire [16-1:0] node4121;
	wire [16-1:0] node4124;
	wire [16-1:0] node4126;
	wire [16-1:0] node4127;
	wire [16-1:0] node4131;
	wire [16-1:0] node4132;
	wire [16-1:0] node4133;
	wire [16-1:0] node4134;
	wire [16-1:0] node4137;
	wire [16-1:0] node4141;
	wire [16-1:0] node4143;
	wire [16-1:0] node4146;
	wire [16-1:0] node4147;
	wire [16-1:0] node4148;
	wire [16-1:0] node4149;
	wire [16-1:0] node4152;
	wire [16-1:0] node4154;
	wire [16-1:0] node4155;
	wire [16-1:0] node4159;
	wire [16-1:0] node4160;
	wire [16-1:0] node4164;
	wire [16-1:0] node4165;
	wire [16-1:0] node4166;
	wire [16-1:0] node4167;
	wire [16-1:0] node4168;
	wire [16-1:0] node4173;
	wire [16-1:0] node4176;
	wire [16-1:0] node4177;
	wire [16-1:0] node4180;
	wire [16-1:0] node4183;
	wire [16-1:0] node4184;
	wire [16-1:0] node4185;
	wire [16-1:0] node4186;
	wire [16-1:0] node4188;
	wire [16-1:0] node4191;
	wire [16-1:0] node4194;
	wire [16-1:0] node4196;
	wire [16-1:0] node4197;
	wire [16-1:0] node4198;
	wire [16-1:0] node4201;
	wire [16-1:0] node4204;
	wire [16-1:0] node4205;
	wire [16-1:0] node4209;
	wire [16-1:0] node4210;
	wire [16-1:0] node4211;
	wire [16-1:0] node4214;
	wire [16-1:0] node4215;
	wire [16-1:0] node4219;
	wire [16-1:0] node4220;
	wire [16-1:0] node4221;
	wire [16-1:0] node4223;
	wire [16-1:0] node4226;
	wire [16-1:0] node4229;
	wire [16-1:0] node4230;
	wire [16-1:0] node4232;
	wire [16-1:0] node4233;
	wire [16-1:0] node4235;
	wire [16-1:0] node4239;
	wire [16-1:0] node4240;
	wire [16-1:0] node4243;
	wire [16-1:0] node4244;
	wire [16-1:0] node4246;
	wire [16-1:0] node4250;
	wire [16-1:0] node4251;
	wire [16-1:0] node4252;
	wire [16-1:0] node4253;
	wire [16-1:0] node4254;
	wire [16-1:0] node4255;
	wire [16-1:0] node4256;
	wire [16-1:0] node4257;
	wire [16-1:0] node4260;
	wire [16-1:0] node4264;
	wire [16-1:0] node4266;
	wire [16-1:0] node4268;
	wire [16-1:0] node4271;
	wire [16-1:0] node4272;
	wire [16-1:0] node4273;
	wire [16-1:0] node4277;
	wire [16-1:0] node4279;
	wire [16-1:0] node4282;
	wire [16-1:0] node4283;
	wire [16-1:0] node4284;
	wire [16-1:0] node4285;
	wire [16-1:0] node4288;
	wire [16-1:0] node4290;
	wire [16-1:0] node4293;
	wire [16-1:0] node4294;
	wire [16-1:0] node4297;
	wire [16-1:0] node4300;
	wire [16-1:0] node4301;
	wire [16-1:0] node4303;
	wire [16-1:0] node4306;
	wire [16-1:0] node4307;
	wire [16-1:0] node4311;
	wire [16-1:0] node4312;
	wire [16-1:0] node4313;
	wire [16-1:0] node4314;
	wire [16-1:0] node4315;
	wire [16-1:0] node4317;
	wire [16-1:0] node4320;
	wire [16-1:0] node4323;
	wire [16-1:0] node4325;
	wire [16-1:0] node4326;
	wire [16-1:0] node4330;
	wire [16-1:0] node4331;
	wire [16-1:0] node4332;
	wire [16-1:0] node4334;
	wire [16-1:0] node4338;
	wire [16-1:0] node4341;
	wire [16-1:0] node4342;
	wire [16-1:0] node4343;
	wire [16-1:0] node4346;
	wire [16-1:0] node4348;
	wire [16-1:0] node4351;
	wire [16-1:0] node4352;
	wire [16-1:0] node4353;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4359;
	wire [16-1:0] node4363;
	wire [16-1:0] node4365;
	wire [16-1:0] node4366;
	wire [16-1:0] node4369;
	wire [16-1:0] node4372;
	wire [16-1:0] node4373;
	wire [16-1:0] node4374;
	wire [16-1:0] node4375;
	wire [16-1:0] node4378;
	wire [16-1:0] node4379;
	wire [16-1:0] node4380;
	wire [16-1:0] node4383;
	wire [16-1:0] node4386;
	wire [16-1:0] node4389;
	wire [16-1:0] node4390;
	wire [16-1:0] node4392;
	wire [16-1:0] node4393;
	wire [16-1:0] node4397;
	wire [16-1:0] node4398;
	wire [16-1:0] node4399;
	wire [16-1:0] node4402;
	wire [16-1:0] node4405;
	wire [16-1:0] node4407;
	wire [16-1:0] node4409;
	wire [16-1:0] node4410;
	wire [16-1:0] node4414;
	wire [16-1:0] node4415;
	wire [16-1:0] node4416;
	wire [16-1:0] node4417;
	wire [16-1:0] node4420;
	wire [16-1:0] node4422;
	wire [16-1:0] node4425;
	wire [16-1:0] node4427;
	wire [16-1:0] node4428;
	wire [16-1:0] node4429;
	wire [16-1:0] node4431;
	wire [16-1:0] node4435;
	wire [16-1:0] node4438;
	wire [16-1:0] node4439;
	wire [16-1:0] node4440;
	wire [16-1:0] node4442;
	wire [16-1:0] node4443;
	wire [16-1:0] node4447;
	wire [16-1:0] node4450;
	wire [16-1:0] node4451;
	wire [16-1:0] node4452;
	wire [16-1:0] node4455;
	wire [16-1:0] node4456;
	wire [16-1:0] node4460;
	wire [16-1:0] node4462;

	assign outp = (inp[1]) ? node2282 : node1;
		assign node1 = (inp[4]) ? node1187 : node2;
			assign node2 = (inp[3]) ? node614 : node3;
				assign node3 = (inp[12]) ? node323 : node4;
					assign node4 = (inp[11]) ? node182 : node5;
						assign node5 = (inp[0]) ? node99 : node6;
							assign node6 = (inp[2]) ? node46 : node7;
								assign node7 = (inp[15]) ? node19 : node8;
									assign node8 = (inp[7]) ? node14 : node9;
										assign node9 = (inp[10]) ? 16'b0000011111111111 : node10;
											assign node10 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
										assign node14 = (inp[13]) ? node16 : 16'b0001111111111111;
											assign node16 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
									assign node19 = (inp[6]) ? node39 : node20;
										assign node20 = (inp[5]) ? node34 : node21;
											assign node21 = (inp[9]) ? node25 : node22;
												assign node22 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node25 = (inp[7]) ? node31 : node26;
													assign node26 = (inp[8]) ? 16'b0000111111111111 : node27;
														assign node27 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node31 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node34 = (inp[13]) ? node36 : 16'b0001111111111111;
												assign node36 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node39 = (inp[8]) ? node41 : 16'b0000111111111111;
											assign node41 = (inp[13]) ? 16'b0000011111111111 : node42;
												assign node42 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
								assign node46 = (inp[15]) ? node70 : node47;
									assign node47 = (inp[10]) ? node61 : node48;
										assign node48 = (inp[7]) ? 16'b0000011111111111 : node49;
											assign node49 = (inp[9]) ? node55 : node50;
												assign node50 = (inp[6]) ? 16'b0001111111111111 : node51;
													assign node51 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node55 = (inp[8]) ? node57 : 16'b0000111111111111;
													assign node57 = (inp[14]) ? 16'b0000011111111111 : 16'b0001111111111111;
										assign node61 = (inp[13]) ? 16'b0000001111111111 : node62;
											assign node62 = (inp[6]) ? node66 : node63;
												assign node63 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node66 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
									assign node70 = (inp[6]) ? node84 : node71;
										assign node71 = (inp[10]) ? 16'b0000001111111111 : node72;
											assign node72 = (inp[7]) ? node80 : node73;
												assign node73 = (inp[13]) ? 16'b0000011111111111 : node74;
													assign node74 = (inp[5]) ? 16'b0000111111111111 : node75;
														assign node75 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node80 = (inp[14]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node84 = (inp[14]) ? node90 : node85;
											assign node85 = (inp[5]) ? node87 : 16'b0000111111111111;
												assign node87 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node90 = (inp[9]) ? node92 : 16'b0000001111111111;
												assign node92 = (inp[5]) ? 16'b0000000011111111 : node93;
													assign node93 = (inp[7]) ? node95 : 16'b0000000111111111;
														assign node95 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node99 = (inp[6]) ? node129 : node100;
								assign node100 = (inp[13]) ? node120 : node101;
									assign node101 = (inp[8]) ? node111 : node102;
										assign node102 = (inp[14]) ? node106 : node103;
											assign node103 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node106 = (inp[9]) ? 16'b0000111111111111 : node107;
												assign node107 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
										assign node111 = (inp[14]) ? 16'b0000001111111111 : node112;
											assign node112 = (inp[9]) ? node116 : node113;
												assign node113 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node116 = (inp[10]) ? 16'b0000011111111111 : 16'b0000001111111111;
									assign node120 = (inp[5]) ? node126 : node121;
										assign node121 = (inp[10]) ? node123 : 16'b0000011111111111;
											assign node123 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node126 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
								assign node129 = (inp[8]) ? node155 : node130;
									assign node130 = (inp[5]) ? node144 : node131;
										assign node131 = (inp[9]) ? node137 : node132;
											assign node132 = (inp[7]) ? node134 : 16'b0001111111111111;
												assign node134 = (inp[14]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node137 = (inp[14]) ? 16'b0000001111111111 : node138;
												assign node138 = (inp[15]) ? node140 : 16'b0000011111111111;
													assign node140 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node144 = (inp[13]) ? node152 : node145;
											assign node145 = (inp[7]) ? node149 : node146;
												assign node146 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node149 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node152 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node155 = (inp[7]) ? node167 : node156;
										assign node156 = (inp[2]) ? node162 : node157;
											assign node157 = (inp[5]) ? node159 : 16'b0000000111111111;
												assign node159 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node162 = (inp[15]) ? 16'b0000001111111111 : node163;
												assign node163 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node167 = (inp[2]) ? node175 : node168;
											assign node168 = (inp[13]) ? 16'b0000000111111111 : node169;
												assign node169 = (inp[5]) ? node171 : 16'b0000001111111111;
													assign node171 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node175 = (inp[15]) ? node179 : node176;
												assign node176 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node179 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
						assign node182 = (inp[13]) ? node244 : node183;
							assign node183 = (inp[10]) ? node211 : node184;
								assign node184 = (inp[6]) ? node198 : node185;
									assign node185 = (inp[7]) ? node191 : node186;
										assign node186 = (inp[9]) ? 16'b0000011111111111 : node187;
											assign node187 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node191 = (inp[14]) ? node193 : 16'b0000111111111111;
											assign node193 = (inp[9]) ? 16'b0000001111111111 : node194;
												assign node194 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node198 = (inp[0]) ? node208 : node199;
										assign node199 = (inp[7]) ? node205 : node200;
											assign node200 = (inp[15]) ? node202 : 16'b0000111111111111;
												assign node202 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node205 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node208 = (inp[7]) ? 16'b0000001111111111 : 16'b0000000111111111;
								assign node211 = (inp[9]) ? node229 : node212;
									assign node212 = (inp[5]) ? node218 : node213;
										assign node213 = (inp[2]) ? node215 : 16'b0001111111111111;
											assign node215 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node218 = (inp[14]) ? node222 : node219;
											assign node219 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node222 = (inp[2]) ? node224 : 16'b0000001111111111;
												assign node224 = (inp[8]) ? node226 : 16'b0000000111111111;
													assign node226 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node229 = (inp[2]) ? node237 : node230;
										assign node230 = (inp[7]) ? node234 : node231;
											assign node231 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node234 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node237 = (inp[5]) ? 16'b0000000001111111 : node238;
											assign node238 = (inp[6]) ? node240 : 16'b0000000111111111;
												assign node240 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node244 = (inp[6]) ? node294 : node245;
								assign node245 = (inp[14]) ? node259 : node246;
									assign node246 = (inp[10]) ? node254 : node247;
										assign node247 = (inp[15]) ? 16'b0000001111111111 : node248;
											assign node248 = (inp[8]) ? 16'b0000011111111111 : node249;
												assign node249 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node254 = (inp[9]) ? node256 : 16'b0000001111111111;
											assign node256 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
									assign node259 = (inp[7]) ? node269 : node260;
										assign node260 = (inp[5]) ? 16'b0000001111111111 : node261;
											assign node261 = (inp[10]) ? 16'b0000001111111111 : node262;
												assign node262 = (inp[0]) ? node264 : 16'b0000011111111111;
													assign node264 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node269 = (inp[10]) ? node285 : node270;
											assign node270 = (inp[2]) ? node276 : node271;
												assign node271 = (inp[0]) ? node273 : 16'b0000011111111111;
													assign node273 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node276 = (inp[5]) ? node278 : 16'b0000000111111111;
													assign node278 = (inp[0]) ? node280 : 16'b0000000111111111;
														assign node280 = (inp[15]) ? 16'b0000000001111111 : node281;
															assign node281 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node285 = (inp[9]) ? node287 : 16'b0000000011111111;
												assign node287 = (inp[15]) ? 16'b0000000001111111 : node288;
													assign node288 = (inp[2]) ? 16'b0000000001111111 : node289;
														assign node289 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node294 = (inp[8]) ? node298 : node295;
									assign node295 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node298 = (inp[2]) ? node312 : node299;
										assign node299 = (inp[7]) ? node305 : node300;
											assign node300 = (inp[14]) ? 16'b0000000011111111 : node301;
												assign node301 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node305 = (inp[10]) ? node309 : node306;
												assign node306 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node309 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node312 = (inp[0]) ? node316 : node313;
											assign node313 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node316 = (inp[7]) ? 16'b0000000000011111 : node317;
												assign node317 = (inp[15]) ? node319 : 16'b0000000001111111;
													assign node319 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node323 = (inp[2]) ? node477 : node324;
						assign node324 = (inp[5]) ? node394 : node325;
							assign node325 = (inp[13]) ? node361 : node326;
								assign node326 = (inp[15]) ? node344 : node327;
									assign node327 = (inp[11]) ? node337 : node328;
										assign node328 = (inp[7]) ? node334 : node329;
											assign node329 = (inp[10]) ? node331 : 16'b0011111111111111;
												assign node331 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node334 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node337 = (inp[9]) ? 16'b0000001111111111 : node338;
											assign node338 = (inp[7]) ? node340 : 16'b0000011111111111;
												assign node340 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
									assign node344 = (inp[6]) ? node358 : node345;
										assign node345 = (inp[7]) ? node353 : node346;
											assign node346 = (inp[10]) ? 16'b0000011111111111 : node347;
												assign node347 = (inp[0]) ? node349 : 16'b0001111111111111;
													assign node349 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node353 = (inp[11]) ? node355 : 16'b0000011111111111;
												assign node355 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node358 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node361 = (inp[15]) ? node375 : node362;
									assign node362 = (inp[11]) ? node366 : node363;
										assign node363 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node366 = (inp[14]) ? node372 : node367;
											assign node367 = (inp[9]) ? 16'b0000000111111111 : node368;
												assign node368 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node372 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node375 = (inp[0]) ? node385 : node376;
										assign node376 = (inp[7]) ? node382 : node377;
											assign node377 = (inp[11]) ? 16'b0000001111111111 : node378;
												assign node378 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node382 = (inp[8]) ? 16'b0000000001111111 : 16'b0000001111111111;
										assign node385 = (inp[6]) ? node389 : node386;
											assign node386 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node389 = (inp[7]) ? node391 : 16'b0000000111111111;
												assign node391 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node394 = (inp[15]) ? node434 : node395;
								assign node395 = (inp[13]) ? node413 : node396;
									assign node396 = (inp[6]) ? node408 : node397;
										assign node397 = (inp[0]) ? node403 : node398;
											assign node398 = (inp[14]) ? node400 : 16'b0000011111111111;
												assign node400 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node403 = (inp[9]) ? 16'b0000001111111111 : node404;
												assign node404 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
										assign node408 = (inp[9]) ? node410 : 16'b0000001111111111;
											assign node410 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node413 = (inp[11]) ? node425 : node414;
										assign node414 = (inp[14]) ? node420 : node415;
											assign node415 = (inp[0]) ? node417 : 16'b0000001111111111;
												assign node417 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node420 = (inp[0]) ? 16'b0000000011111111 : node421;
												assign node421 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node425 = (inp[8]) ? node427 : 16'b0000000111111111;
											assign node427 = (inp[6]) ? 16'b0000000011111111 : node428;
												assign node428 = (inp[14]) ? 16'b0000000011111111 : node429;
													assign node429 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node434 = (inp[9]) ? node456 : node435;
									assign node435 = (inp[10]) ? node447 : node436;
										assign node436 = (inp[8]) ? node440 : node437;
											assign node437 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node440 = (inp[11]) ? 16'b0000000111111111 : node441;
												assign node441 = (inp[0]) ? 16'b0000000111111111 : node442;
													assign node442 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node447 = (inp[6]) ? node449 : 16'b0000011111111111;
											assign node449 = (inp[13]) ? node453 : node450;
												assign node450 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node453 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node456 = (inp[6]) ? node464 : node457;
										assign node457 = (inp[14]) ? node461 : node458;
											assign node458 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node461 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node464 = (inp[7]) ? node472 : node465;
											assign node465 = (inp[14]) ? 16'b0000000001111111 : node466;
												assign node466 = (inp[10]) ? node468 : 16'b0000001111111111;
													assign node468 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node472 = (inp[10]) ? node474 : 16'b0000000001111111;
												assign node474 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node477 = (inp[8]) ? node539 : node478;
							assign node478 = (inp[9]) ? node508 : node479;
								assign node479 = (inp[5]) ? node493 : node480;
									assign node480 = (inp[11]) ? node488 : node481;
										assign node481 = (inp[13]) ? 16'b0000001111111111 : node482;
											assign node482 = (inp[15]) ? node484 : 16'b0000011111111111;
												assign node484 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node488 = (inp[14]) ? 16'b0000001111111111 : node489;
											assign node489 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node493 = (inp[14]) ? node501 : node494;
										assign node494 = (inp[15]) ? 16'b0000000111111111 : node495;
											assign node495 = (inp[10]) ? 16'b0000000111111111 : node496;
												assign node496 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node501 = (inp[0]) ? node505 : node502;
											assign node502 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node505 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node508 = (inp[7]) ? node524 : node509;
									assign node509 = (inp[10]) ? node521 : node510;
										assign node510 = (inp[0]) ? node516 : node511;
											assign node511 = (inp[6]) ? node513 : 16'b0000001111111111;
												assign node513 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node516 = (inp[6]) ? node518 : 16'b0000000111111111;
												assign node518 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node521 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node524 = (inp[15]) ? node534 : node525;
										assign node525 = (inp[14]) ? node531 : node526;
											assign node526 = (inp[0]) ? 16'b0000000011111111 : node527;
												assign node527 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node531 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node534 = (inp[5]) ? 16'b0000000001111111 : node535;
											assign node535 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node539 = (inp[6]) ? node577 : node540;
								assign node540 = (inp[5]) ? node558 : node541;
									assign node541 = (inp[15]) ? node549 : node542;
										assign node542 = (inp[9]) ? 16'b0000000111111111 : node543;
											assign node543 = (inp[14]) ? node545 : 16'b0000001111111111;
												assign node545 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node549 = (inp[11]) ? node553 : node550;
											assign node550 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node553 = (inp[0]) ? 16'b0000000011111111 : node554;
												assign node554 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node558 = (inp[10]) ? node566 : node559;
										assign node559 = (inp[7]) ? node563 : node560;
											assign node560 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node563 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node566 = (inp[7]) ? node574 : node567;
											assign node567 = (inp[13]) ? node571 : node568;
												assign node568 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node571 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node574 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node577 = (inp[7]) ? node597 : node578;
									assign node578 = (inp[15]) ? node590 : node579;
										assign node579 = (inp[13]) ? node585 : node580;
											assign node580 = (inp[11]) ? node582 : 16'b0000000111111111;
												assign node582 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node585 = (inp[9]) ? 16'b0000000001111111 : node586;
												assign node586 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node590 = (inp[0]) ? node594 : node591;
											assign node591 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node594 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node597 = (inp[0]) ? node605 : node598;
										assign node598 = (inp[9]) ? node600 : 16'b0000000011111111;
											assign node600 = (inp[10]) ? node602 : 16'b0000000001111111;
												assign node602 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node605 = (inp[15]) ? node609 : node606;
											assign node606 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node609 = (inp[11]) ? node611 : 16'b0000000000111111;
												assign node611 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000001111;
				assign node614 = (inp[9]) ? node920 : node615;
					assign node615 = (inp[6]) ? node767 : node616;
						assign node616 = (inp[15]) ? node680 : node617;
							assign node617 = (inp[5]) ? node651 : node618;
								assign node618 = (inp[2]) ? node638 : node619;
									assign node619 = (inp[13]) ? node629 : node620;
										assign node620 = (inp[7]) ? node622 : 16'b0000111111111111;
											assign node622 = (inp[10]) ? 16'b0000011111111111 : node623;
												assign node623 = (inp[0]) ? node625 : 16'b0000111111111111;
													assign node625 = (inp[11]) ? 16'b0000111111111111 : 16'b0000011111111111;
										assign node629 = (inp[8]) ? node635 : node630;
											assign node630 = (inp[12]) ? 16'b0000011111111111 : node631;
												assign node631 = (inp[11]) ? 16'b0000011111111111 : 16'b0001111111111111;
											assign node635 = (inp[14]) ? 16'b0000011111111111 : 16'b0000001111111111;
									assign node638 = (inp[14]) ? node644 : node639;
										assign node639 = (inp[12]) ? 16'b0000001111111111 : node640;
											assign node640 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node644 = (inp[13]) ? node646 : 16'b0000011111111111;
											assign node646 = (inp[11]) ? 16'b0000000000111111 : node647;
												assign node647 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node651 = (inp[7]) ? node667 : node652;
									assign node652 = (inp[12]) ? 16'b0000001111111111 : node653;
										assign node653 = (inp[10]) ? node659 : node654;
											assign node654 = (inp[13]) ? node656 : 16'b0000011111111111;
												assign node656 = (inp[8]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node659 = (inp[14]) ? node663 : node660;
												assign node660 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node663 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node667 = (inp[2]) ? node675 : node668;
										assign node668 = (inp[12]) ? node672 : node669;
											assign node669 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node672 = (inp[0]) ? 16'b0000001111111111 : 16'b0000000011111111;
										assign node675 = (inp[11]) ? 16'b0000000111111111 : node676;
											assign node676 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node680 = (inp[14]) ? node730 : node681;
								assign node681 = (inp[5]) ? node713 : node682;
									assign node682 = (inp[10]) ? node696 : node683;
										assign node683 = (inp[11]) ? node691 : node684;
											assign node684 = (inp[13]) ? node686 : 16'b0000011111111111;
												assign node686 = (inp[8]) ? node688 : 16'b0000001111111111;
													assign node688 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node691 = (inp[12]) ? node693 : 16'b0000011111111111;
												assign node693 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node696 = (inp[13]) ? node708 : node697;
											assign node697 = (inp[11]) ? node701 : node698;
												assign node698 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node701 = (inp[8]) ? node703 : 16'b0000011111111111;
													assign node703 = (inp[0]) ? 16'b0000001111111111 : node704;
														assign node704 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node708 = (inp[12]) ? node710 : 16'b0000000111111111;
												assign node710 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node713 = (inp[2]) ? node719 : node714;
										assign node714 = (inp[0]) ? 16'b0000000111111111 : node715;
											assign node715 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node719 = (inp[11]) ? node723 : node720;
											assign node720 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node723 = (inp[7]) ? node727 : node724;
												assign node724 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node727 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000000111111;
								assign node730 = (inp[7]) ? node748 : node731;
									assign node731 = (inp[13]) ? node739 : node732;
										assign node732 = (inp[11]) ? 16'b0000000111111111 : node733;
											assign node733 = (inp[8]) ? 16'b0000000111111111 : node734;
												assign node734 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
										assign node739 = (inp[2]) ? node741 : 16'b0000000111111111;
											assign node741 = (inp[0]) ? 16'b0000000011111111 : node742;
												assign node742 = (inp[5]) ? node744 : 16'b0000000111111111;
													assign node744 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node748 = (inp[0]) ? node756 : node749;
										assign node749 = (inp[11]) ? 16'b0000000111111111 : node750;
											assign node750 = (inp[8]) ? node752 : 16'b0000000111111111;
												assign node752 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node756 = (inp[10]) ? node764 : node757;
											assign node757 = (inp[13]) ? 16'b0000000011111111 : node758;
												assign node758 = (inp[11]) ? node760 : 16'b0000000111111111;
													assign node760 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node764 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
						assign node767 = (inp[13]) ? node843 : node768;
							assign node768 = (inp[8]) ? node804 : node769;
								assign node769 = (inp[5]) ? node791 : node770;
									assign node770 = (inp[15]) ? node780 : node771;
										assign node771 = (inp[10]) ? 16'b0000001111111111 : node772;
											assign node772 = (inp[11]) ? node776 : node773;
												assign node773 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node776 = (inp[0]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node780 = (inp[10]) ? node788 : node781;
											assign node781 = (inp[11]) ? node783 : 16'b0000001111111111;
												assign node783 = (inp[2]) ? 16'b0000001111111111 : node784;
													assign node784 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node788 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node791 = (inp[14]) ? node801 : node792;
										assign node792 = (inp[15]) ? node796 : node793;
											assign node793 = (inp[11]) ? 16'b0000000111111111 : 16'b0001111111111111;
											assign node796 = (inp[11]) ? node798 : 16'b0000001111111111;
												assign node798 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node801 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
								assign node804 = (inp[10]) ? node818 : node805;
									assign node805 = (inp[15]) ? node809 : node806;
										assign node806 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node809 = (inp[14]) ? node811 : 16'b0000001111111111;
											assign node811 = (inp[7]) ? 16'b0000000011111111 : node812;
												assign node812 = (inp[2]) ? node814 : 16'b0000000111111111;
													assign node814 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node818 = (inp[0]) ? node832 : node819;
										assign node819 = (inp[11]) ? node829 : node820;
											assign node820 = (inp[2]) ? node824 : node821;
												assign node821 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node824 = (inp[7]) ? 16'b0000000011111111 : node825;
													assign node825 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node829 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node832 = (inp[15]) ? node838 : node833;
											assign node833 = (inp[12]) ? 16'b0000000011111111 : node834;
												assign node834 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node838 = (inp[12]) ? node840 : 16'b0000000011111111;
												assign node840 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node843 = (inp[5]) ? node889 : node844;
								assign node844 = (inp[15]) ? node856 : node845;
									assign node845 = (inp[7]) ? node851 : node846;
										assign node846 = (inp[14]) ? node848 : 16'b0000001111111111;
											assign node848 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node851 = (inp[2]) ? node853 : 16'b0000000111111111;
											assign node853 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node856 = (inp[11]) ? node872 : node857;
										assign node857 = (inp[10]) ? node863 : node858;
											assign node858 = (inp[14]) ? 16'b0000000001111111 : node859;
												assign node859 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node863 = (inp[2]) ? node865 : 16'b0000000011111111;
												assign node865 = (inp[0]) ? 16'b0000000011111111 : node866;
													assign node866 = (inp[7]) ? node868 : 16'b0000000111111111;
														assign node868 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node872 = (inp[10]) ? node878 : node873;
											assign node873 = (inp[0]) ? node875 : 16'b0000000011111111;
												assign node875 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node878 = (inp[0]) ? 16'b0000000000111111 : node879;
												assign node879 = (inp[14]) ? node885 : node880;
													assign node880 = (inp[2]) ? node882 : 16'b0000000011111111;
														assign node882 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node885 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node889 = (inp[0]) ? node903 : node890;
									assign node890 = (inp[11]) ? node896 : node891;
										assign node891 = (inp[12]) ? 16'b0000000001111111 : node892;
											assign node892 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node896 = (inp[8]) ? node898 : 16'b0000000011111111;
											assign node898 = (inp[15]) ? 16'b0000000011111111 : node899;
												assign node899 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node903 = (inp[14]) ? node911 : node904;
										assign node904 = (inp[10]) ? node908 : node905;
											assign node905 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node908 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node911 = (inp[8]) ? node913 : 16'b0000000001111111;
											assign node913 = (inp[2]) ? node915 : 16'b0000000000111111;
												assign node915 = (inp[7]) ? node917 : 16'b0000000000111111;
													assign node917 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node920 = (inp[10]) ? node1050 : node921;
						assign node921 = (inp[14]) ? node977 : node922;
							assign node922 = (inp[11]) ? node948 : node923;
								assign node923 = (inp[8]) ? node935 : node924;
									assign node924 = (inp[5]) ? node932 : node925;
										assign node925 = (inp[12]) ? 16'b0000001111111111 : node926;
											assign node926 = (inp[15]) ? node928 : 16'b0000111111111111;
												assign node928 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node932 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node935 = (inp[15]) ? node943 : node936;
										assign node936 = (inp[6]) ? 16'b0000000111111111 : node937;
											assign node937 = (inp[5]) ? node939 : 16'b0000001111111111;
												assign node939 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node943 = (inp[5]) ? node945 : 16'b0000000111111111;
											assign node945 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node948 = (inp[15]) ? node964 : node949;
									assign node949 = (inp[0]) ? node959 : node950;
										assign node950 = (inp[13]) ? node956 : node951;
											assign node951 = (inp[5]) ? 16'b0000001111111111 : node952;
												assign node952 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node956 = (inp[7]) ? 16'b0000011111111111 : 16'b0000000111111111;
										assign node959 = (inp[5]) ? node961 : 16'b0000001111111111;
											assign node961 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node964 = (inp[12]) ? node972 : node965;
										assign node965 = (inp[13]) ? node969 : node966;
											assign node966 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node969 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node972 = (inp[13]) ? 16'b0000000011111111 : node973;
											assign node973 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node977 = (inp[7]) ? node1015 : node978;
								assign node978 = (inp[15]) ? node998 : node979;
									assign node979 = (inp[13]) ? node987 : node980;
										assign node980 = (inp[0]) ? 16'b0000000111111111 : node981;
											assign node981 = (inp[12]) ? node983 : 16'b0000111111111111;
												assign node983 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node987 = (inp[2]) ? node991 : node988;
											assign node988 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node991 = (inp[5]) ? node993 : 16'b0000000111111111;
												assign node993 = (inp[6]) ? node995 : 16'b0000000011111111;
													assign node995 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node998 = (inp[0]) ? node1008 : node999;
										assign node999 = (inp[12]) ? 16'b0000000011111111 : node1000;
											assign node1000 = (inp[11]) ? node1004 : node1001;
												assign node1001 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1004 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1008 = (inp[13]) ? node1012 : node1009;
											assign node1009 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1012 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
								assign node1015 = (inp[2]) ? node1037 : node1016;
									assign node1016 = (inp[15]) ? node1024 : node1017;
										assign node1017 = (inp[8]) ? node1019 : 16'b0000000111111111;
											assign node1019 = (inp[6]) ? node1021 : 16'b0000000111111111;
												assign node1021 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1024 = (inp[8]) ? node1030 : node1025;
											assign node1025 = (inp[13]) ? 16'b0000000001111111 : node1026;
												assign node1026 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node1030 = (inp[5]) ? 16'b0000000000111111 : node1031;
												assign node1031 = (inp[11]) ? node1033 : 16'b0000000011111111;
													assign node1033 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1037 = (inp[6]) ? node1043 : node1038;
										assign node1038 = (inp[11]) ? 16'b0000000011111111 : node1039;
											assign node1039 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1043 = (inp[5]) ? node1045 : 16'b0000000001111111;
											assign node1045 = (inp[12]) ? node1047 : 16'b0000000000111111;
												assign node1047 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
						assign node1050 = (inp[14]) ? node1114 : node1051;
							assign node1051 = (inp[6]) ? node1075 : node1052;
								assign node1052 = (inp[8]) ? node1064 : node1053;
									assign node1053 = (inp[11]) ? node1055 : 16'b0000001111111111;
										assign node1055 = (inp[2]) ? node1061 : node1056;
											assign node1056 = (inp[5]) ? 16'b0000000111111111 : node1057;
												assign node1057 = (inp[13]) ? 16'b0000000011111111 : 16'b0000011111111111;
											assign node1061 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node1064 = (inp[15]) ? 16'b0000000011111111 : node1065;
										assign node1065 = (inp[5]) ? node1067 : 16'b0000001111111111;
											assign node1067 = (inp[0]) ? 16'b0000000011111111 : node1068;
												assign node1068 = (inp[11]) ? 16'b0000000111111111 : node1069;
													assign node1069 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1075 = (inp[8]) ? node1093 : node1076;
									assign node1076 = (inp[12]) ? node1088 : node1077;
										assign node1077 = (inp[5]) ? node1083 : node1078;
											assign node1078 = (inp[15]) ? node1080 : 16'b0000001111111111;
												assign node1080 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1083 = (inp[15]) ? node1085 : 16'b0000000111111111;
												assign node1085 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node1088 = (inp[2]) ? node1090 : 16'b0000000011111111;
											assign node1090 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1093 = (inp[5]) ? node1103 : node1094;
										assign node1094 = (inp[11]) ? node1098 : node1095;
											assign node1095 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1098 = (inp[2]) ? node1100 : 16'b0000000001111111;
												assign node1100 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1103 = (inp[0]) ? node1111 : node1104;
											assign node1104 = (inp[11]) ? node1106 : 16'b0000000001111111;
												assign node1106 = (inp[7]) ? node1108 : 16'b0000000001111111;
													assign node1108 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node1111 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1114 = (inp[11]) ? node1146 : node1115;
								assign node1115 = (inp[6]) ? node1131 : node1116;
									assign node1116 = (inp[2]) ? node1122 : node1117;
										assign node1117 = (inp[8]) ? node1119 : 16'b0000000011111111;
											assign node1119 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1122 = (inp[8]) ? 16'b0000000001111111 : node1123;
											assign node1123 = (inp[7]) ? node1125 : 16'b0000000111111111;
												assign node1125 = (inp[5]) ? node1127 : 16'b0000000011111111;
													assign node1127 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1131 = (inp[5]) ? node1139 : node1132;
										assign node1132 = (inp[13]) ? 16'b0000000001111111 : node1133;
											assign node1133 = (inp[15]) ? 16'b0000000001111111 : node1134;
												assign node1134 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1139 = (inp[2]) ? 16'b0000000001111111 : node1140;
											assign node1140 = (inp[15]) ? 16'b0000000000111111 : node1141;
												assign node1141 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node1146 = (inp[7]) ? node1164 : node1147;
									assign node1147 = (inp[5]) ? node1155 : node1148;
										assign node1148 = (inp[13]) ? node1150 : 16'b0000000111111111;
											assign node1150 = (inp[15]) ? node1152 : 16'b0000000011111111;
												assign node1152 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1155 = (inp[6]) ? 16'b0000000011111111 : node1156;
											assign node1156 = (inp[12]) ? 16'b0000000001111111 : node1157;
												assign node1157 = (inp[13]) ? node1159 : 16'b0000000001111111;
													assign node1159 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1164 = (inp[13]) ? node1174 : node1165;
										assign node1165 = (inp[6]) ? node1169 : node1166;
											assign node1166 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1169 = (inp[2]) ? 16'b0000000000001111 : node1170;
												assign node1170 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node1174 = (inp[5]) ? node1182 : node1175;
											assign node1175 = (inp[12]) ? node1179 : node1176;
												assign node1176 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1179 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node1182 = (inp[0]) ? node1184 : 16'b0000000000111111;
												assign node1184 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
			assign node1187 = (inp[10]) ? node1733 : node1188;
				assign node1188 = (inp[3]) ? node1476 : node1189;
					assign node1189 = (inp[13]) ? node1325 : node1190;
						assign node1190 = (inp[15]) ? node1264 : node1191;
							assign node1191 = (inp[11]) ? node1223 : node1192;
								assign node1192 = (inp[6]) ? node1212 : node1193;
									assign node1193 = (inp[12]) ? node1203 : node1194;
										assign node1194 = (inp[8]) ? node1196 : 16'b0000111111111111;
											assign node1196 = (inp[7]) ? node1198 : 16'b0000111111111111;
												assign node1198 = (inp[14]) ? node1200 : 16'b0000011111111111;
													assign node1200 = (inp[5]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node1203 = (inp[14]) ? node1207 : node1204;
											assign node1204 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1207 = (inp[0]) ? node1209 : 16'b0000011111111111;
												assign node1209 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node1212 = (inp[14]) ? node1216 : node1213;
										assign node1213 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1216 = (inp[0]) ? 16'b0000000111111111 : node1217;
											assign node1217 = (inp[12]) ? 16'b0000000111111111 : node1218;
												assign node1218 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
								assign node1223 = (inp[9]) ? node1245 : node1224;
									assign node1224 = (inp[6]) ? node1232 : node1225;
										assign node1225 = (inp[2]) ? 16'b0000001111111111 : node1226;
											assign node1226 = (inp[0]) ? 16'b0000011111111111 : node1227;
												assign node1227 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node1232 = (inp[0]) ? 16'b0000000111111111 : node1233;
											assign node1233 = (inp[12]) ? node1239 : node1234;
												assign node1234 = (inp[5]) ? node1236 : 16'b0000011111111111;
													assign node1236 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1239 = (inp[7]) ? 16'b0000001111111111 : node1240;
													assign node1240 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1245 = (inp[2]) ? node1257 : node1246;
										assign node1246 = (inp[8]) ? node1248 : 16'b0000001111111111;
											assign node1248 = (inp[12]) ? node1252 : node1249;
												assign node1249 = (inp[7]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node1252 = (inp[5]) ? node1254 : 16'b0000000011111111;
													assign node1254 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1257 = (inp[7]) ? node1261 : node1258;
											assign node1258 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1261 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1264 = (inp[7]) ? node1294 : node1265;
								assign node1265 = (inp[12]) ? node1275 : node1266;
									assign node1266 = (inp[5]) ? 16'b0000000111111111 : node1267;
										assign node1267 = (inp[11]) ? 16'b0000001111111111 : node1268;
											assign node1268 = (inp[0]) ? 16'b0000011111111111 : node1269;
												assign node1269 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
									assign node1275 = (inp[8]) ? node1287 : node1276;
										assign node1276 = (inp[11]) ? node1282 : node1277;
											assign node1277 = (inp[5]) ? 16'b0000001111111111 : node1278;
												assign node1278 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1282 = (inp[5]) ? 16'b0000000011111111 : node1283;
												assign node1283 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1287 = (inp[2]) ? 16'b0000000011111111 : node1288;
											assign node1288 = (inp[0]) ? node1290 : 16'b0000001111111111;
												assign node1290 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1294 = (inp[5]) ? node1312 : node1295;
									assign node1295 = (inp[6]) ? node1303 : node1296;
										assign node1296 = (inp[8]) ? node1298 : 16'b0000000111111111;
											assign node1298 = (inp[0]) ? node1300 : 16'b0000011111111111;
												assign node1300 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1303 = (inp[2]) ? node1307 : node1304;
											assign node1304 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1307 = (inp[9]) ? node1309 : 16'b0000000011111111;
												assign node1309 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1312 = (inp[11]) ? node1322 : node1313;
										assign node1313 = (inp[8]) ? node1315 : 16'b0000000011111111;
											assign node1315 = (inp[2]) ? 16'b0000000001111111 : node1316;
												assign node1316 = (inp[14]) ? node1318 : 16'b0000000011111111;
													assign node1318 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1322 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000111111111;
						assign node1325 = (inp[14]) ? node1397 : node1326;
							assign node1326 = (inp[7]) ? node1366 : node1327;
								assign node1327 = (inp[0]) ? node1349 : node1328;
									assign node1328 = (inp[8]) ? node1340 : node1329;
										assign node1329 = (inp[9]) ? node1333 : node1330;
											assign node1330 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1333 = (inp[12]) ? 16'b0000001111111111 : node1334;
												assign node1334 = (inp[6]) ? node1336 : 16'b0000011111111111;
													assign node1336 = (inp[11]) ? 16'b0000000111111111 : 16'b0000111111111111;
										assign node1340 = (inp[5]) ? node1346 : node1341;
											assign node1341 = (inp[15]) ? node1343 : 16'b0000011111111111;
												assign node1343 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1346 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1349 = (inp[2]) ? node1361 : node1350;
										assign node1350 = (inp[8]) ? node1356 : node1351;
											assign node1351 = (inp[9]) ? node1353 : 16'b0000011111111111;
												assign node1353 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1356 = (inp[6]) ? 16'b0000000011111111 : node1357;
												assign node1357 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node1361 = (inp[8]) ? 16'b0000000001111111 : node1362;
											assign node1362 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1366 = (inp[15]) ? node1380 : node1367;
									assign node1367 = (inp[6]) ? node1377 : node1368;
										assign node1368 = (inp[8]) ? node1372 : node1369;
											assign node1369 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1372 = (inp[0]) ? node1374 : 16'b0000011111111111;
												assign node1374 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node1377 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000001111111;
									assign node1380 = (inp[12]) ? node1390 : node1381;
										assign node1381 = (inp[5]) ? node1385 : node1382;
											assign node1382 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1385 = (inp[8]) ? node1387 : 16'b0000000001111111;
												assign node1387 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1390 = (inp[8]) ? node1394 : node1391;
											assign node1391 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node1394 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1397 = (inp[6]) ? node1427 : node1398;
								assign node1398 = (inp[0]) ? node1408 : node1399;
									assign node1399 = (inp[15]) ? 16'b0000000011111111 : node1400;
										assign node1400 = (inp[12]) ? node1404 : node1401;
											assign node1401 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node1404 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1408 = (inp[7]) ? node1420 : node1409;
										assign node1409 = (inp[5]) ? node1415 : node1410;
											assign node1410 = (inp[9]) ? node1412 : 16'b0000000111111111;
												assign node1412 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1415 = (inp[9]) ? 16'b0000000011111111 : node1416;
												assign node1416 = (inp[12]) ? 16'b0000000011111111 : 16'b0000011111111111;
										assign node1420 = (inp[9]) ? node1422 : 16'b0000000011111111;
											assign node1422 = (inp[12]) ? node1424 : 16'b0000000011111111;
												assign node1424 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1427 = (inp[0]) ? node1449 : node1428;
									assign node1428 = (inp[8]) ? node1442 : node1429;
										assign node1429 = (inp[5]) ? node1437 : node1430;
											assign node1430 = (inp[11]) ? 16'b0000000111111111 : node1431;
												assign node1431 = (inp[7]) ? 16'b0000000111111111 : node1432;
													assign node1432 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1437 = (inp[2]) ? node1439 : 16'b0000000001111111;
												assign node1439 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node1442 = (inp[11]) ? node1444 : 16'b0000000000111111;
											assign node1444 = (inp[9]) ? node1446 : 16'b0000000001111111;
												assign node1446 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1449 = (inp[7]) ? node1461 : node1450;
										assign node1450 = (inp[8]) ? node1456 : node1451;
											assign node1451 = (inp[2]) ? node1453 : 16'b0000000011111111;
												assign node1453 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1456 = (inp[2]) ? node1458 : 16'b0000000001111111;
												assign node1458 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1461 = (inp[5]) ? node1471 : node1462;
											assign node1462 = (inp[12]) ? node1466 : node1463;
												assign node1463 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1466 = (inp[15]) ? 16'b0000000000011111 : node1467;
													assign node1467 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1471 = (inp[11]) ? 16'b0000000000011111 : node1472;
												assign node1472 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node1476 = (inp[13]) ? node1634 : node1477;
						assign node1477 = (inp[2]) ? node1559 : node1478;
							assign node1478 = (inp[12]) ? node1520 : node1479;
								assign node1479 = (inp[9]) ? node1497 : node1480;
									assign node1480 = (inp[15]) ? node1492 : node1481;
										assign node1481 = (inp[14]) ? node1485 : node1482;
											assign node1482 = (inp[5]) ? 16'b0000011111111111 : 16'b0001111111111111;
											assign node1485 = (inp[11]) ? 16'b0000000111111111 : node1486;
												assign node1486 = (inp[5]) ? node1488 : 16'b0000011111111111;
													assign node1488 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1492 = (inp[11]) ? 16'b0000000111111111 : node1493;
											assign node1493 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1497 = (inp[0]) ? node1511 : node1498;
										assign node1498 = (inp[8]) ? node1502 : node1499;
											assign node1499 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node1502 = (inp[11]) ? node1508 : node1503;
												assign node1503 = (inp[14]) ? 16'b0000000111111111 : node1504;
													assign node1504 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1508 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1511 = (inp[14]) ? 16'b0000000011111111 : node1512;
											assign node1512 = (inp[5]) ? 16'b0000000111111111 : node1513;
												assign node1513 = (inp[11]) ? node1515 : 16'b0000000111111111;
													assign node1515 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1520 = (inp[14]) ? node1544 : node1521;
									assign node1521 = (inp[5]) ? node1533 : node1522;
										assign node1522 = (inp[15]) ? node1524 : 16'b0000001111111111;
											assign node1524 = (inp[6]) ? node1528 : node1525;
												assign node1525 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1528 = (inp[11]) ? 16'b0000000111111111 : node1529;
													assign node1529 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node1533 = (inp[9]) ? 16'b0000000011111111 : node1534;
											assign node1534 = (inp[11]) ? node1536 : 16'b0000000111111111;
												assign node1536 = (inp[7]) ? node1538 : 16'b0000000111111111;
													assign node1538 = (inp[0]) ? node1540 : 16'b0000000011111111;
														assign node1540 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1544 = (inp[8]) ? node1552 : node1545;
										assign node1545 = (inp[15]) ? node1549 : node1546;
											assign node1546 = (inp[6]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node1549 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1552 = (inp[11]) ? 16'b0000000001111111 : node1553;
											assign node1553 = (inp[9]) ? 16'b0000000001111111 : node1554;
												assign node1554 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1559 = (inp[5]) ? node1595 : node1560;
								assign node1560 = (inp[11]) ? node1580 : node1561;
									assign node1561 = (inp[14]) ? node1573 : node1562;
										assign node1562 = (inp[6]) ? node1566 : node1563;
											assign node1563 = (inp[12]) ? 16'b0000000111111111 : 16'b0000111111111111;
											assign node1566 = (inp[0]) ? 16'b0000001111111111 : node1567;
												assign node1567 = (inp[12]) ? 16'b0000001111111111 : node1568;
													assign node1568 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1573 = (inp[6]) ? node1577 : node1574;
											assign node1574 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1577 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1580 = (inp[0]) ? node1584 : node1581;
										assign node1581 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1584 = (inp[7]) ? node1592 : node1585;
											assign node1585 = (inp[15]) ? node1587 : 16'b0000000011111111;
												assign node1587 = (inp[14]) ? node1589 : 16'b0000000001111111;
													assign node1589 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1592 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1595 = (inp[9]) ? node1615 : node1596;
									assign node1596 = (inp[11]) ? node1602 : node1597;
										assign node1597 = (inp[15]) ? node1599 : 16'b0000000111111111;
											assign node1599 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1602 = (inp[7]) ? node1608 : node1603;
											assign node1603 = (inp[0]) ? 16'b0000000001111111 : node1604;
												assign node1604 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1608 = (inp[6]) ? node1612 : node1609;
												assign node1609 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1612 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1615 = (inp[7]) ? node1621 : node1616;
										assign node1616 = (inp[11]) ? node1618 : 16'b0000000011111111;
											assign node1618 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node1621 = (inp[15]) ? node1627 : node1622;
											assign node1622 = (inp[8]) ? 16'b0000000000111111 : node1623;
												assign node1623 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node1627 = (inp[8]) ? node1629 : 16'b0000000000111111;
												assign node1629 = (inp[0]) ? 16'b0000000000011111 : node1630;
													assign node1630 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1634 = (inp[7]) ? node1676 : node1635;
							assign node1635 = (inp[8]) ? node1651 : node1636;
								assign node1636 = (inp[15]) ? node1642 : node1637;
									assign node1637 = (inp[0]) ? node1639 : 16'b0000001111111111;
										assign node1639 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
									assign node1642 = (inp[6]) ? 16'b0000000001111111 : node1643;
										assign node1643 = (inp[5]) ? node1645 : 16'b0000000111111111;
											assign node1645 = (inp[9]) ? node1647 : 16'b0000000111111111;
												assign node1647 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1651 = (inp[5]) ? node1667 : node1652;
									assign node1652 = (inp[11]) ? node1660 : node1653;
										assign node1653 = (inp[12]) ? node1655 : 16'b0000000111111111;
											assign node1655 = (inp[6]) ? 16'b0000000001111111 : node1656;
												assign node1656 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1660 = (inp[0]) ? 16'b0000000001111111 : node1661;
											assign node1661 = (inp[12]) ? node1663 : 16'b0000000011111111;
												assign node1663 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1667 = (inp[0]) ? node1673 : node1668;
										assign node1668 = (inp[15]) ? 16'b0000000001111111 : node1669;
											assign node1669 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1673 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1676 = (inp[5]) ? node1712 : node1677;
								assign node1677 = (inp[2]) ? node1691 : node1678;
									assign node1678 = (inp[6]) ? node1686 : node1679;
										assign node1679 = (inp[14]) ? 16'b0000000011111111 : node1680;
											assign node1680 = (inp[9]) ? 16'b0000000111111111 : node1681;
												assign node1681 = (inp[12]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node1686 = (inp[8]) ? node1688 : 16'b0000000011111111;
											assign node1688 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1691 = (inp[12]) ? node1705 : node1692;
										assign node1692 = (inp[15]) ? node1700 : node1693;
											assign node1693 = (inp[0]) ? 16'b0000000001111111 : node1694;
												assign node1694 = (inp[6]) ? 16'b0000000011111111 : node1695;
													assign node1695 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1700 = (inp[0]) ? node1702 : 16'b0000000001111111;
												assign node1702 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1705 = (inp[9]) ? node1707 : 16'b0000000001111111;
											assign node1707 = (inp[14]) ? 16'b0000000000011111 : node1708;
												assign node1708 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1712 = (inp[0]) ? node1722 : node1713;
									assign node1713 = (inp[14]) ? node1719 : node1714;
										assign node1714 = (inp[8]) ? 16'b0000000001111111 : node1715;
											assign node1715 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1719 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node1722 = (inp[2]) ? node1728 : node1723;
										assign node1723 = (inp[11]) ? 16'b0000000000111111 : node1724;
											assign node1724 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1728 = (inp[8]) ? 16'b0000000000001111 : node1729;
											assign node1729 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
				assign node1733 = (inp[6]) ? node2003 : node1734;
					assign node1734 = (inp[15]) ? node1864 : node1735;
						assign node1735 = (inp[8]) ? node1807 : node1736;
							assign node1736 = (inp[14]) ? node1772 : node1737;
								assign node1737 = (inp[0]) ? node1759 : node1738;
									assign node1738 = (inp[5]) ? node1750 : node1739;
										assign node1739 = (inp[12]) ? node1743 : node1740;
											assign node1740 = (inp[2]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node1743 = (inp[7]) ? 16'b0000000111111111 : node1744;
												assign node1744 = (inp[9]) ? node1746 : 16'b0000011111111111;
													assign node1746 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1750 = (inp[2]) ? node1756 : node1751;
											assign node1751 = (inp[3]) ? 16'b0000001111111111 : node1752;
												assign node1752 = (inp[12]) ? 16'b0000111111111111 : 16'b0000001111111111;
											assign node1756 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1759 = (inp[11]) ? node1763 : node1760;
										assign node1760 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1763 = (inp[13]) ? node1769 : node1764;
											assign node1764 = (inp[12]) ? 16'b0000001111111111 : node1765;
												assign node1765 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node1769 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1772 = (inp[11]) ? node1788 : node1773;
									assign node1773 = (inp[2]) ? node1783 : node1774;
										assign node1774 = (inp[0]) ? node1778 : node1775;
											assign node1775 = (inp[13]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node1778 = (inp[3]) ? node1780 : 16'b0000001111111111;
												assign node1780 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1783 = (inp[7]) ? 16'b0000000011111111 : node1784;
											assign node1784 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node1788 = (inp[3]) ? node1796 : node1789;
										assign node1789 = (inp[7]) ? 16'b0000000011111111 : node1790;
											assign node1790 = (inp[12]) ? 16'b0000000111111111 : node1791;
												assign node1791 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node1796 = (inp[0]) ? node1804 : node1797;
											assign node1797 = (inp[7]) ? node1799 : 16'b0000000111111111;
												assign node1799 = (inp[5]) ? 16'b0000000011111111 : node1800;
													assign node1800 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1804 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1807 = (inp[9]) ? node1841 : node1808;
								assign node1808 = (inp[2]) ? node1828 : node1809;
									assign node1809 = (inp[12]) ? node1817 : node1810;
										assign node1810 = (inp[0]) ? 16'b0000000111111111 : node1811;
											assign node1811 = (inp[3]) ? node1813 : 16'b0000011111111111;
												assign node1813 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1817 = (inp[13]) ? 16'b0000000011111111 : node1818;
											assign node1818 = (inp[7]) ? node1820 : 16'b0000000111111111;
												assign node1820 = (inp[11]) ? node1822 : 16'b0000000111111111;
													assign node1822 = (inp[3]) ? 16'b0000000011111111 : node1823;
														assign node1823 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1828 = (inp[5]) ? node1836 : node1829;
										assign node1829 = (inp[7]) ? node1831 : 16'b0000001111111111;
											assign node1831 = (inp[13]) ? node1833 : 16'b0000000111111111;
												assign node1833 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node1836 = (inp[3]) ? 16'b0000000001111111 : node1837;
											assign node1837 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1841 = (inp[11]) ? node1853 : node1842;
									assign node1842 = (inp[5]) ? node1844 : 16'b0000000011111111;
										assign node1844 = (inp[0]) ? 16'b0000000011111111 : node1845;
											assign node1845 = (inp[13]) ? node1847 : 16'b0000000111111111;
												assign node1847 = (inp[14]) ? 16'b0000000001111111 : node1848;
													assign node1848 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1853 = (inp[5]) ? node1861 : node1854;
										assign node1854 = (inp[12]) ? node1856 : 16'b0000000011111111;
											assign node1856 = (inp[0]) ? 16'b0000000000111111 : node1857;
												assign node1857 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1861 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node1864 = (inp[8]) ? node1936 : node1865;
							assign node1865 = (inp[5]) ? node1897 : node1866;
								assign node1866 = (inp[9]) ? node1886 : node1867;
									assign node1867 = (inp[12]) ? node1883 : node1868;
										assign node1868 = (inp[11]) ? node1874 : node1869;
											assign node1869 = (inp[13]) ? 16'b0000001111111111 : node1870;
												assign node1870 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1874 = (inp[14]) ? node1880 : node1875;
												assign node1875 = (inp[3]) ? node1877 : 16'b0000001111111111;
													assign node1877 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1880 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node1883 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1886 = (inp[0]) ? node1894 : node1887;
										assign node1887 = (inp[2]) ? node1889 : 16'b0000000111111111;
											assign node1889 = (inp[14]) ? 16'b0000000011111111 : node1890;
												assign node1890 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1894 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1897 = (inp[7]) ? node1921 : node1898;
									assign node1898 = (inp[14]) ? node1908 : node1899;
										assign node1899 = (inp[3]) ? node1903 : node1900;
											assign node1900 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1903 = (inp[12]) ? node1905 : 16'b0000000111111111;
												assign node1905 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1908 = (inp[13]) ? node1916 : node1909;
											assign node1909 = (inp[11]) ? node1911 : 16'b0000000011111111;
												assign node1911 = (inp[2]) ? 16'b0000000001111111 : node1912;
													assign node1912 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1916 = (inp[9]) ? node1918 : 16'b0000000011111111;
												assign node1918 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node1921 = (inp[13]) ? node1925 : node1922;
										assign node1922 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1925 = (inp[2]) ? node1927 : 16'b0000000011111111;
											assign node1927 = (inp[11]) ? node1929 : 16'b0000000001111111;
												assign node1929 = (inp[0]) ? 16'b0000000000011111 : node1930;
													assign node1930 = (inp[12]) ? node1932 : 16'b0000000000111111;
														assign node1932 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1936 = (inp[3]) ? node1972 : node1937;
								assign node1937 = (inp[7]) ? node1957 : node1938;
									assign node1938 = (inp[0]) ? node1946 : node1939;
										assign node1939 = (inp[5]) ? 16'b0000001111111111 : node1940;
											assign node1940 = (inp[14]) ? node1942 : 16'b0000000111111111;
												assign node1942 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1946 = (inp[13]) ? node1950 : node1947;
											assign node1947 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node1950 = (inp[9]) ? node1952 : 16'b0000000011111111;
												assign node1952 = (inp[12]) ? node1954 : 16'b0000000001111111;
													assign node1954 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1957 = (inp[5]) ? node1963 : node1958;
										assign node1958 = (inp[2]) ? node1960 : 16'b0000000011111111;
											assign node1960 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1963 = (inp[2]) ? node1965 : 16'b0000000000111111;
											assign node1965 = (inp[13]) ? node1969 : node1966;
												assign node1966 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node1969 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000011111;
								assign node1972 = (inp[5]) ? node1986 : node1973;
									assign node1973 = (inp[0]) ? node1981 : node1974;
										assign node1974 = (inp[9]) ? node1978 : node1975;
											assign node1975 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1978 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1981 = (inp[7]) ? 16'b0000000000111111 : node1982;
											assign node1982 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node1986 = (inp[14]) ? node1994 : node1987;
										assign node1987 = (inp[7]) ? 16'b0000000000001111 : node1988;
											assign node1988 = (inp[11]) ? 16'b0000000000111111 : node1989;
												assign node1989 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1994 = (inp[9]) ? node1998 : node1995;
											assign node1995 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node1998 = (inp[11]) ? node2000 : 16'b0000000000011111;
												assign node2000 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node2003 = (inp[11]) ? node2149 : node2004;
						assign node2004 = (inp[15]) ? node2068 : node2005;
							assign node2005 = (inp[2]) ? node2041 : node2006;
								assign node2006 = (inp[3]) ? node2022 : node2007;
									assign node2007 = (inp[7]) ? node2019 : node2008;
										assign node2008 = (inp[5]) ? node2014 : node2009;
											assign node2009 = (inp[12]) ? 16'b0000001111111111 : node2010;
												assign node2010 = (inp[13]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node2014 = (inp[9]) ? node2016 : 16'b0000000011111111;
												assign node2016 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2019 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2022 = (inp[5]) ? node2034 : node2023;
										assign node2023 = (inp[12]) ? node2029 : node2024;
											assign node2024 = (inp[0]) ? node2026 : 16'b0000001111111111;
												assign node2026 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2029 = (inp[7]) ? node2031 : 16'b0000000111111111;
												assign node2031 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2034 = (inp[0]) ? node2036 : 16'b0000000011111111;
											assign node2036 = (inp[14]) ? 16'b0000000000011111 : node2037;
												assign node2037 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node2041 = (inp[12]) ? node2053 : node2042;
									assign node2042 = (inp[9]) ? node2044 : 16'b0000001111111111;
										assign node2044 = (inp[14]) ? node2048 : node2045;
											assign node2045 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2048 = (inp[5]) ? 16'b0000000001111111 : node2049;
												assign node2049 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2053 = (inp[8]) ? node2063 : node2054;
										assign node2054 = (inp[7]) ? node2060 : node2055;
											assign node2055 = (inp[14]) ? node2057 : 16'b0000000011111111;
												assign node2057 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2060 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node2063 = (inp[0]) ? node2065 : 16'b0000000001111111;
											assign node2065 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node2068 = (inp[0]) ? node2104 : node2069;
								assign node2069 = (inp[13]) ? node2087 : node2070;
									assign node2070 = (inp[7]) ? node2078 : node2071;
										assign node2071 = (inp[14]) ? node2073 : 16'b0000000111111111;
											assign node2073 = (inp[5]) ? node2075 : 16'b0000000011111111;
												assign node2075 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node2078 = (inp[12]) ? node2080 : 16'b0000000011111111;
											assign node2080 = (inp[2]) ? node2084 : node2081;
												assign node2081 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node2084 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2087 = (inp[3]) ? node2091 : node2088;
										assign node2088 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node2091 = (inp[12]) ? node2093 : 16'b0000000001111111;
											assign node2093 = (inp[14]) ? node2101 : node2094;
												assign node2094 = (inp[7]) ? node2096 : 16'b0000000001111111;
													assign node2096 = (inp[5]) ? 16'b0000000000111111 : node2097;
														assign node2097 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2101 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node2104 = (inp[9]) ? node2130 : node2105;
									assign node2105 = (inp[14]) ? node2113 : node2106;
										assign node2106 = (inp[13]) ? node2108 : 16'b0000000111111111;
											assign node2108 = (inp[7]) ? 16'b0000000001111111 : node2109;
												assign node2109 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2113 = (inp[12]) ? 16'b0000000000011111 : node2114;
											assign node2114 = (inp[8]) ? node2124 : node2115;
												assign node2115 = (inp[2]) ? node2119 : node2116;
													assign node2116 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2119 = (inp[5]) ? node2121 : 16'b0000000001111111;
														assign node2121 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2124 = (inp[7]) ? 16'b0000000000001111 : node2125;
													assign node2125 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2130 = (inp[12]) ? node2140 : node2131;
										assign node2131 = (inp[2]) ? node2137 : node2132;
											assign node2132 = (inp[3]) ? node2134 : 16'b0000000011111111;
												assign node2134 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node2137 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node2140 = (inp[14]) ? node2142 : 16'b0000000000111111;
											assign node2142 = (inp[2]) ? 16'b0000000000011111 : node2143;
												assign node2143 = (inp[7]) ? 16'b0000000000111111 : node2144;
													assign node2144 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
						assign node2149 = (inp[14]) ? node2225 : node2150;
							assign node2150 = (inp[5]) ? node2194 : node2151;
								assign node2151 = (inp[2]) ? node2167 : node2152;
									assign node2152 = (inp[9]) ? node2160 : node2153;
										assign node2153 = (inp[0]) ? node2155 : 16'b0000000111111111;
											assign node2155 = (inp[3]) ? node2157 : 16'b0000000111111111;
												assign node2157 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2160 = (inp[8]) ? node2162 : 16'b0000000011111111;
											assign node2162 = (inp[3]) ? 16'b0000000001111111 : node2163;
												assign node2163 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2167 = (inp[3]) ? node2175 : node2168;
										assign node2168 = (inp[7]) ? node2170 : 16'b0000000011111111;
											assign node2170 = (inp[12]) ? node2172 : 16'b0000000001111111;
												assign node2172 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2175 = (inp[12]) ? node2177 : 16'b0000000001111111;
											assign node2177 = (inp[7]) ? node2189 : node2178;
												assign node2178 = (inp[13]) ? node2182 : node2179;
													assign node2179 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2182 = (inp[8]) ? 16'b0000000000111111 : node2183;
														assign node2183 = (inp[0]) ? 16'b0000000000111111 : node2184;
															assign node2184 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2189 = (inp[0]) ? node2191 : 16'b0000000000111111;
													assign node2191 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node2194 = (inp[9]) ? node2212 : node2195;
									assign node2195 = (inp[0]) ? node2205 : node2196;
										assign node2196 = (inp[8]) ? node2200 : node2197;
											assign node2197 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2200 = (inp[7]) ? 16'b0000000011111111 : node2201;
												assign node2201 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2205 = (inp[13]) ? node2209 : node2206;
											assign node2206 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node2209 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2212 = (inp[13]) ? node2222 : node2213;
										assign node2213 = (inp[0]) ? node2215 : 16'b0000000000111111;
											assign node2215 = (inp[2]) ? 16'b0000000000011111 : node2216;
												assign node2216 = (inp[7]) ? 16'b0000000001111111 : node2217;
													assign node2217 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2222 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000111111;
							assign node2225 = (inp[2]) ? node2249 : node2226;
								assign node2226 = (inp[13]) ? node2238 : node2227;
									assign node2227 = (inp[9]) ? node2231 : node2228;
										assign node2228 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2231 = (inp[0]) ? 16'b0000000000111111 : node2232;
											assign node2232 = (inp[8]) ? node2234 : 16'b0000000001111111;
												assign node2234 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2238 = (inp[3]) ? node2246 : node2239;
										assign node2239 = (inp[5]) ? node2243 : node2240;
											assign node2240 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node2243 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2246 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000000111;
								assign node2249 = (inp[15]) ? node2263 : node2250;
									assign node2250 = (inp[8]) ? node2254 : node2251;
										assign node2251 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2254 = (inp[12]) ? 16'b0000000000011111 : node2255;
											assign node2255 = (inp[0]) ? node2257 : 16'b0000000000111111;
												assign node2257 = (inp[7]) ? 16'b0000000000001111 : node2258;
													assign node2258 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2263 = (inp[8]) ? node2269 : node2264;
										assign node2264 = (inp[3]) ? node2266 : 16'b0000000001111111;
											assign node2266 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node2269 = (inp[7]) ? node2273 : node2270;
											assign node2270 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000000111;
											assign node2273 = (inp[5]) ? node2277 : node2274;
												assign node2274 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node2277 = (inp[12]) ? node2279 : 16'b0000000000000111;
													assign node2279 = (inp[0]) ? 16'b0000000000000011 : 16'b0000000000000111;
		assign node2282 = (inp[8]) ? node3446 : node2283;
			assign node2283 = (inp[14]) ? node2867 : node2284;
				assign node2284 = (inp[6]) ? node2582 : node2285;
					assign node2285 = (inp[13]) ? node2443 : node2286;
						assign node2286 = (inp[7]) ? node2374 : node2287;
							assign node2287 = (inp[5]) ? node2335 : node2288;
								assign node2288 = (inp[4]) ? node2306 : node2289;
									assign node2289 = (inp[15]) ? node2297 : node2290;
										assign node2290 = (inp[2]) ? 16'b0000011111111111 : node2291;
											assign node2291 = (inp[10]) ? 16'b0000111111111111 : node2292;
												assign node2292 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
										assign node2297 = (inp[10]) ? node2301 : node2298;
											assign node2298 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2301 = (inp[12]) ? node2303 : 16'b0000011111111111;
												assign node2303 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node2306 = (inp[11]) ? node2324 : node2307;
										assign node2307 = (inp[12]) ? node2315 : node2308;
											assign node2308 = (inp[2]) ? node2312 : node2309;
												assign node2309 = (inp[9]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node2312 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2315 = (inp[15]) ? 16'b0000001111111111 : node2316;
												assign node2316 = (inp[9]) ? node2318 : 16'b0000111111111111;
													assign node2318 = (inp[0]) ? 16'b0000001111111111 : node2319;
														assign node2319 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2324 = (inp[9]) ? node2332 : node2325;
											assign node2325 = (inp[0]) ? node2329 : node2326;
												assign node2326 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2329 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2332 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node2335 = (inp[12]) ? node2357 : node2336;
									assign node2336 = (inp[9]) ? node2346 : node2337;
										assign node2337 = (inp[4]) ? node2343 : node2338;
											assign node2338 = (inp[11]) ? node2340 : 16'b0000011111111111;
												assign node2340 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2343 = (inp[2]) ? 16'b0000000011111111 : 16'b0000011111111111;
										assign node2346 = (inp[3]) ? node2352 : node2347;
											assign node2347 = (inp[10]) ? 16'b0000001111111111 : node2348;
												assign node2348 = (inp[11]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node2352 = (inp[4]) ? 16'b0000000001111111 : node2353;
												assign node2353 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node2357 = (inp[10]) ? node2365 : node2358;
										assign node2358 = (inp[15]) ? node2360 : 16'b0000011111111111;
											assign node2360 = (inp[0]) ? node2362 : 16'b0000011111111111;
												assign node2362 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2365 = (inp[15]) ? node2369 : node2366;
											assign node2366 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2369 = (inp[11]) ? node2371 : 16'b0000000011111111;
												assign node2371 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
							assign node2374 = (inp[0]) ? node2422 : node2375;
								assign node2375 = (inp[9]) ? node2397 : node2376;
									assign node2376 = (inp[2]) ? node2386 : node2377;
										assign node2377 = (inp[11]) ? node2381 : node2378;
											assign node2378 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2381 = (inp[3]) ? node2383 : 16'b0000011111111111;
												assign node2383 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2386 = (inp[4]) ? node2394 : node2387;
											assign node2387 = (inp[10]) ? node2391 : node2388;
												assign node2388 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2391 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2394 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2397 = (inp[15]) ? node2411 : node2398;
										assign node2398 = (inp[12]) ? node2404 : node2399;
											assign node2399 = (inp[4]) ? 16'b0000001111111111 : node2400;
												assign node2400 = (inp[10]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node2404 = (inp[11]) ? node2408 : node2405;
												assign node2405 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2408 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2411 = (inp[11]) ? node2417 : node2412;
											assign node2412 = (inp[12]) ? node2414 : 16'b0000111111111111;
												assign node2414 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node2417 = (inp[4]) ? node2419 : 16'b0000000011111111;
												assign node2419 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2422 = (inp[12]) ? node2430 : node2423;
									assign node2423 = (inp[5]) ? node2427 : node2424;
										assign node2424 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2427 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node2430 = (inp[10]) ? node2434 : node2431;
										assign node2431 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2434 = (inp[9]) ? node2440 : node2435;
											assign node2435 = (inp[5]) ? node2437 : 16'b0000000011111111;
												assign node2437 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2440 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node2443 = (inp[10]) ? node2507 : node2444;
							assign node2444 = (inp[9]) ? node2484 : node2445;
								assign node2445 = (inp[15]) ? node2467 : node2446;
									assign node2446 = (inp[7]) ? node2456 : node2447;
										assign node2447 = (inp[2]) ? node2451 : node2448;
											assign node2448 = (inp[11]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node2451 = (inp[11]) ? 16'b0000001111111111 : node2452;
												assign node2452 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2456 = (inp[12]) ? node2462 : node2457;
											assign node2457 = (inp[4]) ? node2459 : 16'b0000001111111111;
												assign node2459 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2462 = (inp[4]) ? node2464 : 16'b0000000011111111;
												assign node2464 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node2467 = (inp[2]) ? node2481 : node2468;
										assign node2468 = (inp[0]) ? node2476 : node2469;
											assign node2469 = (inp[4]) ? 16'b0000000111111111 : node2470;
												assign node2470 = (inp[7]) ? 16'b0000001111111111 : node2471;
													assign node2471 = (inp[3]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node2476 = (inp[11]) ? node2478 : 16'b0000000111111111;
												assign node2478 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2481 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000000111111;
								assign node2484 = (inp[15]) ? node2494 : node2485;
									assign node2485 = (inp[5]) ? node2489 : node2486;
										assign node2486 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node2489 = (inp[12]) ? 16'b0000000011111111 : node2490;
											assign node2490 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2494 = (inp[3]) ? node2504 : node2495;
										assign node2495 = (inp[7]) ? node2501 : node2496;
											assign node2496 = (inp[11]) ? node2498 : 16'b0000000111111111;
												assign node2498 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2501 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2504 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
							assign node2507 = (inp[11]) ? node2555 : node2508;
								assign node2508 = (inp[0]) ? node2532 : node2509;
									assign node2509 = (inp[3]) ? node2519 : node2510;
										assign node2510 = (inp[15]) ? node2514 : node2511;
											assign node2511 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2514 = (inp[9]) ? node2516 : 16'b0000001111111111;
												assign node2516 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2519 = (inp[12]) ? node2525 : node2520;
											assign node2520 = (inp[9]) ? 16'b0000000111111111 : node2521;
												assign node2521 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2525 = (inp[9]) ? node2529 : node2526;
												assign node2526 = (inp[7]) ? 16'b0000001111111111 : 16'b0000000011111111;
												assign node2529 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2532 = (inp[3]) ? node2550 : node2533;
										assign node2533 = (inp[9]) ? node2535 : 16'b0000000111111111;
											assign node2535 = (inp[15]) ? node2547 : node2536;
												assign node2536 = (inp[2]) ? node2538 : 16'b0000000111111111;
													assign node2538 = (inp[7]) ? 16'b0000000011111111 : node2539;
														assign node2539 = (inp[12]) ? 16'b0000000011111111 : node2540;
															assign node2540 = (inp[5]) ? node2542 : 16'b0000000111111111;
																assign node2542 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2547 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2550 = (inp[5]) ? 16'b0000000011111111 : node2551;
											assign node2551 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
								assign node2555 = (inp[2]) ? node2569 : node2556;
									assign node2556 = (inp[0]) ? node2562 : node2557;
										assign node2557 = (inp[4]) ? 16'b0000000011111111 : node2558;
											assign node2558 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2562 = (inp[3]) ? node2564 : 16'b0000000011111111;
											assign node2564 = (inp[7]) ? 16'b0000000000111111 : node2565;
												assign node2565 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node2569 = (inp[7]) ? node2575 : node2570;
										assign node2570 = (inp[5]) ? 16'b0000000001111111 : node2571;
											assign node2571 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node2575 = (inp[4]) ? 16'b0000000000111111 : node2576;
											assign node2576 = (inp[15]) ? 16'b0000000000111111 : node2577;
												assign node2577 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
					assign node2582 = (inp[5]) ? node2740 : node2583;
						assign node2583 = (inp[10]) ? node2649 : node2584;
							assign node2584 = (inp[3]) ? node2616 : node2585;
								assign node2585 = (inp[11]) ? node2601 : node2586;
									assign node2586 = (inp[9]) ? node2596 : node2587;
										assign node2587 = (inp[15]) ? node2593 : node2588;
											assign node2588 = (inp[13]) ? 16'b0000011111111111 : node2589;
												assign node2589 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2593 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node2596 = (inp[12]) ? 16'b0000000111111111 : node2597;
											assign node2597 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
									assign node2601 = (inp[15]) ? node2611 : node2602;
										assign node2602 = (inp[4]) ? 16'b0000000111111111 : node2603;
											assign node2603 = (inp[0]) ? node2607 : node2604;
												assign node2604 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2607 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2611 = (inp[7]) ? node2613 : 16'b0000000001111111;
											assign node2613 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node2616 = (inp[15]) ? node2638 : node2617;
									assign node2617 = (inp[0]) ? node2625 : node2618;
										assign node2618 = (inp[4]) ? node2620 : 16'b0000001111111111;
											assign node2620 = (inp[9]) ? node2622 : 16'b0000000111111111;
												assign node2622 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2625 = (inp[13]) ? node2629 : node2626;
											assign node2626 = (inp[9]) ? 16'b0000000111111111 : 16'b0000111111111111;
											assign node2629 = (inp[9]) ? node2635 : node2630;
												assign node2630 = (inp[11]) ? 16'b0000000111111111 : node2631;
													assign node2631 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2635 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2638 = (inp[13]) ? node2644 : node2639;
										assign node2639 = (inp[9]) ? 16'b0000000001111111 : node2640;
											assign node2640 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2644 = (inp[4]) ? node2646 : 16'b0000000011111111;
											assign node2646 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
							assign node2649 = (inp[4]) ? node2691 : node2650;
								assign node2650 = (inp[9]) ? node2668 : node2651;
									assign node2651 = (inp[15]) ? node2659 : node2652;
										assign node2652 = (inp[2]) ? 16'b0000000111111111 : node2653;
											assign node2653 = (inp[0]) ? node2655 : 16'b0000000111111111;
												assign node2655 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2659 = (inp[3]) ? node2661 : 16'b0000000111111111;
											assign node2661 = (inp[0]) ? 16'b0000000011111111 : node2662;
												assign node2662 = (inp[12]) ? node2664 : 16'b0000000111111111;
													assign node2664 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2668 = (inp[3]) ? node2686 : node2669;
										assign node2669 = (inp[0]) ? node2677 : node2670;
											assign node2670 = (inp[13]) ? 16'b0000001111111111 : node2671;
												assign node2671 = (inp[11]) ? 16'b0000001111111111 : node2672;
													assign node2672 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2677 = (inp[7]) ? node2681 : node2678;
												assign node2678 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2681 = (inp[11]) ? 16'b0000000000111111 : node2682;
													assign node2682 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2686 = (inp[15]) ? 16'b0000000000111111 : node2687;
											assign node2687 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node2691 = (inp[13]) ? node2723 : node2692;
									assign node2692 = (inp[15]) ? node2702 : node2693;
										assign node2693 = (inp[9]) ? node2697 : node2694;
											assign node2694 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node2697 = (inp[3]) ? 16'b0000000011111111 : node2698;
												assign node2698 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2702 = (inp[7]) ? node2716 : node2703;
											assign node2703 = (inp[0]) ? node2711 : node2704;
												assign node2704 = (inp[12]) ? 16'b0000000011111111 : node2705;
													assign node2705 = (inp[11]) ? 16'b0000000111111111 : node2706;
														assign node2706 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2711 = (inp[11]) ? node2713 : 16'b0000000011111111;
													assign node2713 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2716 = (inp[9]) ? 16'b0000000011111111 : node2717;
												assign node2717 = (inp[2]) ? 16'b0000000001111111 : node2718;
													assign node2718 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2723 = (inp[7]) ? node2731 : node2724;
										assign node2724 = (inp[3]) ? 16'b0000000001111111 : node2725;
											assign node2725 = (inp[9]) ? node2727 : 16'b0000000111111111;
												assign node2727 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2731 = (inp[2]) ? node2735 : node2732;
											assign node2732 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2735 = (inp[12]) ? 16'b0000000000011111 : node2736;
												assign node2736 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node2740 = (inp[11]) ? node2800 : node2741;
							assign node2741 = (inp[7]) ? node2769 : node2742;
								assign node2742 = (inp[4]) ? node2756 : node2743;
									assign node2743 = (inp[12]) ? node2753 : node2744;
										assign node2744 = (inp[3]) ? node2750 : node2745;
											assign node2745 = (inp[9]) ? 16'b0000001111111111 : node2746;
												assign node2746 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2750 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2753 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2756 = (inp[13]) ? node2766 : node2757;
										assign node2757 = (inp[9]) ? 16'b0000000011111111 : node2758;
											assign node2758 = (inp[0]) ? node2762 : node2759;
												assign node2759 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2762 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node2766 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2769 = (inp[3]) ? node2791 : node2770;
									assign node2770 = (inp[0]) ? node2782 : node2771;
										assign node2771 = (inp[12]) ? node2777 : node2772;
											assign node2772 = (inp[10]) ? 16'b0000000111111111 : node2773;
												assign node2773 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2777 = (inp[4]) ? 16'b0000000011111111 : node2778;
												assign node2778 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2782 = (inp[4]) ? 16'b0000000000111111 : node2783;
											assign node2783 = (inp[12]) ? node2785 : 16'b0000000011111111;
												assign node2785 = (inp[15]) ? node2787 : 16'b0000000011111111;
													assign node2787 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2791 = (inp[10]) ? node2793 : 16'b0000000011111111;
										assign node2793 = (inp[9]) ? node2795 : 16'b0000000001111111;
											assign node2795 = (inp[2]) ? 16'b0000000000111111 : node2796;
												assign node2796 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
							assign node2800 = (inp[9]) ? node2830 : node2801;
								assign node2801 = (inp[0]) ? node2819 : node2802;
									assign node2802 = (inp[4]) ? node2810 : node2803;
										assign node2803 = (inp[3]) ? node2807 : node2804;
											assign node2804 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2807 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2810 = (inp[7]) ? 16'b0000000001111111 : node2811;
											assign node2811 = (inp[2]) ? 16'b0000000001111111 : node2812;
												assign node2812 = (inp[15]) ? node2814 : 16'b0000000111111111;
													assign node2814 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node2819 = (inp[4]) ? node2825 : node2820;
										assign node2820 = (inp[10]) ? 16'b0000000001111111 : node2821;
											assign node2821 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2825 = (inp[15]) ? node2827 : 16'b0000000001111111;
											assign node2827 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node2830 = (inp[13]) ? node2858 : node2831;
									assign node2831 = (inp[15]) ? node2843 : node2832;
										assign node2832 = (inp[12]) ? node2836 : node2833;
											assign node2833 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2836 = (inp[0]) ? node2840 : node2837;
												assign node2837 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2840 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2843 = (inp[3]) ? node2849 : node2844;
											assign node2844 = (inp[7]) ? 16'b0000000011111111 : node2845;
												assign node2845 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2849 = (inp[4]) ? 16'b0000000000011111 : node2850;
												assign node2850 = (inp[2]) ? node2854 : node2851;
													assign node2851 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2854 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2858 = (inp[2]) ? node2860 : 16'b0000000000111111;
										assign node2860 = (inp[15]) ? node2862 : 16'b0000000000111111;
											assign node2862 = (inp[3]) ? 16'b0000000000001111 : node2863;
												assign node2863 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
				assign node2867 = (inp[3]) ? node3145 : node2868;
					assign node2868 = (inp[13]) ? node3034 : node2869;
						assign node2869 = (inp[5]) ? node2947 : node2870;
							assign node2870 = (inp[4]) ? node2910 : node2871;
								assign node2871 = (inp[12]) ? node2895 : node2872;
									assign node2872 = (inp[6]) ? node2884 : node2873;
										assign node2873 = (inp[7]) ? node2879 : node2874;
											assign node2874 = (inp[2]) ? 16'b0000111111111111 : node2875;
												assign node2875 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node2879 = (inp[11]) ? node2881 : 16'b0000011111111111;
												assign node2881 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2884 = (inp[9]) ? node2890 : node2885;
											assign node2885 = (inp[0]) ? 16'b0000001111111111 : node2886;
												assign node2886 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node2890 = (inp[7]) ? node2892 : 16'b0000000011111111;
												assign node2892 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2895 = (inp[7]) ? node2903 : node2896;
										assign node2896 = (inp[15]) ? node2898 : 16'b0000001111111111;
											assign node2898 = (inp[10]) ? node2900 : 16'b0000001111111111;
												assign node2900 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node2903 = (inp[11]) ? 16'b0000000111111111 : node2904;
											assign node2904 = (inp[10]) ? 16'b0000000111111111 : node2905;
												assign node2905 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
								assign node2910 = (inp[7]) ? node2932 : node2911;
									assign node2911 = (inp[2]) ? node2929 : node2912;
										assign node2912 = (inp[9]) ? node2920 : node2913;
											assign node2913 = (inp[15]) ? node2915 : 16'b0000111111111111;
												assign node2915 = (inp[6]) ? node2917 : 16'b0000001111111111;
													assign node2917 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2920 = (inp[0]) ? 16'b0000000111111111 : node2921;
												assign node2921 = (inp[12]) ? node2923 : 16'b0000001111111111;
													assign node2923 = (inp[6]) ? 16'b0000000111111111 : node2924;
														assign node2924 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2929 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node2932 = (inp[9]) ? node2942 : node2933;
										assign node2933 = (inp[12]) ? node2937 : node2934;
											assign node2934 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2937 = (inp[6]) ? 16'b0000000111111111 : node2938;
												assign node2938 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2942 = (inp[6]) ? node2944 : 16'b0000000011111111;
											assign node2944 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
							assign node2947 = (inp[6]) ? node2991 : node2948;
								assign node2948 = (inp[0]) ? node2968 : node2949;
									assign node2949 = (inp[15]) ? node2963 : node2950;
										assign node2950 = (inp[11]) ? node2956 : node2951;
											assign node2951 = (inp[2]) ? 16'b0000001111111111 : node2952;
												assign node2952 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2956 = (inp[9]) ? node2958 : 16'b0000001111111111;
												assign node2958 = (inp[10]) ? 16'b0000000011111111 : node2959;
													assign node2959 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node2963 = (inp[7]) ? node2965 : 16'b0000001111111111;
											assign node2965 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node2968 = (inp[9]) ? node2976 : node2969;
										assign node2969 = (inp[7]) ? 16'b0000000011111111 : node2970;
											assign node2970 = (inp[10]) ? node2972 : 16'b0000000111111111;
												assign node2972 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2976 = (inp[10]) ? node2986 : node2977;
											assign node2977 = (inp[4]) ? node2983 : node2978;
												assign node2978 = (inp[12]) ? 16'b0000000011111111 : node2979;
													assign node2979 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node2983 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2986 = (inp[4]) ? 16'b0000000000111111 : node2987;
												assign node2987 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2991 = (inp[11]) ? node3009 : node2992;
									assign node2992 = (inp[4]) ? node3000 : node2993;
										assign node2993 = (inp[9]) ? 16'b0000000011111111 : node2994;
											assign node2994 = (inp[12]) ? node2996 : 16'b0000000111111111;
												assign node2996 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node3000 = (inp[7]) ? node3004 : node3001;
											assign node3001 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3004 = (inp[12]) ? node3006 : 16'b0000000011111111;
												assign node3006 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3009 = (inp[12]) ? node3019 : node3010;
										assign node3010 = (inp[7]) ? node3014 : node3011;
											assign node3011 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3014 = (inp[2]) ? node3016 : 16'b0000000111111111;
												assign node3016 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3019 = (inp[15]) ? node3025 : node3020;
											assign node3020 = (inp[9]) ? node3022 : 16'b0000000011111111;
												assign node3022 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3025 = (inp[9]) ? node3029 : node3026;
												assign node3026 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node3029 = (inp[0]) ? node3031 : 16'b0000000000011111;
													assign node3031 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node3034 = (inp[0]) ? node3098 : node3035;
							assign node3035 = (inp[12]) ? node3069 : node3036;
								assign node3036 = (inp[6]) ? node3052 : node3037;
									assign node3037 = (inp[7]) ? node3045 : node3038;
										assign node3038 = (inp[4]) ? node3040 : 16'b0000001111111111;
											assign node3040 = (inp[9]) ? 16'b0000001111111111 : node3041;
												assign node3041 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node3045 = (inp[4]) ? node3049 : node3046;
											assign node3046 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node3049 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3052 = (inp[10]) ? node3064 : node3053;
										assign node3053 = (inp[2]) ? node3059 : node3054;
											assign node3054 = (inp[11]) ? 16'b0000000011111111 : node3055;
												assign node3055 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3059 = (inp[11]) ? node3061 : 16'b0000000011111111;
												assign node3061 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3064 = (inp[5]) ? node3066 : 16'b0000000111111111;
											assign node3066 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3069 = (inp[5]) ? node3083 : node3070;
									assign node3070 = (inp[7]) ? node3078 : node3071;
										assign node3071 = (inp[15]) ? node3073 : 16'b0000000111111111;
											assign node3073 = (inp[11]) ? 16'b0000000011111111 : node3074;
												assign node3074 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3078 = (inp[9]) ? node3080 : 16'b0000000011111111;
											assign node3080 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3083 = (inp[2]) ? node3089 : node3084;
										assign node3084 = (inp[15]) ? 16'b0000000001111111 : node3085;
											assign node3085 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3089 = (inp[10]) ? node3095 : node3090;
											assign node3090 = (inp[15]) ? node3092 : 16'b0000000001111111;
												assign node3092 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node3095 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000011111;
							assign node3098 = (inp[4]) ? node3124 : node3099;
								assign node3099 = (inp[2]) ? node3113 : node3100;
									assign node3100 = (inp[10]) ? node3106 : node3101;
										assign node3101 = (inp[5]) ? node3103 : 16'b0000000111111111;
											assign node3103 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3106 = (inp[7]) ? 16'b0000000000111111 : node3107;
											assign node3107 = (inp[6]) ? node3109 : 16'b0000000011111111;
												assign node3109 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3113 = (inp[15]) ? node3117 : node3114;
										assign node3114 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node3117 = (inp[6]) ? node3119 : 16'b0000000000011111;
											assign node3119 = (inp[9]) ? node3121 : 16'b0000000000111111;
												assign node3121 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3124 = (inp[7]) ? node3132 : node3125;
									assign node3125 = (inp[12]) ? 16'b0000000000011111 : node3126;
										assign node3126 = (inp[2]) ? node3128 : 16'b0000000001111111;
											assign node3128 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node3132 = (inp[2]) ? node3140 : node3133;
										assign node3133 = (inp[5]) ? 16'b0000000000011111 : node3134;
											assign node3134 = (inp[15]) ? node3136 : 16'b0000000000111111;
												assign node3136 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3140 = (inp[11]) ? node3142 : 16'b0000000000011111;
											assign node3142 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node3145 = (inp[15]) ? node3287 : node3146;
						assign node3146 = (inp[12]) ? node3214 : node3147;
							assign node3147 = (inp[5]) ? node3183 : node3148;
								assign node3148 = (inp[2]) ? node3162 : node3149;
									assign node3149 = (inp[10]) ? node3157 : node3150;
										assign node3150 = (inp[9]) ? 16'b0000000111111111 : node3151;
											assign node3151 = (inp[13]) ? node3153 : 16'b0000001111111111;
												assign node3153 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node3157 = (inp[7]) ? node3159 : 16'b0000000111111111;
											assign node3159 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3162 = (inp[11]) ? node3172 : node3163;
										assign node3163 = (inp[4]) ? node3167 : node3164;
											assign node3164 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3167 = (inp[6]) ? 16'b0000000011111111 : node3168;
												assign node3168 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3172 = (inp[7]) ? node3180 : node3173;
											assign node3173 = (inp[9]) ? node3177 : node3174;
												assign node3174 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3177 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3180 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3183 = (inp[10]) ? node3201 : node3184;
									assign node3184 = (inp[13]) ? node3196 : node3185;
										assign node3185 = (inp[6]) ? node3191 : node3186;
											assign node3186 = (inp[4]) ? 16'b0000000111111111 : node3187;
												assign node3187 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3191 = (inp[11]) ? 16'b0000000001111111 : node3192;
												assign node3192 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3196 = (inp[9]) ? node3198 : 16'b0000000011111111;
											assign node3198 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3201 = (inp[4]) ? node3207 : node3202;
										assign node3202 = (inp[6]) ? 16'b0000000001111111 : node3203;
											assign node3203 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node3207 = (inp[7]) ? node3211 : node3208;
											assign node3208 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node3211 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node3214 = (inp[2]) ? node3248 : node3215;
								assign node3215 = (inp[6]) ? node3233 : node3216;
									assign node3216 = (inp[5]) ? node3226 : node3217;
										assign node3217 = (inp[9]) ? node3221 : node3218;
											assign node3218 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3221 = (inp[7]) ? node3223 : 16'b0000000111111111;
												assign node3223 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3226 = (inp[11]) ? node3228 : 16'b0000000011111111;
											assign node3228 = (inp[10]) ? 16'b0000000001111111 : node3229;
												assign node3229 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3233 = (inp[4]) ? node3243 : node3234;
										assign node3234 = (inp[7]) ? node3238 : node3235;
											assign node3235 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node3238 = (inp[9]) ? 16'b0000000000111111 : node3239;
												assign node3239 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3243 = (inp[0]) ? node3245 : 16'b0000000001111111;
											assign node3245 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node3248 = (inp[11]) ? node3262 : node3249;
									assign node3249 = (inp[4]) ? node3257 : node3250;
										assign node3250 = (inp[9]) ? 16'b0000000011111111 : node3251;
											assign node3251 = (inp[0]) ? node3253 : 16'b0000000011111111;
												assign node3253 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3257 = (inp[13]) ? node3259 : 16'b0000000001111111;
											assign node3259 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3262 = (inp[9]) ? node3280 : node3263;
										assign node3263 = (inp[7]) ? node3273 : node3264;
											assign node3264 = (inp[13]) ? node3266 : 16'b0000000001111111;
												assign node3266 = (inp[0]) ? 16'b0000000000111111 : node3267;
													assign node3267 = (inp[4]) ? node3269 : 16'b0000000001111111;
														assign node3269 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3273 = (inp[5]) ? 16'b0000000000011111 : node3274;
												assign node3274 = (inp[10]) ? node3276 : 16'b0000000000111111;
													assign node3276 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3280 = (inp[4]) ? 16'b0000000000000111 : node3281;
											assign node3281 = (inp[0]) ? 16'b0000000000011111 : node3282;
												assign node3282 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node3287 = (inp[12]) ? node3361 : node3288;
							assign node3288 = (inp[7]) ? node3312 : node3289;
								assign node3289 = (inp[0]) ? node3303 : node3290;
									assign node3290 = (inp[2]) ? node3292 : 16'b0000000011111111;
										assign node3292 = (inp[6]) ? node3300 : node3293;
											assign node3293 = (inp[10]) ? node3295 : 16'b0000000111111111;
												assign node3295 = (inp[13]) ? node3297 : 16'b0000000011111111;
													assign node3297 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3300 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3303 = (inp[2]) ? node3309 : node3304;
										assign node3304 = (inp[10]) ? 16'b0000000001111111 : node3305;
											assign node3305 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node3309 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3312 = (inp[6]) ? node3336 : node3313;
									assign node3313 = (inp[0]) ? node3321 : node3314;
										assign node3314 = (inp[13]) ? node3316 : 16'b0000001111111111;
											assign node3316 = (inp[5]) ? node3318 : 16'b0000000001111111;
												assign node3318 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3321 = (inp[5]) ? node3327 : node3322;
											assign node3322 = (inp[9]) ? node3324 : 16'b0000000111111111;
												assign node3324 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3327 = (inp[4]) ? node3333 : node3328;
												assign node3328 = (inp[10]) ? 16'b0000000000111111 : node3329;
													assign node3329 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3333 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3336 = (inp[0]) ? node3346 : node3337;
										assign node3337 = (inp[5]) ? node3339 : 16'b0000000000111111;
											assign node3339 = (inp[11]) ? node3341 : 16'b0000000000111111;
												assign node3341 = (inp[9]) ? 16'b0000000000011111 : node3342;
													assign node3342 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3346 = (inp[11]) ? node3348 : 16'b0000000001111111;
											assign node3348 = (inp[2]) ? node3352 : node3349;
												assign node3349 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3352 = (inp[10]) ? node3354 : 16'b0000000000011111;
													assign node3354 = (inp[9]) ? node3358 : node3355;
														assign node3355 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node3358 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node3361 = (inp[0]) ? node3397 : node3362;
								assign node3362 = (inp[13]) ? node3378 : node3363;
									assign node3363 = (inp[11]) ? node3367 : node3364;
										assign node3364 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3367 = (inp[2]) ? node3373 : node3368;
											assign node3368 = (inp[6]) ? 16'b0000000001111111 : node3369;
												assign node3369 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3373 = (inp[7]) ? 16'b0000000000111111 : node3374;
												assign node3374 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3378 = (inp[6]) ? node3386 : node3379;
										assign node3379 = (inp[9]) ? 16'b0000000000011111 : node3380;
											assign node3380 = (inp[10]) ? 16'b0000000001111111 : node3381;
												assign node3381 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000111111111;
										assign node3386 = (inp[10]) ? 16'b0000000000000111 : node3387;
											assign node3387 = (inp[2]) ? node3389 : 16'b0000000000111111;
												assign node3389 = (inp[11]) ? node3393 : node3390;
													assign node3390 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node3393 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node3397 = (inp[11]) ? node3419 : node3398;
									assign node3398 = (inp[7]) ? node3408 : node3399;
										assign node3399 = (inp[5]) ? node3405 : node3400;
											assign node3400 = (inp[4]) ? node3402 : 16'b0000000001111111;
												assign node3402 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node3405 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node3408 = (inp[4]) ? node3416 : node3409;
											assign node3409 = (inp[2]) ? node3411 : 16'b0000000000111111;
												assign node3411 = (inp[13]) ? 16'b0000000000001111 : node3412;
													assign node3412 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3416 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000011111;
									assign node3419 = (inp[4]) ? node3429 : node3420;
										assign node3420 = (inp[9]) ? node3426 : node3421;
											assign node3421 = (inp[7]) ? node3423 : 16'b0000000000111111;
												assign node3423 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3426 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node3429 = (inp[10]) ? node3437 : node3430;
											assign node3430 = (inp[9]) ? node3432 : 16'b0000000000011111;
												assign node3432 = (inp[13]) ? node3434 : 16'b0000000000001111;
													assign node3434 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node3437 = (inp[13]) ? node3439 : 16'b0000000000011111;
												assign node3439 = (inp[2]) ? node3441 : 16'b0000000000001111;
													assign node3441 = (inp[5]) ? node3443 : 16'b0000000000000111;
														assign node3443 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
			assign node3446 = (inp[5]) ? node3982 : node3447;
				assign node3447 = (inp[6]) ? node3701 : node3448;
					assign node3448 = (inp[2]) ? node3570 : node3449;
						assign node3449 = (inp[12]) ? node3517 : node3450;
							assign node3450 = (inp[13]) ? node3486 : node3451;
								assign node3451 = (inp[3]) ? node3467 : node3452;
									assign node3452 = (inp[4]) ? node3460 : node3453;
										assign node3453 = (inp[0]) ? 16'b0000011111111111 : node3454;
											assign node3454 = (inp[14]) ? 16'b0000111111111111 : node3455;
												assign node3455 = (inp[9]) ? 16'b0000111111111111 : 16'b0011111111111111;
										assign node3460 = (inp[14]) ? node3464 : node3461;
											assign node3461 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3464 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node3467 = (inp[0]) ? node3475 : node3468;
										assign node3468 = (inp[15]) ? node3472 : node3469;
											assign node3469 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3472 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3475 = (inp[7]) ? node3481 : node3476;
											assign node3476 = (inp[9]) ? 16'b0000000011111111 : node3477;
												assign node3477 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node3481 = (inp[15]) ? 16'b0000000111111111 : node3482;
												assign node3482 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node3486 = (inp[0]) ? node3506 : node3487;
									assign node3487 = (inp[7]) ? node3499 : node3488;
										assign node3488 = (inp[15]) ? node3494 : node3489;
											assign node3489 = (inp[3]) ? 16'b0000001111111111 : node3490;
												assign node3490 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3494 = (inp[3]) ? 16'b0000000111111111 : node3495;
												assign node3495 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3499 = (inp[4]) ? 16'b0000000011111111 : node3500;
											assign node3500 = (inp[14]) ? node3502 : 16'b0000000111111111;
												assign node3502 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node3506 = (inp[3]) ? node3512 : node3507;
										assign node3507 = (inp[7]) ? node3509 : 16'b0000000111111111;
											assign node3509 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node3512 = (inp[9]) ? node3514 : 16'b0000000000111111;
											assign node3514 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node3517 = (inp[3]) ? node3545 : node3518;
								assign node3518 = (inp[9]) ? node3532 : node3519;
									assign node3519 = (inp[10]) ? node3523 : node3520;
										assign node3520 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node3523 = (inp[4]) ? 16'b0000000011111111 : node3524;
											assign node3524 = (inp[0]) ? node3526 : 16'b0000001111111111;
												assign node3526 = (inp[14]) ? 16'b0000000111111111 : node3527;
													assign node3527 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3532 = (inp[4]) ? node3536 : node3533;
										assign node3533 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3536 = (inp[14]) ? 16'b0000000001111111 : node3537;
											assign node3537 = (inp[0]) ? 16'b0000000011111111 : node3538;
												assign node3538 = (inp[15]) ? node3540 : 16'b0000000111111111;
													assign node3540 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node3545 = (inp[0]) ? node3557 : node3546;
									assign node3546 = (inp[14]) ? node3550 : node3547;
										assign node3547 = (inp[4]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node3550 = (inp[9]) ? 16'b0000000001111111 : node3551;
											assign node3551 = (inp[13]) ? node3553 : 16'b0000000011111111;
												assign node3553 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node3557 = (inp[10]) ? node3565 : node3558;
										assign node3558 = (inp[15]) ? node3560 : 16'b0000000111111111;
											assign node3560 = (inp[9]) ? 16'b0000000001111111 : node3561;
												assign node3561 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node3565 = (inp[13]) ? node3567 : 16'b0000000000111111;
											assign node3567 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
						assign node3570 = (inp[13]) ? node3634 : node3571;
							assign node3571 = (inp[0]) ? node3601 : node3572;
								assign node3572 = (inp[14]) ? node3586 : node3573;
									assign node3573 = (inp[10]) ? node3583 : node3574;
										assign node3574 = (inp[9]) ? node3578 : node3575;
											assign node3575 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3578 = (inp[4]) ? 16'b0000000111111111 : node3579;
												assign node3579 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3583 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
									assign node3586 = (inp[10]) ? node3596 : node3587;
										assign node3587 = (inp[4]) ? node3593 : node3588;
											assign node3588 = (inp[11]) ? node3590 : 16'b0000000111111111;
												assign node3590 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3593 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node3596 = (inp[11]) ? 16'b0000000001111111 : node3597;
											assign node3597 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3601 = (inp[11]) ? node3617 : node3602;
									assign node3602 = (inp[3]) ? node3610 : node3603;
										assign node3603 = (inp[4]) ? node3605 : 16'b0000111111111111;
											assign node3605 = (inp[12]) ? 16'b0000000111111111 : node3606;
												assign node3606 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node3610 = (inp[9]) ? node3614 : node3611;
											assign node3611 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3614 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3617 = (inp[4]) ? node3631 : node3618;
										assign node3618 = (inp[3]) ? node3624 : node3619;
											assign node3619 = (inp[12]) ? 16'b0000000011111111 : node3620;
												assign node3620 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node3624 = (inp[7]) ? 16'b0000000001111111 : node3625;
												assign node3625 = (inp[9]) ? node3627 : 16'b0000000111111111;
													assign node3627 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3631 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node3634 = (inp[3]) ? node3666 : node3635;
								assign node3635 = (inp[15]) ? node3651 : node3636;
									assign node3636 = (inp[10]) ? node3642 : node3637;
										assign node3637 = (inp[12]) ? node3639 : 16'b0000000111111111;
											assign node3639 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3642 = (inp[9]) ? node3646 : node3643;
											assign node3643 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node3646 = (inp[11]) ? 16'b0000000000111111 : node3647;
												assign node3647 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node3651 = (inp[9]) ? node3661 : node3652;
										assign node3652 = (inp[10]) ? node3656 : node3653;
											assign node3653 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3656 = (inp[14]) ? node3658 : 16'b0000000001111111;
												assign node3658 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node3661 = (inp[12]) ? 16'b0000000000111111 : node3662;
											assign node3662 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3666 = (inp[10]) ? node3682 : node3667;
									assign node3667 = (inp[9]) ? node3673 : node3668;
										assign node3668 = (inp[15]) ? node3670 : 16'b0000000111111111;
											assign node3670 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3673 = (inp[14]) ? node3679 : node3674;
											assign node3674 = (inp[7]) ? node3676 : 16'b0000000011111111;
												assign node3676 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3679 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3682 = (inp[0]) ? node3694 : node3683;
										assign node3683 = (inp[9]) ? node3689 : node3684;
											assign node3684 = (inp[15]) ? node3686 : 16'b0000000011111111;
												assign node3686 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3689 = (inp[11]) ? node3691 : 16'b0000000000111111;
												assign node3691 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3694 = (inp[15]) ? node3696 : 16'b0000000000111111;
											assign node3696 = (inp[4]) ? 16'b0000000000011111 : node3697;
												assign node3697 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node3701 = (inp[15]) ? node3823 : node3702;
						assign node3702 = (inp[7]) ? node3756 : node3703;
							assign node3703 = (inp[10]) ? node3729 : node3704;
								assign node3704 = (inp[14]) ? node3716 : node3705;
									assign node3705 = (inp[9]) ? 16'b0000000011111111 : node3706;
										assign node3706 = (inp[13]) ? node3712 : node3707;
											assign node3707 = (inp[2]) ? node3709 : 16'b0000001111111111;
												assign node3709 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3712 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node3716 = (inp[3]) ? node3724 : node3717;
										assign node3717 = (inp[11]) ? 16'b0000000111111111 : node3718;
											assign node3718 = (inp[12]) ? 16'b0000000011111111 : node3719;
												assign node3719 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node3724 = (inp[12]) ? node3726 : 16'b0000000011111111;
											assign node3726 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3729 = (inp[2]) ? node3743 : node3730;
									assign node3730 = (inp[13]) ? node3736 : node3731;
										assign node3731 = (inp[0]) ? 16'b0000000111111111 : node3732;
											assign node3732 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node3736 = (inp[11]) ? 16'b0000000001111111 : node3737;
											assign node3737 = (inp[14]) ? 16'b0000000111111111 : node3738;
												assign node3738 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3743 = (inp[9]) ? node3751 : node3744;
										assign node3744 = (inp[3]) ? 16'b0000000001111111 : node3745;
											assign node3745 = (inp[14]) ? node3747 : 16'b0000000111111111;
												assign node3747 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3751 = (inp[0]) ? 16'b0000000000111111 : node3752;
											assign node3752 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node3756 = (inp[11]) ? node3774 : node3757;
								assign node3757 = (inp[2]) ? node3769 : node3758;
									assign node3758 = (inp[4]) ? node3764 : node3759;
										assign node3759 = (inp[14]) ? node3761 : 16'b0000000111111111;
											assign node3761 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3764 = (inp[14]) ? node3766 : 16'b0000000011111111;
											assign node3766 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3769 = (inp[0]) ? 16'b0000000000111111 : node3770;
										assign node3770 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node3774 = (inp[14]) ? node3794 : node3775;
									assign node3775 = (inp[13]) ? node3781 : node3776;
										assign node3776 = (inp[3]) ? 16'b0000000011111111 : node3777;
											assign node3777 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3781 = (inp[12]) ? node3787 : node3782;
											assign node3782 = (inp[2]) ? 16'b0000000001111111 : node3783;
												assign node3783 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3787 = (inp[10]) ? 16'b0000000000111111 : node3788;
												assign node3788 = (inp[2]) ? node3790 : 16'b0000000001111111;
													assign node3790 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3794 = (inp[13]) ? node3810 : node3795;
										assign node3795 = (inp[2]) ? node3803 : node3796;
											assign node3796 = (inp[10]) ? 16'b0000000001111111 : node3797;
												assign node3797 = (inp[3]) ? node3799 : 16'b0000000011111111;
													assign node3799 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3803 = (inp[4]) ? node3807 : node3804;
												assign node3804 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node3807 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3810 = (inp[0]) ? node3816 : node3811;
											assign node3811 = (inp[3]) ? node3813 : 16'b0000000000111111;
												assign node3813 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3816 = (inp[2]) ? node3818 : 16'b0000000000011111;
												assign node3818 = (inp[9]) ? node3820 : 16'b0000000000011111;
													assign node3820 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000000111;
						assign node3823 = (inp[12]) ? node3911 : node3824;
							assign node3824 = (inp[9]) ? node3870 : node3825;
								assign node3825 = (inp[0]) ? node3851 : node3826;
									assign node3826 = (inp[2]) ? node3840 : node3827;
										assign node3827 = (inp[10]) ? node3835 : node3828;
											assign node3828 = (inp[14]) ? node3830 : 16'b0000001111111111;
												assign node3830 = (inp[4]) ? 16'b0000000011111111 : node3831;
													assign node3831 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node3835 = (inp[11]) ? 16'b0000000011111111 : node3836;
												assign node3836 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3840 = (inp[14]) ? node3844 : node3841;
											assign node3841 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3844 = (inp[7]) ? 16'b0000000000111111 : node3845;
												assign node3845 = (inp[4]) ? 16'b0000000011111111 : node3846;
													assign node3846 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3851 = (inp[13]) ? node3863 : node3852;
										assign node3852 = (inp[7]) ? node3856 : node3853;
											assign node3853 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node3856 = (inp[3]) ? 16'b0000000001111111 : node3857;
												assign node3857 = (inp[11]) ? 16'b0000000001111111 : node3858;
													assign node3858 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3863 = (inp[11]) ? node3867 : node3864;
											assign node3864 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node3867 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
								assign node3870 = (inp[3]) ? node3880 : node3871;
									assign node3871 = (inp[0]) ? node3877 : node3872;
										assign node3872 = (inp[14]) ? 16'b0000000001111111 : node3873;
											assign node3873 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3877 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3880 = (inp[13]) ? node3898 : node3881;
										assign node3881 = (inp[7]) ? node3887 : node3882;
											assign node3882 = (inp[0]) ? node3884 : 16'b0000000001111111;
												assign node3884 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3887 = (inp[11]) ? node3891 : node3888;
												assign node3888 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3891 = (inp[2]) ? node3893 : 16'b0000000000111111;
													assign node3893 = (inp[4]) ? 16'b0000000000011111 : node3894;
														assign node3894 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3898 = (inp[2]) ? node3904 : node3899;
											assign node3899 = (inp[10]) ? 16'b0000000000011111 : node3900;
												assign node3900 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node3904 = (inp[0]) ? node3908 : node3905;
												assign node3905 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3908 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node3911 = (inp[14]) ? node3947 : node3912;
								assign node3912 = (inp[4]) ? node3932 : node3913;
									assign node3913 = (inp[3]) ? node3921 : node3914;
										assign node3914 = (inp[9]) ? node3916 : 16'b0000000011111111;
											assign node3916 = (inp[2]) ? 16'b0000000000111111 : node3917;
												assign node3917 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node3921 = (inp[13]) ? node3923 : 16'b0000000001111111;
											assign node3923 = (inp[9]) ? node3925 : 16'b0000000000111111;
												assign node3925 = (inp[11]) ? node3927 : 16'b0000000000111111;
													assign node3927 = (inp[7]) ? node3929 : 16'b0000000000011111;
														assign node3929 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3932 = (inp[13]) ? node3938 : node3933;
										assign node3933 = (inp[11]) ? 16'b0000000000111111 : node3934;
											assign node3934 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3938 = (inp[3]) ? node3940 : 16'b0000000000001111;
											assign node3940 = (inp[9]) ? node3944 : node3941;
												assign node3941 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3944 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node3947 = (inp[10]) ? node3959 : node3948;
									assign node3948 = (inp[3]) ? node3954 : node3949;
										assign node3949 = (inp[9]) ? node3951 : 16'b0000000001111111;
											assign node3951 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3954 = (inp[13]) ? node3956 : 16'b0000000000111111;
											assign node3956 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000001111;
									assign node3959 = (inp[7]) ? node3967 : node3960;
										assign node3960 = (inp[9]) ? node3962 : 16'b0000000000111111;
											assign node3962 = (inp[11]) ? node3964 : 16'b0000000000001111;
												assign node3964 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3967 = (inp[4]) ? node3975 : node3968;
											assign node3968 = (inp[2]) ? node3970 : 16'b0000000000111111;
												assign node3970 = (inp[0]) ? 16'b0000000000001111 : node3971;
													assign node3971 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node3975 = (inp[0]) ? node3979 : node3976;
												assign node3976 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node3979 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node3982 = (inp[10]) ? node4250 : node3983;
					assign node3983 = (inp[11]) ? node4111 : node3984;
						assign node3984 = (inp[12]) ? node4050 : node3985;
							assign node3985 = (inp[4]) ? node4021 : node3986;
								assign node3986 = (inp[15]) ? node4006 : node3987;
									assign node3987 = (inp[14]) ? node3995 : node3988;
										assign node3988 = (inp[2]) ? node3990 : 16'b0000011111111111;
											assign node3990 = (inp[6]) ? 16'b0000000111111111 : node3991;
												assign node3991 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node3995 = (inp[2]) ? node4001 : node3996;
											assign node3996 = (inp[7]) ? node3998 : 16'b0000000111111111;
												assign node3998 = (inp[0]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node4001 = (inp[6]) ? node4003 : 16'b0000000011111111;
												assign node4003 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4006 = (inp[3]) ? node4014 : node4007;
										assign node4007 = (inp[13]) ? node4009 : 16'b0000000111111111;
											assign node4009 = (inp[0]) ? 16'b0000000011111111 : node4010;
												assign node4010 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4014 = (inp[7]) ? node4018 : node4015;
											assign node4015 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4018 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node4021 = (inp[13]) ? node4035 : node4022;
									assign node4022 = (inp[2]) ? node4028 : node4023;
										assign node4023 = (inp[6]) ? 16'b0000000001111111 : node4024;
											assign node4024 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4028 = (inp[15]) ? 16'b0000000001111111 : node4029;
											assign node4029 = (inp[14]) ? node4031 : 16'b0000000011111111;
												assign node4031 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node4035 = (inp[15]) ? node4043 : node4036;
										assign node4036 = (inp[3]) ? node4038 : 16'b0000000011111111;
											assign node4038 = (inp[9]) ? 16'b0000000001111111 : node4039;
												assign node4039 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4043 = (inp[2]) ? 16'b0000000001111111 : node4044;
											assign node4044 = (inp[14]) ? node4046 : 16'b0000000000111111;
												assign node4046 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
							assign node4050 = (inp[0]) ? node4072 : node4051;
								assign node4051 = (inp[15]) ? node4061 : node4052;
									assign node4052 = (inp[7]) ? 16'b0000000011111111 : node4053;
										assign node4053 = (inp[3]) ? node4057 : node4054;
											assign node4054 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4057 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node4061 = (inp[9]) ? node4069 : node4062;
										assign node4062 = (inp[3]) ? 16'b0000000000111111 : node4063;
											assign node4063 = (inp[4]) ? 16'b0000000011111111 : node4064;
												assign node4064 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node4069 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4072 = (inp[4]) ? node4088 : node4073;
									assign node4073 = (inp[13]) ? node4079 : node4074;
										assign node4074 = (inp[2]) ? 16'b0000000001111111 : node4075;
											assign node4075 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4079 = (inp[3]) ? node4083 : node4080;
											assign node4080 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node4083 = (inp[9]) ? node4085 : 16'b0000000000111111;
												assign node4085 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4088 = (inp[6]) ? node4102 : node4089;
										assign node4089 = (inp[14]) ? node4091 : 16'b0000000001111111;
											assign node4091 = (inp[9]) ? node4095 : node4092;
												assign node4092 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node4095 = (inp[3]) ? 16'b0000000000011111 : node4096;
													assign node4096 = (inp[2]) ? node4098 : 16'b0000000000111111;
														assign node4098 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4102 = (inp[15]) ? node4108 : node4103;
											assign node4103 = (inp[14]) ? 16'b0000000001111111 : node4104;
												assign node4104 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4108 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node4111 = (inp[13]) ? node4183 : node4112;
							assign node4112 = (inp[0]) ? node4146 : node4113;
								assign node4113 = (inp[14]) ? node4131 : node4114;
									assign node4114 = (inp[9]) ? node4124 : node4115;
										assign node4115 = (inp[15]) ? node4121 : node4116;
											assign node4116 = (inp[7]) ? 16'b0000000011111111 : node4117;
												assign node4117 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4121 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4124 = (inp[4]) ? node4126 : 16'b0000000011111111;
											assign node4126 = (inp[12]) ? 16'b0000000001111111 : node4127;
												assign node4127 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4131 = (inp[3]) ? node4141 : node4132;
										assign node4132 = (inp[4]) ? 16'b0000000001111111 : node4133;
											assign node4133 = (inp[9]) ? node4137 : node4134;
												assign node4134 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4137 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4141 = (inp[2]) ? node4143 : 16'b0000000001111111;
											assign node4143 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node4146 = (inp[3]) ? node4164 : node4147;
									assign node4147 = (inp[2]) ? node4159 : node4148;
										assign node4148 = (inp[9]) ? node4152 : node4149;
											assign node4149 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4152 = (inp[15]) ? node4154 : 16'b0000000001111111;
												assign node4154 = (inp[14]) ? 16'b0000000000111111 : node4155;
													assign node4155 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4159 = (inp[4]) ? 16'b0000000000011111 : node4160;
											assign node4160 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4164 = (inp[9]) ? node4176 : node4165;
										assign node4165 = (inp[2]) ? node4173 : node4166;
											assign node4166 = (inp[4]) ? 16'b0000000000111111 : node4167;
												assign node4167 = (inp[6]) ? 16'b0000000001111111 : node4168;
													assign node4168 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4173 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node4176 = (inp[7]) ? node4180 : node4177;
											assign node4177 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4180 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node4183 = (inp[7]) ? node4209 : node4184;
								assign node4184 = (inp[3]) ? node4194 : node4185;
									assign node4185 = (inp[2]) ? node4191 : node4186;
										assign node4186 = (inp[6]) ? node4188 : 16'b0000000001111111;
											assign node4188 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4191 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4194 = (inp[14]) ? node4196 : 16'b0000000000111111;
										assign node4196 = (inp[12]) ? node4204 : node4197;
											assign node4197 = (inp[15]) ? node4201 : node4198;
												assign node4198 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node4201 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4204 = (inp[6]) ? 16'b0000000000001111 : node4205;
												assign node4205 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node4209 = (inp[14]) ? node4219 : node4210;
									assign node4210 = (inp[2]) ? node4214 : node4211;
										assign node4211 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4214 = (inp[6]) ? 16'b0000000000011111 : node4215;
											assign node4215 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4219 = (inp[0]) ? node4229 : node4220;
										assign node4220 = (inp[3]) ? node4226 : node4221;
											assign node4221 = (inp[9]) ? node4223 : 16'b0000000000111111;
												assign node4223 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4226 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node4229 = (inp[4]) ? node4239 : node4230;
											assign node4230 = (inp[3]) ? node4232 : 16'b0000000000011111;
												assign node4232 = (inp[6]) ? 16'b0000000000001111 : node4233;
													assign node4233 = (inp[2]) ? node4235 : 16'b0000000000011111;
														assign node4235 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4239 = (inp[9]) ? node4243 : node4240;
												assign node4240 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4243 = (inp[6]) ? 16'b0000000000000011 : node4244;
													assign node4244 = (inp[2]) ? node4246 : 16'b0000000000001111;
														assign node4246 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000000111;
					assign node4250 = (inp[9]) ? node4372 : node4251;
						assign node4251 = (inp[14]) ? node4311 : node4252;
							assign node4252 = (inp[2]) ? node4282 : node4253;
								assign node4253 = (inp[4]) ? node4271 : node4254;
									assign node4254 = (inp[11]) ? node4264 : node4255;
										assign node4255 = (inp[0]) ? 16'b0000000011111111 : node4256;
											assign node4256 = (inp[3]) ? node4260 : node4257;
												assign node4257 = (inp[13]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node4260 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4264 = (inp[13]) ? node4266 : 16'b0000000111111111;
											assign node4266 = (inp[6]) ? node4268 : 16'b0000000001111111;
												assign node4268 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node4271 = (inp[13]) ? node4277 : node4272;
										assign node4272 = (inp[7]) ? 16'b0000000001111111 : node4273;
											assign node4273 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4277 = (inp[15]) ? node4279 : 16'b0000000111111111;
											assign node4279 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000011111;
								assign node4282 = (inp[13]) ? node4300 : node4283;
									assign node4283 = (inp[4]) ? node4293 : node4284;
										assign node4284 = (inp[12]) ? node4288 : node4285;
											assign node4285 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4288 = (inp[6]) ? node4290 : 16'b0000000001111111;
												assign node4290 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node4293 = (inp[12]) ? node4297 : node4294;
											assign node4294 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node4297 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node4300 = (inp[15]) ? node4306 : node4301;
										assign node4301 = (inp[7]) ? node4303 : 16'b0000000001111111;
											assign node4303 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node4306 = (inp[3]) ? 16'b0000000000001111 : node4307;
											assign node4307 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node4311 = (inp[15]) ? node4341 : node4312;
								assign node4312 = (inp[7]) ? node4330 : node4313;
									assign node4313 = (inp[2]) ? node4323 : node4314;
										assign node4314 = (inp[4]) ? node4320 : node4315;
											assign node4315 = (inp[13]) ? node4317 : 16'b0000011111111111;
												assign node4317 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4320 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4323 = (inp[13]) ? node4325 : 16'b0000000001111111;
											assign node4325 = (inp[3]) ? 16'b0000000000111111 : node4326;
												assign node4326 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node4330 = (inp[0]) ? node4338 : node4331;
										assign node4331 = (inp[2]) ? 16'b0000000000111111 : node4332;
											assign node4332 = (inp[12]) ? node4334 : 16'b0000000001111111;
												assign node4334 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node4338 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node4341 = (inp[6]) ? node4351 : node4342;
									assign node4342 = (inp[4]) ? node4346 : node4343;
										assign node4343 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4346 = (inp[13]) ? node4348 : 16'b0000000000111111;
											assign node4348 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node4351 = (inp[11]) ? node4363 : node4352;
										assign node4352 = (inp[4]) ? node4356 : node4353;
											assign node4353 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4356 = (inp[3]) ? 16'b0000000000011111 : node4357;
												assign node4357 = (inp[12]) ? node4359 : 16'b0000000000011111;
													assign node4359 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node4363 = (inp[0]) ? node4365 : 16'b0000000000011111;
											assign node4365 = (inp[12]) ? node4369 : node4366;
												assign node4366 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node4369 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node4372 = (inp[4]) ? node4414 : node4373;
							assign node4373 = (inp[2]) ? node4389 : node4374;
								assign node4374 = (inp[11]) ? node4378 : node4375;
									assign node4375 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node4378 = (inp[13]) ? node4386 : node4379;
										assign node4379 = (inp[12]) ? node4383 : node4380;
											assign node4380 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4383 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node4386 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000001111;
								assign node4389 = (inp[6]) ? node4397 : node4390;
									assign node4390 = (inp[7]) ? node4392 : 16'b0000000001111111;
										assign node4392 = (inp[12]) ? 16'b0000000000011111 : node4393;
											assign node4393 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4397 = (inp[13]) ? node4405 : node4398;
										assign node4398 = (inp[3]) ? node4402 : node4399;
											assign node4399 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4402 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4405 = (inp[3]) ? node4407 : 16'b0000000000011111;
											assign node4407 = (inp[15]) ? node4409 : 16'b0000000000011111;
												assign node4409 = (inp[0]) ? 16'b0000000000001111 : node4410;
													assign node4410 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node4414 = (inp[13]) ? node4438 : node4415;
								assign node4415 = (inp[12]) ? node4425 : node4416;
									assign node4416 = (inp[6]) ? node4420 : node4417;
										assign node4417 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4420 = (inp[3]) ? node4422 : 16'b0000000000111111;
											assign node4422 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node4425 = (inp[14]) ? node4427 : 16'b0000000000011111;
										assign node4427 = (inp[15]) ? node4435 : node4428;
											assign node4428 = (inp[6]) ? 16'b0000000000001111 : node4429;
												assign node4429 = (inp[7]) ? node4431 : 16'b0000000000011111;
													assign node4431 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4435 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node4438 = (inp[6]) ? node4450 : node4439;
									assign node4439 = (inp[2]) ? node4447 : node4440;
										assign node4440 = (inp[15]) ? node4442 : 16'b0000000000011111;
											assign node4442 = (inp[3]) ? 16'b0000000000001111 : node4443;
												assign node4443 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node4447 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node4450 = (inp[12]) ? node4460 : node4451;
										assign node4451 = (inp[14]) ? node4455 : node4452;
											assign node4452 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4455 = (inp[2]) ? 16'b0000000000000111 : node4456;
												assign node4456 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node4460 = (inp[15]) ? node4462 : 16'b0000000000001111;
											assign node4462 = (inp[3]) ? 16'b0000000000000001 : 16'b0000000000000011;

endmodule