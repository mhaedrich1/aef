module dtc_split66_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node302;

	assign outp = (inp[3]) ? node230 : node1;
		assign node1 = (inp[9]) ? node107 : node2;
			assign node2 = (inp[4]) ? node74 : node3;
				assign node3 = (inp[0]) ? node23 : node4;
					assign node4 = (inp[6]) ? node10 : node5;
						assign node5 = (inp[1]) ? 3'b001 : node6;
							assign node6 = (inp[5]) ? 3'b000 : 3'b001;
						assign node10 = (inp[11]) ? node12 : 3'b000;
							assign node12 = (inp[2]) ? node14 : 3'b000;
								assign node14 = (inp[10]) ? node16 : 3'b000;
									assign node16 = (inp[8]) ? node18 : 3'b000;
										assign node18 = (inp[7]) ? node20 : 3'b000;
											assign node20 = (inp[5]) ? 3'b000 : 3'b001;
					assign node23 = (inp[6]) ? 3'b001 : node24;
						assign node24 = (inp[5]) ? node50 : node25;
							assign node25 = (inp[1]) ? 3'b000 : node26;
								assign node26 = (inp[7]) ? node40 : node27;
									assign node27 = (inp[10]) ? node33 : node28;
										assign node28 = (inp[8]) ? node30 : 3'b001;
											assign node30 = (inp[2]) ? 3'b001 : 3'b000;
										assign node33 = (inp[2]) ? node37 : node34;
											assign node34 = (inp[8]) ? 3'b000 : 3'b001;
											assign node37 = (inp[8]) ? 3'b000 : 3'b000;
									assign node40 = (inp[2]) ? node46 : node41;
										assign node41 = (inp[8]) ? 3'b000 : node42;
											assign node42 = (inp[10]) ? 3'b001 : 3'b000;
										assign node46 = (inp[8]) ? 3'b001 : 3'b000;
							assign node50 = (inp[1]) ? 3'b001 : node51;
								assign node51 = (inp[7]) ? node61 : node52;
									assign node52 = (inp[10]) ? node54 : 3'b000;
										assign node54 = (inp[2]) ? node58 : node55;
											assign node55 = (inp[8]) ? 3'b000 : 3'b000;
											assign node58 = (inp[8]) ? 3'b001 : 3'b000;
									assign node61 = (inp[10]) ? node67 : node62;
										assign node62 = (inp[2]) ? node64 : 3'b001;
											assign node64 = (inp[8]) ? 3'b001 : 3'b000;
										assign node67 = (inp[2]) ? 3'b000 : node68;
											assign node68 = (inp[11]) ? 3'b000 : 3'b000;
				assign node74 = (inp[0]) ? node76 : 3'b000;
					assign node76 = (inp[10]) ? node88 : node77;
						assign node77 = (inp[6]) ? node83 : node78;
							assign node78 = (inp[5]) ? 3'b000 : node79;
								assign node79 = (inp[1]) ? 3'b001 : 3'b000;
							assign node83 = (inp[1]) ? 3'b000 : node84;
								assign node84 = (inp[5]) ? 3'b001 : 3'b000;
						assign node88 = (inp[6]) ? node102 : node89;
							assign node89 = (inp[5]) ? node97 : node90;
								assign node90 = (inp[1]) ? 3'b001 : node91;
									assign node91 = (inp[2]) ? node93 : 3'b000;
										assign node93 = (inp[7]) ? 3'b001 : 3'b000;
								assign node97 = (inp[1]) ? 3'b000 : node98;
									assign node98 = (inp[7]) ? 3'b001 : 3'b000;
							assign node102 = (inp[5]) ? node104 : 3'b000;
								assign node104 = (inp[1]) ? 3'b000 : 3'b001;
			assign node107 = (inp[6]) ? node183 : node108;
				assign node108 = (inp[4]) ? node154 : node109;
					assign node109 = (inp[0]) ? node119 : node110;
						assign node110 = (inp[1]) ? node116 : node111;
							assign node111 = (inp[5]) ? 3'b100 : node112;
								assign node112 = (inp[7]) ? 3'b110 : 3'b010;
							assign node116 = (inp[5]) ? 3'b010 : 3'b110;
						assign node119 = (inp[5]) ? node141 : node120;
							assign node120 = (inp[7]) ? node130 : node121;
								assign node121 = (inp[1]) ? 3'b001 : node122;
									assign node122 = (inp[8]) ? 3'b001 : node123;
										assign node123 = (inp[11]) ? node125 : 3'b001;
											assign node125 = (inp[2]) ? 3'b001 : 3'b110;
								assign node130 = (inp[1]) ? 3'b101 : node131;
									assign node131 = (inp[2]) ? node137 : node132;
										assign node132 = (inp[11]) ? node134 : 3'b001;
											assign node134 = (inp[8]) ? 3'b001 : 3'b110;
										assign node137 = (inp[11]) ? 3'b001 : 3'b110;
							assign node141 = (inp[1]) ? 3'b110 : node142;
								assign node142 = (inp[11]) ? node148 : node143;
									assign node143 = (inp[8]) ? node145 : 3'b001;
										assign node145 = (inp[2]) ? 3'b110 : 3'b001;
									assign node148 = (inp[8]) ? 3'b001 : node149;
										assign node149 = (inp[2]) ? 3'b001 : 3'b110;
					assign node154 = (inp[0]) ? node166 : node155;
						assign node155 = (inp[7]) ? 3'b000 : node156;
							assign node156 = (inp[5]) ? 3'b000 : node157;
								assign node157 = (inp[2]) ? node159 : 3'b000;
									assign node159 = (inp[11]) ? 3'b000 : node160;
										assign node160 = (inp[1]) ? 3'b100 : 3'b000;
						assign node166 = (inp[5]) ? node176 : node167;
							assign node167 = (inp[1]) ? 3'b010 : node168;
								assign node168 = (inp[7]) ? node170 : 3'b100;
									assign node170 = (inp[2]) ? node172 : 3'b100;
										assign node172 = (inp[10]) ? 3'b010 : 3'b100;
							assign node176 = (inp[1]) ? 3'b100 : node177;
								assign node177 = (inp[10]) ? node179 : 3'b100;
									assign node179 = (inp[7]) ? 3'b010 : 3'b100;
				assign node183 = (inp[0]) ? node199 : node184;
					assign node184 = (inp[4]) ? 3'b001 : node185;
						assign node185 = (inp[11]) ? node187 : 3'b001;
							assign node187 = (inp[2]) ? node189 : 3'b001;
								assign node189 = (inp[8]) ? node191 : 3'b001;
									assign node191 = (inp[7]) ? node193 : 3'b001;
										assign node193 = (inp[10]) ? node195 : 3'b001;
											assign node195 = (inp[5]) ? 3'b001 : 3'b011;
					assign node199 = (inp[4]) ? node213 : node200;
						assign node200 = (inp[1]) ? node210 : node201;
							assign node201 = (inp[7]) ? node203 : 3'b011;
								assign node203 = (inp[10]) ? node205 : 3'b011;
									assign node205 = (inp[5]) ? 3'b111 : node206;
										assign node206 = (inp[2]) ? 3'b111 : 3'b011;
							assign node210 = (inp[5]) ? 3'b011 : 3'b111;
						assign node213 = (inp[5]) ? node223 : node214;
							assign node214 = (inp[1]) ? 3'b101 : node215;
								assign node215 = (inp[2]) ? node217 : 3'b001;
									assign node217 = (inp[7]) ? node219 : 3'b001;
										assign node219 = (inp[10]) ? 3'b101 : 3'b001;
							assign node223 = (inp[1]) ? 3'b001 : node224;
								assign node224 = (inp[7]) ? node226 : 3'b010;
									assign node226 = (inp[10]) ? 3'b110 : 3'b010;
		assign node230 = (inp[6]) ? node232 : 3'b000;
			assign node232 = (inp[0]) ? node248 : node233;
				assign node233 = (inp[4]) ? node237 : node234;
					assign node234 = (inp[9]) ? 3'b100 : 3'b000;
					assign node237 = (inp[9]) ? 3'b000 : node238;
						assign node238 = (inp[1]) ? node240 : 3'b010;
							assign node240 = (inp[10]) ? node242 : 3'b010;
								assign node242 = (inp[2]) ? 3'b100 : node243;
									assign node243 = (inp[5]) ? 3'b100 : 3'b010;
				assign node248 = (inp[4]) ? node252 : node249;
					assign node249 = (inp[9]) ? 3'b010 : 3'b001;
					assign node252 = (inp[9]) ? node288 : node253;
						assign node253 = (inp[1]) ? node263 : node254;
							assign node254 = (inp[7]) ? node256 : 3'b010;
								assign node256 = (inp[10]) ? 3'b010 : node257;
									assign node257 = (inp[2]) ? 3'b110 : node258;
										assign node258 = (inp[11]) ? 3'b010 : 3'b110;
							assign node263 = (inp[7]) ? node265 : 3'b110;
								assign node265 = (inp[10]) ? node277 : node266;
									assign node266 = (inp[2]) ? node272 : node267;
										assign node267 = (inp[11]) ? node269 : 3'b110;
											assign node269 = (inp[8]) ? 3'b110 : 3'b010;
										assign node272 = (inp[8]) ? node274 : 3'b110;
											assign node274 = (inp[11]) ? 3'b110 : 3'b001;
									assign node277 = (inp[8]) ? node283 : node278;
										assign node278 = (inp[2]) ? 3'b010 : node279;
											assign node279 = (inp[11]) ? 3'b110 : 3'b010;
										assign node283 = (inp[2]) ? node285 : 3'b010;
											assign node285 = (inp[11]) ? 3'b010 : 3'b110;
						assign node288 = (inp[10]) ? 3'b000 : node289;
							assign node289 = (inp[7]) ? node291 : 3'b000;
								assign node291 = (inp[11]) ? node299 : node292;
									assign node292 = (inp[1]) ? node294 : 3'b100;
										assign node294 = (inp[2]) ? node296 : 3'b100;
											assign node296 = (inp[8]) ? 3'b010 : 3'b100;
									assign node299 = (inp[1]) ? node301 : 3'b000;
										assign node301 = (inp[8]) ? 3'b100 : node302;
											assign node302 = (inp[2]) ? 3'b100 : 3'b000;

endmodule