module dtc_split66_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node946;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1093;
	wire [3-1:0] node1097;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1136;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1156;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1251;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1356;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1383;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1389;
	wire [3-1:0] node1391;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1413;
	wire [3-1:0] node1414;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1443;
	wire [3-1:0] node1445;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1454;
	wire [3-1:0] node1457;
	wire [3-1:0] node1459;
	wire [3-1:0] node1462;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1481;
	wire [3-1:0] node1482;
	wire [3-1:0] node1485;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1493;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1515;
	wire [3-1:0] node1516;
	wire [3-1:0] node1517;
	wire [3-1:0] node1520;
	wire [3-1:0] node1523;
	wire [3-1:0] node1525;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1559;
	wire [3-1:0] node1562;
	wire [3-1:0] node1563;
	wire [3-1:0] node1564;
	wire [3-1:0] node1568;
	wire [3-1:0] node1571;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1575;
	wire [3-1:0] node1576;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1583;
	wire [3-1:0] node1586;
	wire [3-1:0] node1588;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1594;
	wire [3-1:0] node1595;
	wire [3-1:0] node1598;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1605;
	wire [3-1:0] node1608;
	wire [3-1:0] node1609;
	wire [3-1:0] node1610;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1616;
	wire [3-1:0] node1619;
	wire [3-1:0] node1621;
	wire [3-1:0] node1624;
	wire [3-1:0] node1625;
	wire [3-1:0] node1628;
	wire [3-1:0] node1630;
	wire [3-1:0] node1633;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1637;
	wire [3-1:0] node1640;
	wire [3-1:0] node1641;
	wire [3-1:0] node1644;
	wire [3-1:0] node1647;
	wire [3-1:0] node1648;
	wire [3-1:0] node1649;
	wire [3-1:0] node1652;
	wire [3-1:0] node1655;
	wire [3-1:0] node1656;
	wire [3-1:0] node1660;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1666;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1676;
	wire [3-1:0] node1679;
	wire [3-1:0] node1680;
	wire [3-1:0] node1683;
	wire [3-1:0] node1686;
	wire [3-1:0] node1687;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1693;
	wire [3-1:0] node1694;
	wire [3-1:0] node1698;
	wire [3-1:0] node1701;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;
	wire [3-1:0] node1704;
	wire [3-1:0] node1705;
	wire [3-1:0] node1706;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1711;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1719;
	wire [3-1:0] node1720;
	wire [3-1:0] node1721;
	wire [3-1:0] node1724;
	wire [3-1:0] node1727;
	wire [3-1:0] node1729;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1738;
	wire [3-1:0] node1741;
	wire [3-1:0] node1742;
	wire [3-1:0] node1745;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1750;
	wire [3-1:0] node1753;
	wire [3-1:0] node1757;
	wire [3-1:0] node1758;
	wire [3-1:0] node1759;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1766;
	wire [3-1:0] node1767;
	wire [3-1:0] node1768;
	wire [3-1:0] node1772;
	wire [3-1:0] node1773;
	wire [3-1:0] node1776;
	wire [3-1:0] node1779;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1783;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1790;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1795;
	wire [3-1:0] node1799;
	wire [3-1:0] node1800;
	wire [3-1:0] node1804;
	wire [3-1:0] node1805;
	wire [3-1:0] node1806;
	wire [3-1:0] node1807;
	wire [3-1:0] node1809;
	wire [3-1:0] node1812;
	wire [3-1:0] node1813;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1825;
	wire [3-1:0] node1828;
	wire [3-1:0] node1829;
	wire [3-1:0] node1830;
	wire [3-1:0] node1831;
	wire [3-1:0] node1832;
	wire [3-1:0] node1835;
	wire [3-1:0] node1838;
	wire [3-1:0] node1840;
	wire [3-1:0] node1843;
	wire [3-1:0] node1844;
	wire [3-1:0] node1847;
	wire [3-1:0] node1849;
	wire [3-1:0] node1852;
	wire [3-1:0] node1853;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1860;
	wire [3-1:0] node1861;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1864;
	wire [3-1:0] node1866;
	wire [3-1:0] node1869;
	wire [3-1:0] node1871;
	wire [3-1:0] node1874;
	wire [3-1:0] node1875;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1883;
	wire [3-1:0] node1884;
	wire [3-1:0] node1885;
	wire [3-1:0] node1886;
	wire [3-1:0] node1889;
	wire [3-1:0] node1892;
	wire [3-1:0] node1894;
	wire [3-1:0] node1897;
	wire [3-1:0] node1899;
	wire [3-1:0] node1901;
	wire [3-1:0] node1904;
	wire [3-1:0] node1905;
	wire [3-1:0] node1906;
	wire [3-1:0] node1908;
	wire [3-1:0] node1910;
	wire [3-1:0] node1913;
	wire [3-1:0] node1914;
	wire [3-1:0] node1915;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1924;
	wire [3-1:0] node1925;
	wire [3-1:0] node1926;
	wire [3-1:0] node1927;
	wire [3-1:0] node1930;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1937;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1943;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1953;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1959;
	wire [3-1:0] node1960;
	wire [3-1:0] node1965;
	wire [3-1:0] node1966;
	wire [3-1:0] node1967;
	wire [3-1:0] node1968;
	wire [3-1:0] node1972;
	wire [3-1:0] node1973;
	wire [3-1:0] node1978;
	wire [3-1:0] node1979;
	wire [3-1:0] node1980;
	wire [3-1:0] node1981;
	wire [3-1:0] node1982;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1986;
	wire [3-1:0] node1989;
	wire [3-1:0] node1991;
	wire [3-1:0] node1994;
	wire [3-1:0] node1995;
	wire [3-1:0] node1997;
	wire [3-1:0] node2000;
	wire [3-1:0] node2002;
	wire [3-1:0] node2005;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2008;
	wire [3-1:0] node2012;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2018;
	wire [3-1:0] node2019;
	wire [3-1:0] node2022;
	wire [3-1:0] node2025;
	wire [3-1:0] node2026;
	wire [3-1:0] node2027;
	wire [3-1:0] node2029;
	wire [3-1:0] node2032;
	wire [3-1:0] node2034;
	wire [3-1:0] node2037;
	wire [3-1:0] node2038;
	wire [3-1:0] node2041;
	wire [3-1:0] node2044;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2047;
	wire [3-1:0] node2048;
	wire [3-1:0] node2051;
	wire [3-1:0] node2054;
	wire [3-1:0] node2056;
	wire [3-1:0] node2059;
	wire [3-1:0] node2060;
	wire [3-1:0] node2061;
	wire [3-1:0] node2064;
	wire [3-1:0] node2067;
	wire [3-1:0] node2068;
	wire [3-1:0] node2071;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2076;
	wire [3-1:0] node2079;
	wire [3-1:0] node2082;
	wire [3-1:0] node2083;
	wire [3-1:0] node2084;
	wire [3-1:0] node2085;
	wire [3-1:0] node2088;
	wire [3-1:0] node2092;
	wire [3-1:0] node2093;
	wire [3-1:0] node2094;
	wire [3-1:0] node2097;
	wire [3-1:0] node2100;
	wire [3-1:0] node2101;
	wire [3-1:0] node2104;
	wire [3-1:0] node2107;
	wire [3-1:0] node2108;
	wire [3-1:0] node2109;
	wire [3-1:0] node2110;
	wire [3-1:0] node2111;
	wire [3-1:0] node2112;
	wire [3-1:0] node2115;
	wire [3-1:0] node2118;
	wire [3-1:0] node2119;
	wire [3-1:0] node2122;
	wire [3-1:0] node2125;
	wire [3-1:0] node2126;
	wire [3-1:0] node2127;
	wire [3-1:0] node2128;
	wire [3-1:0] node2132;
	wire [3-1:0] node2134;
	wire [3-1:0] node2137;
	wire [3-1:0] node2138;
	wire [3-1:0] node2141;
	wire [3-1:0] node2144;
	wire [3-1:0] node2145;
	wire [3-1:0] node2148;
	wire [3-1:0] node2151;
	wire [3-1:0] node2152;
	wire [3-1:0] node2153;
	wire [3-1:0] node2154;
	wire [3-1:0] node2155;
	wire [3-1:0] node2159;
	wire [3-1:0] node2160;
	wire [3-1:0] node2165;
	wire [3-1:0] node2166;
	wire [3-1:0] node2167;
	wire [3-1:0] node2168;
	wire [3-1:0] node2172;
	wire [3-1:0] node2173;
	wire [3-1:0] node2178;
	wire [3-1:0] node2179;
	wire [3-1:0] node2180;
	wire [3-1:0] node2181;
	wire [3-1:0] node2184;
	wire [3-1:0] node2187;
	wire [3-1:0] node2188;
	wire [3-1:0] node2189;
	wire [3-1:0] node2193;
	wire [3-1:0] node2194;
	wire [3-1:0] node2198;
	wire [3-1:0] node2199;
	wire [3-1:0] node2200;
	wire [3-1:0] node2201;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2210;
	wire [3-1:0] node2211;

	assign outp = (inp[5]) ? node1324 : node1;
		assign node1 = (inp[8]) ? node729 : node2;
			assign node2 = (inp[4]) ? node424 : node3;
				assign node3 = (inp[6]) ? node223 : node4;
					assign node4 = (inp[0]) ? node112 : node5;
						assign node5 = (inp[9]) ? node59 : node6;
							assign node6 = (inp[1]) ? node30 : node7;
								assign node7 = (inp[3]) ? node19 : node8;
									assign node8 = (inp[11]) ? node12 : node9;
										assign node9 = (inp[10]) ? 3'b010 : 3'b000;
										assign node12 = (inp[2]) ? node16 : node13;
											assign node13 = (inp[10]) ? 3'b011 : 3'b000;
											assign node16 = (inp[7]) ? 3'b000 : 3'b011;
									assign node19 = (inp[10]) ? node25 : node20;
										assign node20 = (inp[7]) ? node22 : 3'b010;
											assign node22 = (inp[11]) ? 3'b000 : 3'b011;
										assign node25 = (inp[2]) ? node27 : 3'b001;
											assign node27 = (inp[7]) ? 3'b000 : 3'b000;
								assign node30 = (inp[2]) ? node44 : node31;
									assign node31 = (inp[7]) ? node39 : node32;
										assign node32 = (inp[10]) ? node36 : node33;
											assign node33 = (inp[3]) ? 3'b010 : 3'b000;
											assign node36 = (inp[3]) ? 3'b000 : 3'b010;
										assign node39 = (inp[11]) ? 3'b011 : node40;
											assign node40 = (inp[3]) ? 3'b011 : 3'b000;
									assign node44 = (inp[3]) ? node52 : node45;
										assign node45 = (inp[11]) ? node49 : node46;
											assign node46 = (inp[10]) ? 3'b011 : 3'b001;
											assign node49 = (inp[10]) ? 3'b001 : 3'b011;
										assign node52 = (inp[10]) ? node56 : node53;
											assign node53 = (inp[7]) ? 3'b000 : 3'b011;
											assign node56 = (inp[7]) ? 3'b000 : 3'b000;
							assign node59 = (inp[1]) ? node83 : node60;
								assign node60 = (inp[10]) ? node72 : node61;
									assign node61 = (inp[11]) ? node65 : node62;
										assign node62 = (inp[3]) ? 3'b011 : 3'b001;
										assign node65 = (inp[3]) ? node69 : node66;
											assign node66 = (inp[7]) ? 3'b010 : 3'b001;
											assign node69 = (inp[7]) ? 3'b001 : 3'b011;
									assign node72 = (inp[3]) ? node78 : node73;
										assign node73 = (inp[11]) ? node75 : 3'b011;
											assign node75 = (inp[7]) ? 3'b001 : 3'b010;
										assign node78 = (inp[11]) ? 3'b010 : node79;
											assign node79 = (inp[2]) ? 3'b001 : 3'b000;
								assign node83 = (inp[2]) ? node97 : node84;
									assign node84 = (inp[7]) ? node92 : node85;
										assign node85 = (inp[10]) ? node89 : node86;
											assign node86 = (inp[3]) ? 3'b011 : 3'b001;
											assign node89 = (inp[3]) ? 3'b000 : 3'b010;
										assign node92 = (inp[3]) ? 3'b010 : node93;
											assign node93 = (inp[11]) ? 3'b000 : 3'b001;
									assign node97 = (inp[3]) ? node105 : node98;
										assign node98 = (inp[10]) ? node102 : node99;
											assign node99 = (inp[7]) ? 3'b000 : 3'b000;
											assign node102 = (inp[11]) ? 3'b000 : 3'b010;
										assign node105 = (inp[10]) ? node109 : node106;
											assign node106 = (inp[11]) ? 3'b000 : 3'b010;
											assign node109 = (inp[7]) ? 3'b011 : 3'b000;
						assign node112 = (inp[9]) ? node168 : node113;
							assign node113 = (inp[1]) ? node141 : node114;
								assign node114 = (inp[7]) ? node126 : node115;
									assign node115 = (inp[10]) ? node119 : node116;
										assign node116 = (inp[3]) ? 3'b011 : 3'b001;
										assign node119 = (inp[3]) ? node123 : node120;
											assign node120 = (inp[11]) ? 3'b010 : 3'b011;
											assign node123 = (inp[11]) ? 3'b001 : 3'b000;
									assign node126 = (inp[3]) ? node134 : node127;
										assign node127 = (inp[10]) ? node131 : node128;
											assign node128 = (inp[11]) ? 3'b010 : 3'b001;
											assign node131 = (inp[11]) ? 3'b001 : 3'b011;
										assign node134 = (inp[11]) ? node138 : node135;
											assign node135 = (inp[10]) ? 3'b000 : 3'b010;
											assign node138 = (inp[10]) ? 3'b010 : 3'b001;
								assign node141 = (inp[3]) ? node155 : node142;
									assign node142 = (inp[2]) ? node148 : node143;
										assign node143 = (inp[11]) ? node145 : 3'b001;
											assign node145 = (inp[7]) ? 3'b010 : 3'b001;
										assign node148 = (inp[11]) ? node152 : node149;
											assign node149 = (inp[10]) ? 3'b010 : 3'b000;
											assign node152 = (inp[7]) ? 3'b000 : 3'b000;
									assign node155 = (inp[10]) ? node163 : node156;
										assign node156 = (inp[11]) ? node160 : node157;
											assign node157 = (inp[2]) ? 3'b011 : 3'b010;
											assign node160 = (inp[2]) ? 3'b000 : 3'b001;
										assign node163 = (inp[2]) ? 3'b001 : node164;
											assign node164 = (inp[7]) ? 3'b010 : 3'b000;
							assign node168 = (inp[2]) ? node196 : node169;
								assign node169 = (inp[10]) ? node181 : node170;
									assign node170 = (inp[3]) ? node176 : node171;
										assign node171 = (inp[7]) ? node173 : 3'b000;
											assign node173 = (inp[11]) ? 3'b011 : 3'b000;
										assign node176 = (inp[7]) ? node178 : 3'b010;
											assign node178 = (inp[11]) ? 3'b000 : 3'b011;
									assign node181 = (inp[3]) ? node189 : node182;
										assign node182 = (inp[7]) ? node186 : node183;
											assign node183 = (inp[11]) ? 3'b011 : 3'b010;
											assign node186 = (inp[11]) ? 3'b000 : 3'b010;
										assign node189 = (inp[11]) ? node193 : node190;
											assign node190 = (inp[7]) ? 3'b000 : 3'b000;
											assign node193 = (inp[7]) ? 3'b011 : 3'b000;
								assign node196 = (inp[1]) ? node210 : node197;
									assign node197 = (inp[10]) ? node205 : node198;
										assign node198 = (inp[7]) ? node202 : node199;
											assign node199 = (inp[3]) ? 3'b010 : 3'b000;
											assign node202 = (inp[3]) ? 3'b000 : 3'b011;
										assign node205 = (inp[7]) ? 3'b000 : node206;
											assign node206 = (inp[11]) ? 3'b011 : 3'b001;
									assign node210 = (inp[7]) ? node216 : node211;
										assign node211 = (inp[10]) ? node213 : 3'b011;
											assign node213 = (inp[11]) ? 3'b010 : 3'b011;
										assign node216 = (inp[3]) ? node220 : node217;
											assign node217 = (inp[10]) ? 3'b011 : 3'b001;
											assign node220 = (inp[11]) ? 3'b001 : 3'b000;
					assign node223 = (inp[10]) ? node323 : node224;
						assign node224 = (inp[3]) ? node274 : node225;
							assign node225 = (inp[11]) ? node245 : node226;
								assign node226 = (inp[7]) ? node234 : node227;
									assign node227 = (inp[9]) ? 3'b101 : node228;
										assign node228 = (inp[0]) ? node230 : 3'b100;
											assign node230 = (inp[2]) ? 3'b101 : 3'b100;
									assign node234 = (inp[2]) ? node240 : node235;
										assign node235 = (inp[9]) ? node237 : 3'b111;
											assign node237 = (inp[0]) ? 3'b110 : 3'b111;
										assign node240 = (inp[1]) ? 3'b110 : node241;
											assign node241 = (inp[9]) ? 3'b110 : 3'b110;
								assign node245 = (inp[1]) ? node259 : node246;
									assign node246 = (inp[0]) ? node252 : node247;
										assign node247 = (inp[7]) ? 3'b100 : node248;
											assign node248 = (inp[9]) ? 3'b101 : 3'b100;
										assign node252 = (inp[9]) ? node256 : node253;
											assign node253 = (inp[7]) ? 3'b100 : 3'b101;
											assign node256 = (inp[7]) ? 3'b101 : 3'b100;
									assign node259 = (inp[2]) ? node267 : node260;
										assign node260 = (inp[0]) ? node264 : node261;
											assign node261 = (inp[7]) ? 3'b100 : 3'b100;
											assign node264 = (inp[7]) ? 3'b100 : 3'b101;
										assign node267 = (inp[9]) ? node271 : node268;
											assign node268 = (inp[7]) ? 3'b100 : 3'b100;
											assign node271 = (inp[0]) ? 3'b100 : 3'b100;
							assign node274 = (inp[11]) ? node302 : node275;
								assign node275 = (inp[7]) ? node289 : node276;
									assign node276 = (inp[0]) ? node282 : node277;
										assign node277 = (inp[2]) ? 3'b110 : node278;
											assign node278 = (inp[1]) ? 3'b110 : 3'b111;
										assign node282 = (inp[9]) ? node286 : node283;
											assign node283 = (inp[2]) ? 3'b111 : 3'b110;
											assign node286 = (inp[2]) ? 3'b110 : 3'b111;
									assign node289 = (inp[1]) ? node295 : node290;
										assign node290 = (inp[2]) ? node292 : 3'b100;
											assign node292 = (inp[9]) ? 3'b100 : 3'b100;
										assign node295 = (inp[9]) ? node299 : node296;
											assign node296 = (inp[0]) ? 3'b100 : 3'b101;
											assign node299 = (inp[0]) ? 3'b101 : 3'b100;
								assign node302 = (inp[9]) ? node312 : node303;
									assign node303 = (inp[0]) ? node307 : node304;
										assign node304 = (inp[1]) ? 3'b111 : 3'b110;
										assign node307 = (inp[2]) ? 3'b111 : node308;
											assign node308 = (inp[1]) ? 3'b110 : 3'b111;
									assign node312 = (inp[1]) ? node316 : node313;
										assign node313 = (inp[0]) ? 3'b110 : 3'b111;
										assign node316 = (inp[0]) ? node320 : node317;
											assign node317 = (inp[2]) ? 3'b111 : 3'b110;
											assign node320 = (inp[2]) ? 3'b110 : 3'b111;
						assign node323 = (inp[3]) ? node375 : node324;
							assign node324 = (inp[7]) ? node354 : node325;
								assign node325 = (inp[9]) ? node339 : node326;
									assign node326 = (inp[1]) ? node334 : node327;
										assign node327 = (inp[0]) ? node331 : node328;
											assign node328 = (inp[2]) ? 3'b111 : 3'b110;
											assign node331 = (inp[11]) ? 3'b110 : 3'b110;
										assign node334 = (inp[0]) ? node336 : 3'b110;
											assign node336 = (inp[11]) ? 3'b110 : 3'b111;
									assign node339 = (inp[2]) ? node347 : node340;
										assign node340 = (inp[11]) ? node344 : node341;
											assign node341 = (inp[0]) ? 3'b110 : 3'b111;
											assign node344 = (inp[0]) ? 3'b111 : 3'b110;
										assign node347 = (inp[11]) ? node351 : node348;
											assign node348 = (inp[0]) ? 3'b111 : 3'b110;
											assign node351 = (inp[0]) ? 3'b110 : 3'b110;
								assign node354 = (inp[11]) ? node362 : node355;
									assign node355 = (inp[0]) ? 3'b101 : node356;
										assign node356 = (inp[1]) ? node358 : 3'b100;
											assign node358 = (inp[9]) ? 3'b101 : 3'b100;
									assign node362 = (inp[0]) ? node368 : node363;
										assign node363 = (inp[2]) ? node365 : 3'b110;
											assign node365 = (inp[1]) ? 3'b111 : 3'b110;
										assign node368 = (inp[9]) ? node372 : node369;
											assign node369 = (inp[2]) ? 3'b110 : 3'b111;
											assign node372 = (inp[2]) ? 3'b111 : 3'b110;
							assign node375 = (inp[11]) ? node401 : node376;
								assign node376 = (inp[7]) ? node388 : node377;
									assign node377 = (inp[9]) ? node383 : node378;
										assign node378 = (inp[0]) ? 3'b100 : node379;
											assign node379 = (inp[1]) ? 3'b100 : 3'b101;
										assign node383 = (inp[1]) ? 3'b101 : node384;
											assign node384 = (inp[0]) ? 3'b101 : 3'b100;
									assign node388 = (inp[2]) ? node394 : node389;
										assign node389 = (inp[0]) ? node391 : 3'b111;
											assign node391 = (inp[9]) ? 3'b110 : 3'b110;
										assign node394 = (inp[1]) ? node398 : node395;
											assign node395 = (inp[9]) ? 3'b111 : 3'b110;
											assign node398 = (inp[0]) ? 3'b110 : 3'b110;
								assign node401 = (inp[1]) ? node409 : node402;
									assign node402 = (inp[9]) ? node406 : node403;
										assign node403 = (inp[0]) ? 3'b101 : 3'b100;
										assign node406 = (inp[0]) ? 3'b100 : 3'b101;
									assign node409 = (inp[0]) ? node417 : node410;
										assign node410 = (inp[7]) ? node414 : node411;
											assign node411 = (inp[2]) ? 3'b100 : 3'b100;
											assign node414 = (inp[2]) ? 3'b101 : 3'b100;
										assign node417 = (inp[9]) ? node421 : node418;
											assign node418 = (inp[7]) ? 3'b101 : 3'b100;
											assign node421 = (inp[2]) ? 3'b100 : 3'b101;
				assign node424 = (inp[11]) ? node582 : node425;
					assign node425 = (inp[10]) ? node517 : node426;
						assign node426 = (inp[9]) ? node478 : node427;
							assign node427 = (inp[7]) ? node455 : node428;
								assign node428 = (inp[3]) ? node444 : node429;
									assign node429 = (inp[6]) ? node437 : node430;
										assign node430 = (inp[2]) ? node434 : node431;
											assign node431 = (inp[0]) ? 3'b101 : 3'b100;
											assign node434 = (inp[0]) ? 3'b100 : 3'b101;
										assign node437 = (inp[0]) ? node441 : node438;
											assign node438 = (inp[1]) ? 3'b100 : 3'b100;
											assign node441 = (inp[2]) ? 3'b100 : 3'b100;
									assign node444 = (inp[2]) ? node450 : node445;
										assign node445 = (inp[0]) ? node447 : 3'b100;
											assign node447 = (inp[1]) ? 3'b100 : 3'b101;
										assign node450 = (inp[0]) ? node452 : 3'b101;
											assign node452 = (inp[1]) ? 3'b101 : 3'b100;
								assign node455 = (inp[0]) ? node467 : node456;
									assign node456 = (inp[2]) ? node462 : node457;
										assign node457 = (inp[1]) ? node459 : 3'b100;
											assign node459 = (inp[3]) ? 3'b100 : 3'b100;
										assign node462 = (inp[3]) ? node464 : 3'b101;
											assign node464 = (inp[6]) ? 3'b100 : 3'b100;
									assign node467 = (inp[2]) ? node473 : node468;
										assign node468 = (inp[3]) ? node470 : 3'b101;
											assign node470 = (inp[1]) ? 3'b100 : 3'b101;
										assign node473 = (inp[3]) ? node475 : 3'b100;
											assign node475 = (inp[6]) ? 3'b100 : 3'b100;
							assign node478 = (inp[0]) ? node498 : node479;
								assign node479 = (inp[2]) ? node487 : node480;
									assign node480 = (inp[3]) ? node482 : 3'b100;
										assign node482 = (inp[7]) ? node484 : 3'b100;
											assign node484 = (inp[6]) ? 3'b100 : 3'b101;
									assign node487 = (inp[3]) ? node493 : node488;
										assign node488 = (inp[7]) ? 3'b101 : node489;
											assign node489 = (inp[1]) ? 3'b100 : 3'b101;
										assign node493 = (inp[7]) ? node495 : 3'b101;
											assign node495 = (inp[1]) ? 3'b100 : 3'b100;
								assign node498 = (inp[2]) ? node506 : node499;
									assign node499 = (inp[1]) ? node501 : 3'b101;
										assign node501 = (inp[7]) ? 3'b101 : node502;
											assign node502 = (inp[3]) ? 3'b100 : 3'b100;
									assign node506 = (inp[3]) ? node512 : node507;
										assign node507 = (inp[6]) ? node509 : 3'b100;
											assign node509 = (inp[1]) ? 3'b101 : 3'b100;
										assign node512 = (inp[6]) ? 3'b101 : node513;
											assign node513 = (inp[1]) ? 3'b100 : 3'b100;
						assign node517 = (inp[3]) ? node549 : node518;
							assign node518 = (inp[0]) ? node534 : node519;
								assign node519 = (inp[2]) ? node527 : node520;
									assign node520 = (inp[1]) ? 3'b110 : node521;
										assign node521 = (inp[6]) ? node523 : 3'b110;
											assign node523 = (inp[7]) ? 3'b111 : 3'b110;
									assign node527 = (inp[7]) ? node529 : 3'b111;
										assign node529 = (inp[6]) ? node531 : 3'b111;
											assign node531 = (inp[1]) ? 3'b111 : 3'b110;
								assign node534 = (inp[2]) ? node542 : node535;
									assign node535 = (inp[7]) ? node537 : 3'b111;
										assign node537 = (inp[1]) ? 3'b111 : node538;
											assign node538 = (inp[6]) ? 3'b110 : 3'b111;
									assign node542 = (inp[6]) ? node544 : 3'b110;
										assign node544 = (inp[7]) ? node546 : 3'b110;
											assign node546 = (inp[1]) ? 3'b110 : 3'b111;
							assign node549 = (inp[1]) ? node571 : node550;
								assign node550 = (inp[9]) ? node560 : node551;
									assign node551 = (inp[2]) ? node553 : 3'b110;
										assign node553 = (inp[7]) ? node557 : node554;
											assign node554 = (inp[6]) ? 3'b110 : 3'b110;
											assign node557 = (inp[0]) ? 3'b110 : 3'b111;
									assign node560 = (inp[6]) ? node566 : node561;
										assign node561 = (inp[7]) ? 3'b111 : node562;
											assign node562 = (inp[2]) ? 3'b110 : 3'b111;
										assign node566 = (inp[2]) ? 3'b111 : node567;
											assign node567 = (inp[0]) ? 3'b110 : 3'b110;
								assign node571 = (inp[2]) ? node573 : 3'b111;
									assign node573 = (inp[7]) ? 3'b111 : node574;
										assign node574 = (inp[0]) ? node578 : node575;
											assign node575 = (inp[6]) ? 3'b111 : 3'b110;
											assign node578 = (inp[6]) ? 3'b110 : 3'b111;
					assign node582 = (inp[10]) ? node656 : node583;
						assign node583 = (inp[2]) ? node627 : node584;
							assign node584 = (inp[0]) ? node606 : node585;
								assign node585 = (inp[1]) ? node593 : node586;
									assign node586 = (inp[6]) ? node588 : 3'b110;
										assign node588 = (inp[3]) ? 3'b110 : node589;
											assign node589 = (inp[9]) ? 3'b110 : 3'b111;
									assign node593 = (inp[3]) ? node601 : node594;
										assign node594 = (inp[9]) ? node598 : node595;
											assign node595 = (inp[7]) ? 3'b111 : 3'b110;
											assign node598 = (inp[7]) ? 3'b110 : 3'b111;
										assign node601 = (inp[6]) ? 3'b110 : node602;
											assign node602 = (inp[9]) ? 3'b111 : 3'b110;
								assign node606 = (inp[3]) ? node620 : node607;
									assign node607 = (inp[6]) ? node613 : node608;
										assign node608 = (inp[1]) ? node610 : 3'b111;
											assign node610 = (inp[7]) ? 3'b110 : 3'b111;
										assign node613 = (inp[1]) ? node617 : node614;
											assign node614 = (inp[7]) ? 3'b110 : 3'b111;
											assign node617 = (inp[7]) ? 3'b111 : 3'b110;
									assign node620 = (inp[7]) ? 3'b111 : node621;
										assign node621 = (inp[6]) ? 3'b111 : node622;
											assign node622 = (inp[1]) ? 3'b110 : 3'b111;
							assign node627 = (inp[0]) ? node645 : node628;
								assign node628 = (inp[1]) ? node634 : node629;
									assign node629 = (inp[7]) ? node631 : 3'b111;
										assign node631 = (inp[3]) ? 3'b111 : 3'b110;
									assign node634 = (inp[7]) ? node640 : node635;
										assign node635 = (inp[3]) ? 3'b110 : node636;
											assign node636 = (inp[6]) ? 3'b110 : 3'b111;
										assign node640 = (inp[3]) ? 3'b111 : node641;
											assign node641 = (inp[6]) ? 3'b111 : 3'b110;
								assign node645 = (inp[3]) ? 3'b110 : node646;
									assign node646 = (inp[7]) ? node648 : 3'b110;
										assign node648 = (inp[1]) ? node652 : node649;
											assign node649 = (inp[6]) ? 3'b111 : 3'b110;
											assign node652 = (inp[6]) ? 3'b110 : 3'b111;
						assign node656 = (inp[7]) ? node692 : node657;
							assign node657 = (inp[2]) ? node675 : node658;
								assign node658 = (inp[0]) ? node668 : node659;
									assign node659 = (inp[3]) ? 3'b100 : node660;
										assign node660 = (inp[6]) ? node664 : node661;
											assign node661 = (inp[1]) ? 3'b100 : 3'b101;
											assign node664 = (inp[1]) ? 3'b101 : 3'b100;
									assign node668 = (inp[3]) ? 3'b101 : node669;
										assign node669 = (inp[9]) ? node671 : 3'b101;
											assign node671 = (inp[6]) ? 3'b100 : 3'b100;
								assign node675 = (inp[0]) ? node683 : node676;
									assign node676 = (inp[3]) ? 3'b101 : node677;
										assign node677 = (inp[9]) ? 3'b101 : node678;
											assign node678 = (inp[1]) ? 3'b100 : 3'b100;
									assign node683 = (inp[3]) ? 3'b100 : node684;
										assign node684 = (inp[1]) ? node688 : node685;
											assign node685 = (inp[6]) ? 3'b100 : 3'b101;
											assign node688 = (inp[6]) ? 3'b101 : 3'b100;
							assign node692 = (inp[9]) ? node710 : node693;
								assign node693 = (inp[0]) ? node703 : node694;
									assign node694 = (inp[2]) ? node698 : node695;
										assign node695 = (inp[1]) ? 3'b100 : 3'b101;
										assign node698 = (inp[1]) ? 3'b101 : node699;
											assign node699 = (inp[6]) ? 3'b101 : 3'b100;
									assign node703 = (inp[2]) ? 3'b100 : node704;
										assign node704 = (inp[1]) ? 3'b101 : node705;
											assign node705 = (inp[6]) ? 3'b100 : 3'b100;
								assign node710 = (inp[0]) ? node718 : node711;
									assign node711 = (inp[2]) ? node713 : 3'b100;
										assign node713 = (inp[1]) ? 3'b101 : node714;
											assign node714 = (inp[6]) ? 3'b101 : 3'b100;
									assign node718 = (inp[2]) ? node724 : node719;
										assign node719 = (inp[1]) ? 3'b101 : node720;
											assign node720 = (inp[6]) ? 3'b100 : 3'b100;
										assign node724 = (inp[1]) ? 3'b100 : node725;
											assign node725 = (inp[6]) ? 3'b100 : 3'b100;
			assign node729 = (inp[4]) ? node1085 : node730;
				assign node730 = (inp[6]) ? node918 : node731;
					assign node731 = (inp[10]) ? node815 : node732;
						assign node732 = (inp[0]) ? node776 : node733;
							assign node733 = (inp[7]) ? node749 : node734;
								assign node734 = (inp[3]) ? node742 : node735;
									assign node735 = (inp[9]) ? node739 : node736;
										assign node736 = (inp[1]) ? 3'b101 : 3'b100;
										assign node739 = (inp[1]) ? 3'b100 : 3'b101;
									assign node742 = (inp[9]) ? node746 : node743;
										assign node743 = (inp[11]) ? 3'b111 : 3'b110;
										assign node746 = (inp[1]) ? 3'b110 : 3'b111;
								assign node749 = (inp[3]) ? node763 : node750;
									assign node750 = (inp[9]) ? node756 : node751;
										assign node751 = (inp[1]) ? 3'b111 : node752;
											assign node752 = (inp[11]) ? 3'b110 : 3'b110;
										assign node756 = (inp[1]) ? node760 : node757;
											assign node757 = (inp[2]) ? 3'b110 : 3'b111;
											assign node760 = (inp[11]) ? 3'b110 : 3'b110;
									assign node763 = (inp[1]) ? node771 : node764;
										assign node764 = (inp[9]) ? node768 : node765;
											assign node765 = (inp[2]) ? 3'b100 : 3'b101;
											assign node768 = (inp[2]) ? 3'b101 : 3'b100;
										assign node771 = (inp[11]) ? 3'b100 : node772;
											assign node772 = (inp[9]) ? 3'b100 : 3'b100;
							assign node776 = (inp[1]) ? node798 : node777;
								assign node777 = (inp[9]) ? node787 : node778;
									assign node778 = (inp[7]) ? node782 : node779;
										assign node779 = (inp[3]) ? 3'b110 : 3'b100;
										assign node782 = (inp[3]) ? 3'b101 : node783;
											assign node783 = (inp[11]) ? 3'b111 : 3'b110;
									assign node787 = (inp[7]) ? node791 : node788;
										assign node788 = (inp[3]) ? 3'b111 : 3'b101;
										assign node791 = (inp[3]) ? node795 : node792;
											assign node792 = (inp[11]) ? 3'b110 : 3'b111;
											assign node795 = (inp[2]) ? 3'b101 : 3'b100;
								assign node798 = (inp[9]) ? node806 : node799;
									assign node799 = (inp[3]) ? node803 : node800;
										assign node800 = (inp[7]) ? 3'b111 : 3'b101;
										assign node803 = (inp[7]) ? 3'b101 : 3'b111;
									assign node806 = (inp[7]) ? node810 : node807;
										assign node807 = (inp[3]) ? 3'b110 : 3'b100;
										assign node810 = (inp[3]) ? 3'b101 : node811;
											assign node811 = (inp[2]) ? 3'b111 : 3'b110;
						assign node815 = (inp[1]) ? node869 : node816;
							assign node816 = (inp[9]) ? node846 : node817;
								assign node817 = (inp[11]) ? node833 : node818;
									assign node818 = (inp[2]) ? node826 : node819;
										assign node819 = (inp[0]) ? node823 : node820;
											assign node820 = (inp[3]) ? 3'b100 : 3'b100;
											assign node823 = (inp[3]) ? 3'b100 : 3'b100;
										assign node826 = (inp[7]) ? node830 : node827;
											assign node827 = (inp[3]) ? 3'b111 : 3'b101;
											assign node830 = (inp[3]) ? 3'b100 : 3'b111;
									assign node833 = (inp[2]) ? node839 : node834;
										assign node834 = (inp[3]) ? node836 : 3'b110;
											assign node836 = (inp[7]) ? 3'b101 : 3'b111;
										assign node839 = (inp[3]) ? node843 : node840;
											assign node840 = (inp[7]) ? 3'b110 : 3'b100;
											assign node843 = (inp[7]) ? 3'b100 : 3'b110;
								assign node846 = (inp[7]) ? node858 : node847;
									assign node847 = (inp[3]) ? node853 : node848;
										assign node848 = (inp[11]) ? 3'b100 : node849;
											assign node849 = (inp[2]) ? 3'b100 : 3'b101;
										assign node853 = (inp[11]) ? node855 : 3'b110;
											assign node855 = (inp[2]) ? 3'b111 : 3'b110;
									assign node858 = (inp[3]) ? node864 : node859;
										assign node859 = (inp[2]) ? node861 : 3'b111;
											assign node861 = (inp[11]) ? 3'b111 : 3'b110;
										assign node864 = (inp[2]) ? 3'b101 : node865;
											assign node865 = (inp[11]) ? 3'b100 : 3'b101;
							assign node869 = (inp[9]) ? node895 : node870;
								assign node870 = (inp[0]) ? node882 : node871;
									assign node871 = (inp[3]) ? node875 : node872;
										assign node872 = (inp[7]) ? 3'b111 : 3'b101;
										assign node875 = (inp[7]) ? node879 : node876;
											assign node876 = (inp[11]) ? 3'b110 : 3'b110;
											assign node879 = (inp[2]) ? 3'b101 : 3'b100;
									assign node882 = (inp[7]) ? node888 : node883;
										assign node883 = (inp[3]) ? node885 : 3'b100;
											assign node885 = (inp[11]) ? 3'b110 : 3'b110;
										assign node888 = (inp[3]) ? node892 : node889;
											assign node889 = (inp[11]) ? 3'b111 : 3'b110;
											assign node892 = (inp[11]) ? 3'b100 : 3'b101;
								assign node895 = (inp[0]) ? node909 : node896;
									assign node896 = (inp[3]) ? node904 : node897;
										assign node897 = (inp[7]) ? node901 : node898;
											assign node898 = (inp[11]) ? 3'b100 : 3'b100;
											assign node901 = (inp[11]) ? 3'b110 : 3'b110;
										assign node904 = (inp[7]) ? node906 : 3'b110;
											assign node906 = (inp[2]) ? 3'b100 : 3'b101;
									assign node909 = (inp[2]) ? 3'b111 : node910;
										assign node910 = (inp[11]) ? node914 : node911;
											assign node911 = (inp[7]) ? 3'b100 : 3'b110;
											assign node914 = (inp[3]) ? 3'b101 : 3'b100;
					assign node918 = (inp[1]) ? node1000 : node919;
						assign node919 = (inp[10]) ? node961 : node920;
							assign node920 = (inp[9]) ? node942 : node921;
								assign node921 = (inp[7]) ? node931 : node922;
									assign node922 = (inp[3]) ? node926 : node923;
										assign node923 = (inp[11]) ? 3'b010 : 3'b000;
										assign node926 = (inp[11]) ? node928 : 3'b010;
											assign node928 = (inp[0]) ? 3'b001 : 3'b000;
									assign node931 = (inp[11]) ? node937 : node932;
										assign node932 = (inp[3]) ? 3'b010 : node933;
											assign node933 = (inp[2]) ? 3'b001 : 3'b000;
										assign node937 = (inp[3]) ? node939 : 3'b011;
											assign node939 = (inp[2]) ? 3'b001 : 3'b000;
								assign node942 = (inp[11]) ? node954 : node943;
									assign node943 = (inp[3]) ? node949 : node944;
										assign node944 = (inp[2]) ? node946 : 3'b001;
											assign node946 = (inp[7]) ? 3'b000 : 3'b001;
										assign node949 = (inp[2]) ? 3'b011 : node950;
											assign node950 = (inp[7]) ? 3'b010 : 3'b011;
									assign node954 = (inp[3]) ? node958 : node955;
										assign node955 = (inp[7]) ? 3'b010 : 3'b011;
										assign node958 = (inp[2]) ? 3'b000 : 3'b001;
							assign node961 = (inp[9]) ? node983 : node962;
								assign node962 = (inp[2]) ? node972 : node963;
									assign node963 = (inp[3]) ? node969 : node964;
										assign node964 = (inp[11]) ? node966 : 3'b001;
											assign node966 = (inp[7]) ? 3'b011 : 3'b010;
										assign node969 = (inp[11]) ? 3'b000 : 3'b010;
									assign node972 = (inp[3]) ? node980 : node973;
										assign node973 = (inp[11]) ? node977 : node974;
											assign node974 = (inp[7]) ? 3'b000 : 3'b001;
											assign node977 = (inp[7]) ? 3'b011 : 3'b010;
										assign node980 = (inp[11]) ? 3'b001 : 3'b011;
								assign node983 = (inp[3]) ? node993 : node984;
									assign node984 = (inp[11]) ? node990 : node985;
										assign node985 = (inp[2]) ? node987 : 3'b000;
											assign node987 = (inp[7]) ? 3'b001 : 3'b000;
										assign node990 = (inp[7]) ? 3'b010 : 3'b011;
									assign node993 = (inp[2]) ? node997 : node994;
										assign node994 = (inp[11]) ? 3'b001 : 3'b011;
										assign node997 = (inp[11]) ? 3'b000 : 3'b010;
						assign node1000 = (inp[10]) ? node1050 : node1001;
							assign node1001 = (inp[9]) ? node1021 : node1002;
								assign node1002 = (inp[7]) ? node1012 : node1003;
									assign node1003 = (inp[11]) ? node1007 : node1004;
										assign node1004 = (inp[3]) ? 3'b010 : 3'b000;
										assign node1007 = (inp[2]) ? 3'b001 : node1008;
											assign node1008 = (inp[3]) ? 3'b000 : 3'b010;
									assign node1012 = (inp[2]) ? 3'b001 : node1013;
										assign node1013 = (inp[3]) ? node1017 : node1014;
											assign node1014 = (inp[11]) ? 3'b011 : 3'b000;
											assign node1017 = (inp[11]) ? 3'b000 : 3'b011;
								assign node1021 = (inp[7]) ? node1037 : node1022;
									assign node1022 = (inp[2]) ? node1030 : node1023;
										assign node1023 = (inp[0]) ? node1027 : node1024;
											assign node1024 = (inp[3]) ? 3'b001 : 3'b001;
											assign node1027 = (inp[3]) ? 3'b001 : 3'b001;
										assign node1030 = (inp[3]) ? node1034 : node1031;
											assign node1031 = (inp[11]) ? 3'b011 : 3'b001;
											assign node1034 = (inp[11]) ? 3'b000 : 3'b011;
									assign node1037 = (inp[11]) ? node1045 : node1038;
										assign node1038 = (inp[3]) ? node1042 : node1039;
											assign node1039 = (inp[2]) ? 3'b000 : 3'b001;
											assign node1042 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1045 = (inp[3]) ? node1047 : 3'b010;
											assign node1047 = (inp[2]) ? 3'b000 : 3'b001;
							assign node1050 = (inp[9]) ? node1066 : node1051;
								assign node1051 = (inp[11]) ? node1059 : node1052;
									assign node1052 = (inp[3]) ? 3'b011 : node1053;
										assign node1053 = (inp[2]) ? node1055 : 3'b001;
											assign node1055 = (inp[7]) ? 3'b000 : 3'b001;
									assign node1059 = (inp[3]) ? node1063 : node1060;
										assign node1060 = (inp[7]) ? 3'b011 : 3'b010;
										assign node1063 = (inp[2]) ? 3'b001 : 3'b000;
								assign node1066 = (inp[11]) ? node1078 : node1067;
									assign node1067 = (inp[3]) ? node1073 : node1068;
										assign node1068 = (inp[7]) ? node1070 : 3'b000;
											assign node1070 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1073 = (inp[7]) ? node1075 : 3'b010;
											assign node1075 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1078 = (inp[3]) ? node1082 : node1079;
										assign node1079 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1082 = (inp[2]) ? 3'b000 : 3'b001;
				assign node1085 = (inp[11]) ? node1229 : node1086;
					assign node1086 = (inp[7]) ? node1146 : node1087;
						assign node1087 = (inp[6]) ? node1113 : node1088;
							assign node1088 = (inp[1]) ? node1102 : node1089;
								assign node1089 = (inp[2]) ? node1097 : node1090;
									assign node1090 = (inp[9]) ? 3'b000 : node1091;
										assign node1091 = (inp[3]) ? node1093 : 3'b000;
											assign node1093 = (inp[10]) ? 3'b001 : 3'b000;
									assign node1097 = (inp[3]) ? node1099 : 3'b001;
										assign node1099 = (inp[10]) ? 3'b000 : 3'b001;
								assign node1102 = (inp[2]) ? node1108 : node1103;
									assign node1103 = (inp[10]) ? node1105 : 3'b001;
										assign node1105 = (inp[3]) ? 3'b000 : 3'b001;
									assign node1108 = (inp[3]) ? node1110 : 3'b000;
										assign node1110 = (inp[10]) ? 3'b001 : 3'b000;
							assign node1113 = (inp[0]) ? node1127 : node1114;
								assign node1114 = (inp[9]) ? node1122 : node1115;
									assign node1115 = (inp[10]) ? node1119 : node1116;
										assign node1116 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1119 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1122 = (inp[2]) ? 3'b010 : node1123;
										assign node1123 = (inp[10]) ? 3'b011 : 3'b010;
								assign node1127 = (inp[3]) ? node1141 : node1128;
									assign node1128 = (inp[1]) ? node1136 : node1129;
										assign node1129 = (inp[10]) ? node1133 : node1130;
											assign node1130 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1133 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1136 = (inp[2]) ? node1138 : 3'b010;
											assign node1138 = (inp[10]) ? 3'b010 : 3'b011;
									assign node1141 = (inp[10]) ? 3'b010 : node1142;
										assign node1142 = (inp[2]) ? 3'b011 : 3'b010;
						assign node1146 = (inp[3]) ? node1192 : node1147;
							assign node1147 = (inp[9]) ? node1163 : node1148;
								assign node1148 = (inp[10]) ? node1156 : node1149;
									assign node1149 = (inp[2]) ? 3'b011 : node1150;
										assign node1150 = (inp[6]) ? 3'b010 : node1151;
											assign node1151 = (inp[1]) ? 3'b011 : 3'b010;
									assign node1156 = (inp[2]) ? node1158 : 3'b011;
										assign node1158 = (inp[1]) ? 3'b010 : node1159;
											assign node1159 = (inp[6]) ? 3'b010 : 3'b011;
								assign node1163 = (inp[0]) ? node1177 : node1164;
									assign node1164 = (inp[6]) ? node1172 : node1165;
										assign node1165 = (inp[2]) ? node1169 : node1166;
											assign node1166 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1169 = (inp[1]) ? 3'b010 : 3'b011;
										assign node1172 = (inp[2]) ? node1174 : 3'b010;
											assign node1174 = (inp[1]) ? 3'b010 : 3'b011;
									assign node1177 = (inp[6]) ? node1185 : node1178;
										assign node1178 = (inp[10]) ? node1182 : node1179;
											assign node1179 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1182 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1185 = (inp[2]) ? node1189 : node1186;
											assign node1186 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1189 = (inp[10]) ? 3'b010 : 3'b011;
							assign node1192 = (inp[6]) ? node1222 : node1193;
								assign node1193 = (inp[2]) ? node1207 : node1194;
									assign node1194 = (inp[9]) ? node1202 : node1195;
										assign node1195 = (inp[0]) ? node1199 : node1196;
											assign node1196 = (inp[1]) ? 3'b010 : 3'b010;
											assign node1199 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1202 = (inp[0]) ? 3'b010 : node1203;
											assign node1203 = (inp[10]) ? 3'b010 : 3'b010;
									assign node1207 = (inp[9]) ? node1215 : node1208;
										assign node1208 = (inp[0]) ? node1212 : node1209;
											assign node1209 = (inp[10]) ? 3'b010 : 3'b010;
											assign node1212 = (inp[10]) ? 3'b010 : 3'b010;
										assign node1215 = (inp[0]) ? node1219 : node1216;
											assign node1216 = (inp[1]) ? 3'b010 : 3'b010;
											assign node1219 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1222 = (inp[2]) ? node1226 : node1223;
									assign node1223 = (inp[10]) ? 3'b011 : 3'b010;
									assign node1226 = (inp[10]) ? 3'b010 : 3'b011;
					assign node1229 = (inp[7]) ? node1297 : node1230;
						assign node1230 = (inp[6]) ? node1266 : node1231;
							assign node1231 = (inp[3]) ? node1259 : node1232;
								assign node1232 = (inp[1]) ? node1248 : node1233;
									assign node1233 = (inp[9]) ? node1241 : node1234;
										assign node1234 = (inp[2]) ? node1238 : node1235;
											assign node1235 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1238 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1241 = (inp[2]) ? node1245 : node1242;
											assign node1242 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1245 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1248 = (inp[9]) ? node1254 : node1249;
										assign node1249 = (inp[2]) ? node1251 : 3'b011;
											assign node1251 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1254 = (inp[2]) ? 3'b011 : node1255;
											assign node1255 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1259 = (inp[2]) ? node1263 : node1260;
									assign node1260 = (inp[1]) ? 3'b011 : 3'b010;
									assign node1263 = (inp[1]) ? 3'b010 : 3'b011;
							assign node1266 = (inp[1]) ? node1274 : node1267;
								assign node1267 = (inp[3]) ? node1271 : node1268;
									assign node1268 = (inp[2]) ? 3'b001 : 3'b000;
									assign node1271 = (inp[2]) ? 3'b000 : 3'b001;
								assign node1274 = (inp[0]) ? node1284 : node1275;
									assign node1275 = (inp[10]) ? node1277 : 3'b001;
										assign node1277 = (inp[3]) ? node1281 : node1278;
											assign node1278 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1281 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1284 = (inp[9]) ? node1290 : node1285;
										assign node1285 = (inp[2]) ? node1287 : 3'b000;
											assign node1287 = (inp[3]) ? 3'b000 : 3'b001;
										assign node1290 = (inp[3]) ? node1294 : node1291;
											assign node1291 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1294 = (inp[2]) ? 3'b000 : 3'b001;
						assign node1297 = (inp[2]) ? node1311 : node1298;
							assign node1298 = (inp[6]) ? 3'b001 : node1299;
								assign node1299 = (inp[1]) ? node1305 : node1300;
									assign node1300 = (inp[3]) ? 3'b000 : node1301;
										assign node1301 = (inp[10]) ? 3'b000 : 3'b001;
									assign node1305 = (inp[10]) ? 3'b001 : node1306;
										assign node1306 = (inp[3]) ? 3'b001 : 3'b000;
							assign node1311 = (inp[6]) ? 3'b000 : node1312;
								assign node1312 = (inp[1]) ? node1318 : node1313;
									assign node1313 = (inp[10]) ? 3'b001 : node1314;
										assign node1314 = (inp[3]) ? 3'b001 : 3'b000;
									assign node1318 = (inp[3]) ? 3'b000 : node1319;
										assign node1319 = (inp[10]) ? 3'b000 : 3'b001;
		assign node1324 = (inp[4]) ? node1978 : node1325;
			assign node1325 = (inp[6]) ? node1701 : node1326;
				assign node1326 = (inp[8]) ? node1528 : node1327;
					assign node1327 = (inp[1]) ? node1433 : node1328;
						assign node1328 = (inp[11]) ? node1386 : node1329;
							assign node1329 = (inp[9]) ? node1359 : node1330;
								assign node1330 = (inp[2]) ? node1344 : node1331;
									assign node1331 = (inp[0]) ? node1337 : node1332;
										assign node1332 = (inp[7]) ? node1334 : 3'b101;
											assign node1334 = (inp[3]) ? 3'b100 : 3'b100;
										assign node1337 = (inp[3]) ? node1341 : node1338;
											assign node1338 = (inp[10]) ? 3'b111 : 3'b101;
											assign node1341 = (inp[10]) ? 3'b100 : 3'b111;
									assign node1344 = (inp[0]) ? node1352 : node1345;
										assign node1345 = (inp[7]) ? node1349 : node1346;
											assign node1346 = (inp[3]) ? 3'b100 : 3'b111;
											assign node1349 = (inp[10]) ? 3'b101 : 3'b111;
										assign node1352 = (inp[7]) ? node1356 : node1353;
											assign node1353 = (inp[3]) ? 3'b101 : 3'b100;
											assign node1356 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1359 = (inp[2]) ? node1375 : node1360;
									assign node1360 = (inp[0]) ? node1368 : node1361;
										assign node1361 = (inp[3]) ? node1365 : node1362;
											assign node1362 = (inp[10]) ? 3'b111 : 3'b101;
											assign node1365 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1368 = (inp[3]) ? node1372 : node1369;
											assign node1369 = (inp[10]) ? 3'b110 : 3'b100;
											assign node1372 = (inp[10]) ? 3'b100 : 3'b110;
									assign node1375 = (inp[7]) ? node1381 : node1376;
										assign node1376 = (inp[3]) ? node1378 : 3'b100;
											assign node1378 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1381 = (inp[0]) ? node1383 : 3'b100;
											assign node1383 = (inp[3]) ? 3'b101 : 3'b101;
							assign node1386 = (inp[3]) ? node1408 : node1387;
								assign node1387 = (inp[10]) ? node1395 : node1388;
									assign node1388 = (inp[7]) ? 3'b101 : node1389;
										assign node1389 = (inp[2]) ? node1391 : 3'b111;
											assign node1391 = (inp[0]) ? 3'b110 : 3'b110;
									assign node1395 = (inp[7]) ? node1401 : node1396;
										assign node1396 = (inp[0]) ? 3'b100 : node1397;
											assign node1397 = (inp[2]) ? 3'b100 : 3'b101;
										assign node1401 = (inp[2]) ? node1405 : node1402;
											assign node1402 = (inp[9]) ? 3'b110 : 3'b110;
											assign node1405 = (inp[9]) ? 3'b110 : 3'b110;
								assign node1408 = (inp[2]) ? node1418 : node1409;
									assign node1409 = (inp[10]) ? node1413 : node1410;
										assign node1410 = (inp[7]) ? 3'b110 : 3'b100;
										assign node1413 = (inp[7]) ? 3'b101 : node1414;
											assign node1414 = (inp[0]) ? 3'b110 : 3'b110;
									assign node1418 = (inp[0]) ? node1426 : node1419;
										assign node1419 = (inp[9]) ? node1423 : node1420;
											assign node1420 = (inp[10]) ? 3'b101 : 3'b100;
											assign node1423 = (inp[10]) ? 3'b100 : 3'b111;
										assign node1426 = (inp[7]) ? node1430 : node1427;
											assign node1427 = (inp[9]) ? 3'b111 : 3'b101;
											assign node1430 = (inp[10]) ? 3'b100 : 3'b111;
						assign node1433 = (inp[10]) ? node1473 : node1434;
							assign node1434 = (inp[3]) ? node1450 : node1435;
								assign node1435 = (inp[11]) ? node1443 : node1436;
									assign node1436 = (inp[0]) ? node1440 : node1437;
										assign node1437 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1440 = (inp[9]) ? 3'b100 : 3'b101;
									assign node1443 = (inp[7]) ? node1445 : 3'b110;
										assign node1445 = (inp[0]) ? node1447 : 3'b101;
											assign node1447 = (inp[9]) ? 3'b101 : 3'b100;
								assign node1450 = (inp[11]) ? node1462 : node1451;
									assign node1451 = (inp[2]) ? node1457 : node1452;
										assign node1452 = (inp[9]) ? node1454 : 3'b110;
											assign node1454 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1457 = (inp[7]) ? node1459 : 3'b111;
											assign node1459 = (inp[0]) ? 3'b111 : 3'b110;
									assign node1462 = (inp[7]) ? node1468 : node1463;
										assign node1463 = (inp[0]) ? 3'b100 : node1464;
											assign node1464 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1468 = (inp[9]) ? 3'b110 : node1469;
											assign node1469 = (inp[0]) ? 3'b111 : 3'b110;
							assign node1473 = (inp[3]) ? node1501 : node1474;
								assign node1474 = (inp[7]) ? node1488 : node1475;
									assign node1475 = (inp[11]) ? node1481 : node1476;
										assign node1476 = (inp[2]) ? 3'b110 : node1477;
											assign node1477 = (inp[0]) ? 3'b110 : 3'b111;
										assign node1481 = (inp[9]) ? node1485 : node1482;
											assign node1482 = (inp[0]) ? 3'b100 : 3'b100;
											assign node1485 = (inp[0]) ? 3'b100 : 3'b101;
									assign node1488 = (inp[11]) ? node1496 : node1489;
										assign node1489 = (inp[2]) ? node1493 : node1490;
											assign node1490 = (inp[9]) ? 3'b110 : 3'b110;
											assign node1493 = (inp[0]) ? 3'b110 : 3'b110;
										assign node1496 = (inp[0]) ? 3'b110 : node1497;
											assign node1497 = (inp[9]) ? 3'b111 : 3'b110;
								assign node1501 = (inp[7]) ? node1515 : node1502;
									assign node1502 = (inp[11]) ? node1508 : node1503;
										assign node1503 = (inp[2]) ? 3'b100 : node1504;
											assign node1504 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1508 = (inp[0]) ? node1512 : node1509;
											assign node1509 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1512 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1515 = (inp[11]) ? node1523 : node1516;
										assign node1516 = (inp[0]) ? node1520 : node1517;
											assign node1517 = (inp[9]) ? 3'b101 : 3'b100;
											assign node1520 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1523 = (inp[0]) ? node1525 : 3'b100;
											assign node1525 = (inp[9]) ? 3'b100 : 3'b101;
					assign node1528 = (inp[1]) ? node1608 : node1529;
						assign node1529 = (inp[9]) ? node1571 : node1530;
							assign node1530 = (inp[11]) ? node1554 : node1531;
								assign node1531 = (inp[10]) ? node1545 : node1532;
									assign node1532 = (inp[2]) ? node1538 : node1533;
										assign node1533 = (inp[0]) ? 3'b110 : node1534;
											assign node1534 = (inp[7]) ? 3'b100 : 3'b110;
										assign node1538 = (inp[7]) ? node1542 : node1539;
											assign node1539 = (inp[3]) ? 3'b110 : 3'b101;
											assign node1542 = (inp[3]) ? 3'b101 : 3'b111;
									assign node1545 = (inp[3]) ? node1549 : node1546;
										assign node1546 = (inp[7]) ? 3'b110 : 3'b100;
										assign node1549 = (inp[7]) ? 3'b100 : node1550;
											assign node1550 = (inp[2]) ? 3'b110 : 3'b111;
								assign node1554 = (inp[10]) ? node1562 : node1555;
									assign node1555 = (inp[7]) ? node1559 : node1556;
										assign node1556 = (inp[3]) ? 3'b110 : 3'b100;
										assign node1559 = (inp[2]) ? 3'b100 : 3'b101;
									assign node1562 = (inp[7]) ? node1568 : node1563;
										assign node1563 = (inp[3]) ? 3'b110 : node1564;
											assign node1564 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1568 = (inp[3]) ? 3'b100 : 3'b110;
							assign node1571 = (inp[2]) ? node1591 : node1572;
								assign node1572 = (inp[3]) ? node1580 : node1573;
									assign node1573 = (inp[7]) ? node1575 : 3'b101;
										assign node1575 = (inp[10]) ? 3'b111 : node1576;
											assign node1576 = (inp[11]) ? 3'b110 : 3'b111;
									assign node1580 = (inp[7]) ? node1586 : node1581;
										assign node1581 = (inp[10]) ? node1583 : 3'b111;
											assign node1583 = (inp[11]) ? 3'b111 : 3'b110;
										assign node1586 = (inp[11]) ? node1588 : 3'b101;
											assign node1588 = (inp[10]) ? 3'b101 : 3'b100;
								assign node1591 = (inp[11]) ? node1601 : node1592;
									assign node1592 = (inp[10]) ? node1594 : 3'b100;
										assign node1594 = (inp[0]) ? node1598 : node1595;
											assign node1595 = (inp[7]) ? 3'b101 : 3'b101;
											assign node1598 = (inp[7]) ? 3'b101 : 3'b101;
									assign node1601 = (inp[7]) ? node1605 : node1602;
										assign node1602 = (inp[3]) ? 3'b111 : 3'b101;
										assign node1605 = (inp[3]) ? 3'b101 : 3'b111;
						assign node1608 = (inp[9]) ? node1660 : node1609;
							assign node1609 = (inp[11]) ? node1633 : node1610;
								assign node1610 = (inp[0]) ? node1624 : node1611;
									assign node1611 = (inp[2]) ? node1619 : node1612;
										assign node1612 = (inp[3]) ? node1616 : node1613;
											assign node1613 = (inp[7]) ? 3'b111 : 3'b101;
											assign node1616 = (inp[7]) ? 3'b101 : 3'b110;
										assign node1619 = (inp[3]) ? node1621 : 3'b110;
											assign node1621 = (inp[10]) ? 3'b101 : 3'b111;
									assign node1624 = (inp[7]) ? node1628 : node1625;
										assign node1625 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1628 = (inp[2]) ? node1630 : 3'b111;
											assign node1630 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1633 = (inp[10]) ? node1647 : node1634;
									assign node1634 = (inp[2]) ? node1640 : node1635;
										assign node1635 = (inp[0]) ? node1637 : 3'b110;
											assign node1637 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1640 = (inp[7]) ? node1644 : node1641;
											assign node1641 = (inp[3]) ? 3'b111 : 3'b101;
											assign node1644 = (inp[3]) ? 3'b101 : 3'b111;
									assign node1647 = (inp[2]) ? node1655 : node1648;
										assign node1648 = (inp[3]) ? node1652 : node1649;
											assign node1649 = (inp[7]) ? 3'b111 : 3'b101;
											assign node1652 = (inp[7]) ? 3'b101 : 3'b111;
										assign node1655 = (inp[7]) ? 3'b111 : node1656;
											assign node1656 = (inp[3]) ? 3'b111 : 3'b100;
							assign node1660 = (inp[10]) ? node1686 : node1661;
								assign node1661 = (inp[7]) ? node1671 : node1662;
									assign node1662 = (inp[3]) ? node1666 : node1663;
										assign node1663 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1666 = (inp[11]) ? node1668 : 3'b110;
											assign node1668 = (inp[2]) ? 3'b110 : 3'b111;
									assign node1671 = (inp[3]) ? node1679 : node1672;
										assign node1672 = (inp[11]) ? node1676 : node1673;
											assign node1673 = (inp[2]) ? 3'b111 : 3'b110;
											assign node1676 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1679 = (inp[11]) ? node1683 : node1680;
											assign node1680 = (inp[2]) ? 3'b101 : 3'b100;
											assign node1683 = (inp[2]) ? 3'b100 : 3'b101;
								assign node1686 = (inp[7]) ? node1698 : node1687;
									assign node1687 = (inp[3]) ? node1693 : node1688;
										assign node1688 = (inp[0]) ? 3'b100 : node1689;
											assign node1689 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1693 = (inp[2]) ? 3'b110 : node1694;
											assign node1694 = (inp[11]) ? 3'b110 : 3'b111;
									assign node1698 = (inp[3]) ? 3'b100 : 3'b110;
				assign node1701 = (inp[3]) ? node1859 : node1702;
					assign node1702 = (inp[8]) ? node1804 : node1703;
						assign node1703 = (inp[10]) ? node1757 : node1704;
							assign node1704 = (inp[11]) ? node1732 : node1705;
								assign node1705 = (inp[7]) ? node1719 : node1706;
									assign node1706 = (inp[0]) ? node1714 : node1707;
										assign node1707 = (inp[9]) ? node1711 : node1708;
											assign node1708 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1711 = (inp[2]) ? 3'b010 : 3'b010;
										assign node1714 = (inp[9]) ? 3'b011 : node1715;
											assign node1715 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1719 = (inp[1]) ? node1727 : node1720;
										assign node1720 = (inp[2]) ? node1724 : node1721;
											assign node1721 = (inp[0]) ? 3'b000 : 3'b000;
											assign node1724 = (inp[0]) ? 3'b000 : 3'b001;
										assign node1727 = (inp[9]) ? node1729 : 3'b001;
											assign node1729 = (inp[0]) ? 3'b000 : 3'b001;
								assign node1732 = (inp[0]) ? node1748 : node1733;
									assign node1733 = (inp[1]) ? node1741 : node1734;
										assign node1734 = (inp[7]) ? node1738 : node1735;
											assign node1735 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1738 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1741 = (inp[2]) ? node1745 : node1742;
											assign node1742 = (inp[7]) ? 3'b000 : 3'b000;
											assign node1745 = (inp[9]) ? 3'b000 : 3'b000;
									assign node1748 = (inp[2]) ? 3'b000 : node1749;
										assign node1749 = (inp[7]) ? node1753 : node1750;
											assign node1750 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1753 = (inp[9]) ? 3'b001 : 3'b000;
							assign node1757 = (inp[7]) ? node1779 : node1758;
								assign node1758 = (inp[11]) ? node1766 : node1759;
									assign node1759 = (inp[9]) ? node1761 : 3'b000;
										assign node1761 = (inp[0]) ? 3'b000 : node1762;
											assign node1762 = (inp[1]) ? 3'b001 : 3'b000;
									assign node1766 = (inp[9]) ? node1772 : node1767;
										assign node1767 = (inp[1]) ? 3'b011 : node1768;
											assign node1768 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1772 = (inp[2]) ? node1776 : node1773;
											assign node1773 = (inp[1]) ? 3'b010 : 3'b010;
											assign node1776 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1779 = (inp[2]) ? node1793 : node1780;
									assign node1780 = (inp[11]) ? node1786 : node1781;
										assign node1781 = (inp[0]) ? node1783 : 3'b011;
											assign node1783 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1786 = (inp[0]) ? node1790 : node1787;
											assign node1787 = (inp[1]) ? 3'b010 : 3'b010;
											assign node1790 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1793 = (inp[1]) ? node1799 : node1794;
										assign node1794 = (inp[0]) ? 3'b010 : node1795;
											assign node1795 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1799 = (inp[9]) ? 3'b010 : node1800;
											assign node1800 = (inp[0]) ? 3'b011 : 3'b010;
						assign node1804 = (inp[2]) ? node1828 : node1805;
							assign node1805 = (inp[9]) ? node1817 : node1806;
								assign node1806 = (inp[10]) ? node1812 : node1807;
									assign node1807 = (inp[11]) ? node1809 : 3'b010;
										assign node1809 = (inp[7]) ? 3'b011 : 3'b010;
									assign node1812 = (inp[7]) ? 3'b011 : node1813;
										assign node1813 = (inp[11]) ? 3'b010 : 3'b011;
								assign node1817 = (inp[10]) ? node1823 : node1818;
									assign node1818 = (inp[11]) ? node1820 : 3'b011;
										assign node1820 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1823 = (inp[11]) ? node1825 : 3'b010;
										assign node1825 = (inp[7]) ? 3'b010 : 3'b011;
							assign node1828 = (inp[11]) ? node1852 : node1829;
								assign node1829 = (inp[0]) ? node1843 : node1830;
									assign node1830 = (inp[7]) ? node1838 : node1831;
										assign node1831 = (inp[9]) ? node1835 : node1832;
											assign node1832 = (inp[10]) ? 3'b010 : 3'b011;
											assign node1835 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1838 = (inp[1]) ? node1840 : 3'b010;
											assign node1840 = (inp[10]) ? 3'b010 : 3'b010;
									assign node1843 = (inp[9]) ? node1847 : node1844;
										assign node1844 = (inp[7]) ? 3'b011 : 3'b010;
										assign node1847 = (inp[7]) ? node1849 : 3'b011;
											assign node1849 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1852 = (inp[7]) ? node1856 : node1853;
									assign node1853 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1856 = (inp[9]) ? 3'b010 : 3'b011;
					assign node1859 = (inp[8]) ? node1951 : node1860;
						assign node1860 = (inp[10]) ? node1904 : node1861;
							assign node1861 = (inp[11]) ? node1883 : node1862;
								assign node1862 = (inp[7]) ? node1874 : node1863;
									assign node1863 = (inp[0]) ? node1869 : node1864;
										assign node1864 = (inp[9]) ? node1866 : 3'b000;
											assign node1866 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1869 = (inp[2]) ? node1871 : 3'b000;
											assign node1871 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1874 = (inp[1]) ? node1878 : node1875;
										assign node1875 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1878 = (inp[9]) ? 3'b010 : node1879;
											assign node1879 = (inp[0]) ? 3'b010 : 3'b011;
								assign node1883 = (inp[1]) ? node1897 : node1884;
									assign node1884 = (inp[9]) ? node1892 : node1885;
										assign node1885 = (inp[0]) ? node1889 : node1886;
											assign node1886 = (inp[2]) ? 3'b010 : 3'b011;
											assign node1889 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1892 = (inp[0]) ? node1894 : 3'b011;
											assign node1894 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1897 = (inp[2]) ? node1899 : 3'b010;
										assign node1899 = (inp[9]) ? node1901 : 3'b011;
											assign node1901 = (inp[0]) ? 3'b010 : 3'b011;
							assign node1904 = (inp[11]) ? node1924 : node1905;
								assign node1905 = (inp[7]) ? node1913 : node1906;
									assign node1906 = (inp[9]) ? node1908 : 3'b011;
										assign node1908 = (inp[2]) ? node1910 : 3'b011;
											assign node1910 = (inp[0]) ? 3'b010 : 3'b010;
									assign node1913 = (inp[0]) ? node1919 : node1914;
										assign node1914 = (inp[9]) ? 3'b001 : node1915;
											assign node1915 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1919 = (inp[1]) ? 3'b000 : node1920;
											assign node1920 = (inp[9]) ? 3'b001 : 3'b000;
								assign node1924 = (inp[2]) ? node1940 : node1925;
									assign node1925 = (inp[1]) ? node1933 : node1926;
										assign node1926 = (inp[7]) ? node1930 : node1927;
											assign node1927 = (inp[9]) ? 3'b000 : 3'b000;
											assign node1930 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1933 = (inp[7]) ? node1937 : node1934;
											assign node1934 = (inp[9]) ? 3'b000 : 3'b000;
											assign node1937 = (inp[0]) ? 3'b000 : 3'b000;
									assign node1940 = (inp[1]) ? node1946 : node1941;
										assign node1941 = (inp[0]) ? node1943 : 3'b000;
											assign node1943 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1946 = (inp[0]) ? 3'b000 : node1947;
											assign node1947 = (inp[9]) ? 3'b001 : 3'b000;
						assign node1951 = (inp[9]) ? node1965 : node1952;
							assign node1952 = (inp[11]) ? 3'b001 : node1953;
								assign node1953 = (inp[10]) ? node1959 : node1954;
									assign node1954 = (inp[7]) ? 3'b000 : node1955;
										assign node1955 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1959 = (inp[7]) ? 3'b001 : node1960;
										assign node1960 = (inp[2]) ? 3'b001 : 3'b000;
							assign node1965 = (inp[11]) ? 3'b000 : node1966;
								assign node1966 = (inp[10]) ? node1972 : node1967;
									assign node1967 = (inp[7]) ? 3'b001 : node1968;
										assign node1968 = (inp[2]) ? 3'b001 : 3'b000;
									assign node1972 = (inp[7]) ? 3'b000 : node1973;
										assign node1973 = (inp[2]) ? 3'b000 : 3'b001;
			assign node1978 = (inp[8]) ? node2178 : node1979;
				assign node1979 = (inp[10]) ? node2107 : node1980;
					assign node1980 = (inp[6]) ? node2044 : node1981;
						assign node1981 = (inp[7]) ? node2005 : node1982;
							assign node1982 = (inp[0]) ? node1994 : node1983;
								assign node1983 = (inp[3]) ? node1989 : node1984;
									assign node1984 = (inp[11]) ? node1986 : 3'b000;
										assign node1986 = (inp[1]) ? 3'b001 : 3'b000;
									assign node1989 = (inp[1]) ? node1991 : 3'b001;
										assign node1991 = (inp[11]) ? 3'b000 : 3'b001;
								assign node1994 = (inp[3]) ? node2000 : node1995;
									assign node1995 = (inp[11]) ? node1997 : 3'b001;
										assign node1997 = (inp[1]) ? 3'b000 : 3'b001;
									assign node2000 = (inp[1]) ? node2002 : 3'b000;
										assign node2002 = (inp[11]) ? 3'b001 : 3'b000;
							assign node2005 = (inp[2]) ? node2025 : node2006;
								assign node2006 = (inp[9]) ? node2012 : node2007;
									assign node2007 = (inp[11]) ? 3'b011 : node2008;
										assign node2008 = (inp[0]) ? 3'b011 : 3'b010;
									assign node2012 = (inp[3]) ? node2018 : node2013;
										assign node2013 = (inp[1]) ? 3'b010 : node2014;
											assign node2014 = (inp[11]) ? 3'b010 : 3'b011;
										assign node2018 = (inp[0]) ? node2022 : node2019;
											assign node2019 = (inp[11]) ? 3'b011 : 3'b010;
											assign node2022 = (inp[11]) ? 3'b010 : 3'b011;
								assign node2025 = (inp[9]) ? node2037 : node2026;
									assign node2026 = (inp[3]) ? node2032 : node2027;
										assign node2027 = (inp[1]) ? node2029 : 3'b010;
											assign node2029 = (inp[11]) ? 3'b010 : 3'b010;
										assign node2032 = (inp[11]) ? node2034 : 3'b010;
											assign node2034 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2037 = (inp[11]) ? node2041 : node2038;
										assign node2038 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2041 = (inp[0]) ? 3'b010 : 3'b011;
						assign node2044 = (inp[7]) ? node2074 : node2045;
							assign node2045 = (inp[11]) ? node2059 : node2046;
								assign node2046 = (inp[3]) ? node2054 : node2047;
									assign node2047 = (inp[0]) ? node2051 : node2048;
										assign node2048 = (inp[1]) ? 3'b011 : 3'b010;
										assign node2051 = (inp[1]) ? 3'b010 : 3'b011;
									assign node2054 = (inp[0]) ? node2056 : 3'b011;
										assign node2056 = (inp[1]) ? 3'b011 : 3'b010;
								assign node2059 = (inp[9]) ? node2067 : node2060;
									assign node2060 = (inp[3]) ? node2064 : node2061;
										assign node2061 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2064 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2067 = (inp[0]) ? node2071 : node2068;
										assign node2068 = (inp[3]) ? 3'b011 : 3'b010;
										assign node2071 = (inp[3]) ? 3'b010 : 3'b011;
							assign node2074 = (inp[9]) ? node2082 : node2075;
								assign node2075 = (inp[11]) ? node2079 : node2076;
									assign node2076 = (inp[0]) ? 3'b011 : 3'b010;
									assign node2079 = (inp[0]) ? 3'b010 : 3'b011;
								assign node2082 = (inp[1]) ? node2092 : node2083;
									assign node2083 = (inp[3]) ? 3'b010 : node2084;
										assign node2084 = (inp[11]) ? node2088 : node2085;
											assign node2085 = (inp[0]) ? 3'b011 : 3'b010;
											assign node2088 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2092 = (inp[2]) ? node2100 : node2093;
										assign node2093 = (inp[0]) ? node2097 : node2094;
											assign node2094 = (inp[11]) ? 3'b011 : 3'b010;
											assign node2097 = (inp[11]) ? 3'b010 : 3'b011;
										assign node2100 = (inp[0]) ? node2104 : node2101;
											assign node2101 = (inp[11]) ? 3'b011 : 3'b010;
											assign node2104 = (inp[11]) ? 3'b010 : 3'b011;
					assign node2107 = (inp[6]) ? node2151 : node2108;
						assign node2108 = (inp[7]) ? node2144 : node2109;
							assign node2109 = (inp[1]) ? node2125 : node2110;
								assign node2110 = (inp[3]) ? node2118 : node2111;
									assign node2111 = (inp[0]) ? node2115 : node2112;
										assign node2112 = (inp[11]) ? 3'b011 : 3'b010;
										assign node2115 = (inp[11]) ? 3'b010 : 3'b011;
									assign node2118 = (inp[0]) ? node2122 : node2119;
										assign node2119 = (inp[11]) ? 3'b010 : 3'b011;
										assign node2122 = (inp[11]) ? 3'b011 : 3'b010;
								assign node2125 = (inp[2]) ? node2137 : node2126;
									assign node2126 = (inp[9]) ? node2132 : node2127;
										assign node2127 = (inp[11]) ? 3'b010 : node2128;
											assign node2128 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2132 = (inp[11]) ? node2134 : 3'b010;
											assign node2134 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2137 = (inp[0]) ? node2141 : node2138;
										assign node2138 = (inp[3]) ? 3'b011 : 3'b010;
										assign node2141 = (inp[3]) ? 3'b010 : 3'b011;
							assign node2144 = (inp[1]) ? node2148 : node2145;
								assign node2145 = (inp[0]) ? 3'b001 : 3'b000;
								assign node2148 = (inp[0]) ? 3'b000 : 3'b001;
						assign node2151 = (inp[0]) ? node2165 : node2152;
							assign node2152 = (inp[7]) ? 3'b001 : node2153;
								assign node2153 = (inp[3]) ? node2159 : node2154;
									assign node2154 = (inp[1]) ? 3'b000 : node2155;
										assign node2155 = (inp[11]) ? 3'b000 : 3'b001;
									assign node2159 = (inp[11]) ? 3'b001 : node2160;
										assign node2160 = (inp[1]) ? 3'b001 : 3'b000;
							assign node2165 = (inp[7]) ? 3'b000 : node2166;
								assign node2166 = (inp[3]) ? node2172 : node2167;
									assign node2167 = (inp[11]) ? 3'b001 : node2168;
										assign node2168 = (inp[1]) ? 3'b001 : 3'b000;
									assign node2172 = (inp[1]) ? 3'b000 : node2173;
										assign node2173 = (inp[11]) ? 3'b000 : 3'b001;
				assign node2178 = (inp[6]) ? node2198 : node2179;
					assign node2179 = (inp[7]) ? node2187 : node2180;
						assign node2180 = (inp[3]) ? node2184 : node2181;
							assign node2181 = (inp[1]) ? 3'b011 : 3'b010;
							assign node2184 = (inp[1]) ? 3'b010 : 3'b011;
						assign node2187 = (inp[1]) ? node2193 : node2188;
							assign node2188 = (inp[11]) ? 3'b001 : node2189;
								assign node2189 = (inp[10]) ? 3'b001 : 3'b000;
							assign node2193 = (inp[11]) ? 3'b000 : node2194;
								assign node2194 = (inp[10]) ? 3'b000 : 3'b001;
					assign node2198 = (inp[10]) ? node2210 : node2199;
						assign node2199 = (inp[11]) ? node2205 : node2200;
							assign node2200 = (inp[3]) ? 3'b001 : node2201;
								assign node2201 = (inp[7]) ? 3'b001 : 3'b000;
							assign node2205 = (inp[3]) ? 3'b000 : node2206;
								assign node2206 = (inp[7]) ? 3'b000 : 3'b001;
						assign node2210 = (inp[7]) ? 3'b000 : node2211;
							assign node2211 = (inp[3]) ? 3'b000 : 3'b001;

endmodule