module dtc_split25_bm72 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;

	assign outp = (inp[6]) ? node62 : node1;
		assign node1 = (inp[3]) ? node33 : node2;
			assign node2 = (inp[9]) ? node18 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[7]) ? node8 : node5;
						assign node5 = (inp[4]) ? 3'b010 : 3'b001;
						assign node8 = (inp[4]) ? 3'b101 : 3'b101;
					assign node11 = (inp[4]) ? node15 : node12;
						assign node12 = (inp[7]) ? 3'b001 : 3'b010;
						assign node15 = (inp[7]) ? 3'b010 : 3'b000;
				assign node18 = (inp[10]) ? node26 : node19;
					assign node19 = (inp[0]) ? node23 : node20;
						assign node20 = (inp[4]) ? 3'b010 : 3'b000;
						assign node23 = (inp[7]) ? 3'b010 : 3'b000;
					assign node26 = (inp[0]) ? node30 : node27;
						assign node27 = (inp[5]) ? 3'b000 : 3'b010;
						assign node30 = (inp[8]) ? 3'b000 : 3'b000;
			assign node33 = (inp[9]) ? node49 : node34;
				assign node34 = (inp[4]) ? node42 : node35;
					assign node35 = (inp[0]) ? node39 : node36;
						assign node36 = (inp[1]) ? 3'b110 : 3'b000;
						assign node39 = (inp[10]) ? 3'b000 : 3'b100;
					assign node42 = (inp[0]) ? node46 : node43;
						assign node43 = (inp[7]) ? 3'b100 : 3'b000;
						assign node46 = (inp[10]) ? 3'b000 : 3'b000;
				assign node49 = (inp[7]) ? node55 : node50;
					assign node50 = (inp[4]) ? 3'b000 : node51;
						assign node51 = (inp[5]) ? 3'b000 : 3'b000;
					assign node55 = (inp[0]) ? node59 : node56;
						assign node56 = (inp[11]) ? 3'b000 : 3'b100;
						assign node59 = (inp[4]) ? 3'b000 : 3'b000;
		assign node62 = (inp[3]) ? node94 : node63;
			assign node63 = (inp[9]) ? node79 : node64;
				assign node64 = (inp[0]) ? node72 : node65;
					assign node65 = (inp[4]) ? node69 : node66;
						assign node66 = (inp[7]) ? 3'b111 : 3'b111;
						assign node69 = (inp[11]) ? 3'b111 : 3'b111;
					assign node72 = (inp[7]) ? node76 : node73;
						assign node73 = (inp[4]) ? 3'b101 : 3'b001;
						assign node76 = (inp[4]) ? 3'b001 : 3'b111;
				assign node79 = (inp[0]) ? node87 : node80;
					assign node80 = (inp[4]) ? node84 : node81;
						assign node81 = (inp[7]) ? 3'b111 : 3'b001;
						assign node84 = (inp[5]) ? 3'b001 : 3'b101;
					assign node87 = (inp[4]) ? node91 : node88;
						assign node88 = (inp[7]) ? 3'b011 : 3'b100;
						assign node91 = (inp[11]) ? 3'b110 : 3'b010;
			assign node94 = (inp[9]) ? node110 : node95;
				assign node95 = (inp[0]) ? node103 : node96;
					assign node96 = (inp[4]) ? node100 : node97;
						assign node97 = (inp[2]) ? 3'b001 : 3'b101;
						assign node100 = (inp[1]) ? 3'b110 : 3'b001;
					assign node103 = (inp[10]) ? node107 : node104;
						assign node104 = (inp[7]) ? 3'b101 : 3'b110;
						assign node107 = (inp[1]) ? 3'b010 : 3'b010;
				assign node110 = (inp[0]) ? node118 : node111;
					assign node111 = (inp[7]) ? node115 : node112;
						assign node112 = (inp[4]) ? 3'b000 : 3'b110;
						assign node115 = (inp[4]) ? 3'b110 : 3'b101;
					assign node118 = (inp[4]) ? node122 : node119;
						assign node119 = (inp[10]) ? 3'b000 : 3'b110;
						assign node122 = (inp[7]) ? 3'b000 : 3'b000;

endmodule