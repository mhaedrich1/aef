module dtc_split33_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node604;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node740;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node818;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;

	assign outp = (inp[9]) ? node282 : node1;
		assign node1 = (inp[3]) ? node213 : node2;
			assign node2 = (inp[6]) ? node128 : node3;
				assign node3 = (inp[7]) ? node65 : node4;
					assign node4 = (inp[10]) ? node36 : node5;
						assign node5 = (inp[4]) ? node21 : node6;
							assign node6 = (inp[5]) ? node14 : node7;
								assign node7 = (inp[11]) ? node11 : node8;
									assign node8 = (inp[8]) ? 3'b001 : 3'b101;
									assign node11 = (inp[8]) ? 3'b101 : 3'b011;
								assign node14 = (inp[11]) ? node18 : node15;
									assign node15 = (inp[8]) ? 3'b110 : 3'b001;
									assign node18 = (inp[8]) ? 3'b001 : 3'b101;
							assign node21 = (inp[11]) ? node29 : node22;
								assign node22 = (inp[5]) ? node26 : node23;
									assign node23 = (inp[8]) ? 3'b010 : 3'b110;
									assign node26 = (inp[8]) ? 3'b100 : 3'b010;
								assign node29 = (inp[5]) ? node33 : node30;
									assign node30 = (inp[8]) ? 3'b110 : 3'b001;
									assign node33 = (inp[8]) ? 3'b010 : 3'b110;
						assign node36 = (inp[4]) ? node50 : node37;
							assign node37 = (inp[5]) ? node43 : node38;
								assign node38 = (inp[11]) ? 3'b111 : node39;
									assign node39 = (inp[8]) ? 3'b011 : 3'b111;
								assign node43 = (inp[8]) ? node47 : node44;
									assign node44 = (inp[11]) ? 3'b111 : 3'b011;
									assign node47 = (inp[11]) ? 3'b011 : 3'b101;
							assign node50 = (inp[5]) ? node58 : node51;
								assign node51 = (inp[11]) ? node55 : node52;
									assign node52 = (inp[8]) ? 3'b001 : 3'b101;
									assign node55 = (inp[8]) ? 3'b101 : 3'b011;
								assign node58 = (inp[8]) ? node62 : node59;
									assign node59 = (inp[11]) ? 3'b101 : 3'b001;
									assign node62 = (inp[1]) ? 3'b110 : 3'b001;
					assign node65 = (inp[10]) ? node93 : node66;
						assign node66 = (inp[4]) ? node82 : node67;
							assign node67 = (inp[5]) ? node75 : node68;
								assign node68 = (inp[8]) ? node72 : node69;
									assign node69 = (inp[11]) ? 3'b001 : 3'b110;
									assign node72 = (inp[11]) ? 3'b110 : 3'b010;
								assign node75 = (inp[11]) ? node79 : node76;
									assign node76 = (inp[8]) ? 3'b100 : 3'b010;
									assign node79 = (inp[8]) ? 3'b010 : 3'b110;
							assign node82 = (inp[11]) ? node88 : node83;
								assign node83 = (inp[8]) ? 3'b000 : node84;
									assign node84 = (inp[5]) ? 3'b000 : 3'b100;
								assign node88 = (inp[1]) ? node90 : 3'b100;
									assign node90 = (inp[8]) ? 3'b000 : 3'b100;
						assign node93 = (inp[4]) ? node111 : node94;
							assign node94 = (inp[5]) ? node102 : node95;
								assign node95 = (inp[8]) ? node99 : node96;
									assign node96 = (inp[11]) ? 3'b011 : 3'b101;
									assign node99 = (inp[11]) ? 3'b101 : 3'b001;
								assign node102 = (inp[1]) ? 3'b001 : node103;
									assign node103 = (inp[8]) ? node107 : node104;
										assign node104 = (inp[11]) ? 3'b101 : 3'b001;
										assign node107 = (inp[11]) ? 3'b001 : 3'b110;
							assign node111 = (inp[8]) ? node119 : node112;
								assign node112 = (inp[11]) ? node116 : node113;
									assign node113 = (inp[5]) ? 3'b010 : 3'b110;
									assign node116 = (inp[5]) ? 3'b110 : 3'b001;
								assign node119 = (inp[2]) ? 3'b010 : node120;
									assign node120 = (inp[5]) ? node124 : node121;
										assign node121 = (inp[11]) ? 3'b110 : 3'b010;
										assign node124 = (inp[11]) ? 3'b010 : 3'b100;
				assign node128 = (inp[10]) ? node146 : node129;
					assign node129 = (inp[7]) ? 3'b000 : node130;
						assign node130 = (inp[4]) ? 3'b000 : node131;
							assign node131 = (inp[5]) ? node139 : node132;
								assign node132 = (inp[8]) ? node136 : node133;
									assign node133 = (inp[11]) ? 3'b010 : 3'b100;
									assign node136 = (inp[11]) ? 3'b100 : 3'b000;
								assign node139 = (inp[8]) ? 3'b000 : node140;
									assign node140 = (inp[11]) ? 3'b100 : 3'b000;
					assign node146 = (inp[4]) ? node190 : node147;
						assign node147 = (inp[7]) ? node173 : node148;
							assign node148 = (inp[1]) ? node158 : node149;
								assign node149 = (inp[5]) ? node153 : node150;
									assign node150 = (inp[11]) ? 3'b001 : 3'b010;
									assign node153 = (inp[2]) ? node155 : 3'b010;
										assign node155 = (inp[11]) ? 3'b110 : 3'b010;
								assign node158 = (inp[0]) ? node168 : node159;
									assign node159 = (inp[2]) ? node163 : node160;
										assign node160 = (inp[5]) ? 3'b010 : 3'b110;
										assign node163 = (inp[5]) ? node165 : 3'b110;
											assign node165 = (inp[11]) ? 3'b110 : 3'b100;
									assign node168 = (inp[8]) ? 3'b110 : node169;
										assign node169 = (inp[5]) ? 3'b110 : 3'b001;
							assign node173 = (inp[2]) ? node185 : node174;
								assign node174 = (inp[11]) ? node180 : node175;
									assign node175 = (inp[5]) ? 3'b000 : node176;
										assign node176 = (inp[1]) ? 3'b100 : 3'b000;
									assign node180 = (inp[0]) ? node182 : 3'b010;
										assign node182 = (inp[1]) ? 3'b000 : 3'b100;
								assign node185 = (inp[11]) ? 3'b100 : node186;
									assign node186 = (inp[8]) ? 3'b000 : 3'b100;
						assign node190 = (inp[7]) ? node204 : node191;
							assign node191 = (inp[5]) ? node199 : node192;
								assign node192 = (inp[8]) ? node196 : node193;
									assign node193 = (inp[11]) ? 3'b010 : 3'b100;
									assign node196 = (inp[11]) ? 3'b100 : 3'b000;
								assign node199 = (inp[11]) ? node201 : 3'b000;
									assign node201 = (inp[8]) ? 3'b000 : 3'b100;
							assign node204 = (inp[11]) ? node206 : 3'b000;
								assign node206 = (inp[5]) ? 3'b000 : node207;
									assign node207 = (inp[0]) ? 3'b000 : node208;
										assign node208 = (inp[8]) ? 3'b000 : 3'b100;
			assign node213 = (inp[6]) ? 3'b000 : node214;
				assign node214 = (inp[10]) ? node236 : node215;
					assign node215 = (inp[7]) ? 3'b000 : node216;
						assign node216 = (inp[4]) ? 3'b000 : node217;
							assign node217 = (inp[8]) ? node229 : node218;
								assign node218 = (inp[0]) ? node224 : node219;
									assign node219 = (inp[11]) ? 3'b100 : node220;
										assign node220 = (inp[2]) ? 3'b000 : 3'b100;
									assign node224 = (inp[5]) ? node226 : 3'b010;
										assign node226 = (inp[11]) ? 3'b100 : 3'b000;
								assign node229 = (inp[5]) ? 3'b000 : node230;
									assign node230 = (inp[11]) ? 3'b100 : 3'b000;
					assign node236 = (inp[4]) ? node270 : node237;
						assign node237 = (inp[7]) ? node257 : node238;
							assign node238 = (inp[2]) ? node246 : node239;
								assign node239 = (inp[0]) ? node241 : 3'b110;
									assign node241 = (inp[11]) ? node243 : 3'b010;
										assign node243 = (inp[1]) ? 3'b110 : 3'b010;
								assign node246 = (inp[11]) ? node254 : node247;
									assign node247 = (inp[8]) ? node251 : node248;
										assign node248 = (inp[5]) ? 3'b010 : 3'b110;
										assign node251 = (inp[5]) ? 3'b100 : 3'b010;
									assign node254 = (inp[5]) ? 3'b110 : 3'b001;
							assign node257 = (inp[11]) ? node263 : node258;
								assign node258 = (inp[5]) ? 3'b000 : node259;
									assign node259 = (inp[8]) ? 3'b000 : 3'b100;
								assign node263 = (inp[5]) ? node267 : node264;
									assign node264 = (inp[8]) ? 3'b100 : 3'b010;
									assign node267 = (inp[8]) ? 3'b000 : 3'b100;
						assign node270 = (inp[11]) ? node272 : 3'b000;
							assign node272 = (inp[7]) ? 3'b000 : node273;
								assign node273 = (inp[1]) ? node275 : 3'b000;
									assign node275 = (inp[5]) ? 3'b100 : node276;
										assign node276 = (inp[8]) ? 3'b100 : 3'b010;
		assign node282 = (inp[6]) ? node540 : node283;
			assign node283 = (inp[3]) ? node357 : node284;
				assign node284 = (inp[7]) ? node306 : node285;
					assign node285 = (inp[10]) ? 3'b111 : node286;
						assign node286 = (inp[4]) ? node288 : 3'b111;
							assign node288 = (inp[11]) ? node296 : node289;
								assign node289 = (inp[5]) ? node293 : node290;
									assign node290 = (inp[8]) ? 3'b011 : 3'b111;
									assign node293 = (inp[8]) ? 3'b101 : 3'b011;
								assign node296 = (inp[8]) ? node298 : 3'b111;
									assign node298 = (inp[5]) ? node300 : 3'b111;
										assign node300 = (inp[1]) ? 3'b011 : node301;
											assign node301 = (inp[0]) ? 3'b011 : 3'b111;
					assign node306 = (inp[10]) ? node338 : node307;
						assign node307 = (inp[4]) ? node321 : node308;
							assign node308 = (inp[5]) ? node314 : node309;
								assign node309 = (inp[8]) ? node311 : 3'b111;
									assign node311 = (inp[11]) ? 3'b111 : 3'b011;
								assign node314 = (inp[11]) ? node318 : node315;
									assign node315 = (inp[8]) ? 3'b101 : 3'b011;
									assign node318 = (inp[8]) ? 3'b011 : 3'b111;
							assign node321 = (inp[11]) ? node329 : node322;
								assign node322 = (inp[8]) ? node326 : node323;
									assign node323 = (inp[5]) ? 3'b001 : 3'b101;
									assign node326 = (inp[5]) ? 3'b110 : 3'b001;
								assign node329 = (inp[5]) ? node335 : node330;
									assign node330 = (inp[8]) ? node332 : 3'b011;
										assign node332 = (inp[2]) ? 3'b101 : 3'b011;
									assign node335 = (inp[8]) ? 3'b001 : 3'b101;
						assign node338 = (inp[4]) ? node340 : 3'b111;
							assign node340 = (inp[8]) ? node342 : 3'b111;
								assign node342 = (inp[11]) ? node352 : node343;
									assign node343 = (inp[5]) ? node349 : node344;
										assign node344 = (inp[0]) ? 3'b011 : node345;
											assign node345 = (inp[1]) ? 3'b011 : 3'b111;
										assign node349 = (inp[2]) ? 3'b101 : 3'b011;
									assign node352 = (inp[0]) ? node354 : 3'b111;
										assign node354 = (inp[2]) ? 3'b011 : 3'b111;
				assign node357 = (inp[10]) ? node443 : node358;
					assign node358 = (inp[7]) ? node396 : node359;
						assign node359 = (inp[4]) ? node377 : node360;
							assign node360 = (inp[5]) ? node366 : node361;
								assign node361 = (inp[11]) ? 3'b011 : node362;
									assign node362 = (inp[8]) ? 3'b001 : 3'b101;
								assign node366 = (inp[11]) ? node370 : node367;
									assign node367 = (inp[2]) ? 3'b110 : 3'b001;
									assign node370 = (inp[8]) ? node372 : 3'b101;
										assign node372 = (inp[2]) ? 3'b001 : node373;
											assign node373 = (inp[1]) ? 3'b001 : 3'b101;
							assign node377 = (inp[5]) ? node387 : node378;
								assign node378 = (inp[11]) ? node382 : node379;
									assign node379 = (inp[8]) ? 3'b010 : 3'b110;
									assign node382 = (inp[8]) ? node384 : 3'b001;
										assign node384 = (inp[0]) ? 3'b110 : 3'b001;
								assign node387 = (inp[11]) ? node391 : node388;
									assign node388 = (inp[8]) ? 3'b100 : 3'b010;
									assign node391 = (inp[0]) ? node393 : 3'b110;
										assign node393 = (inp[8]) ? 3'b010 : 3'b110;
						assign node396 = (inp[4]) ? node424 : node397;
							assign node397 = (inp[5]) ? node409 : node398;
								assign node398 = (inp[11]) ? node404 : node399;
									assign node399 = (inp[8]) ? node401 : 3'b110;
										assign node401 = (inp[0]) ? 3'b010 : 3'b110;
									assign node404 = (inp[2]) ? node406 : 3'b001;
										assign node406 = (inp[0]) ? 3'b110 : 3'b101;
								assign node409 = (inp[8]) ? node417 : node410;
									assign node410 = (inp[11]) ? 3'b110 : node411;
										assign node411 = (inp[2]) ? 3'b010 : node412;
											assign node412 = (inp[1]) ? 3'b010 : 3'b110;
									assign node417 = (inp[11]) ? node419 : 3'b100;
										assign node419 = (inp[0]) ? 3'b010 : node420;
											assign node420 = (inp[2]) ? 3'b010 : 3'b110;
							assign node424 = (inp[11]) ? node436 : node425;
								assign node425 = (inp[8]) ? node431 : node426;
									assign node426 = (inp[5]) ? node428 : 3'b100;
										assign node428 = (inp[0]) ? 3'b000 : 3'b100;
									assign node431 = (inp[1]) ? 3'b000 : node432;
										assign node432 = (inp[0]) ? 3'b000 : 3'b100;
								assign node436 = (inp[8]) ? node438 : 3'b010;
									assign node438 = (inp[5]) ? node440 : 3'b100;
										assign node440 = (inp[1]) ? 3'b000 : 3'b100;
					assign node443 = (inp[4]) ? node491 : node444;
						assign node444 = (inp[7]) ? node464 : node445;
							assign node445 = (inp[11]) ? node459 : node446;
								assign node446 = (inp[8]) ? node452 : node447;
									assign node447 = (inp[5]) ? node449 : 3'b111;
										assign node449 = (inp[2]) ? 3'b111 : 3'b011;
									assign node452 = (inp[5]) ? node454 : 3'b011;
										assign node454 = (inp[1]) ? node456 : 3'b101;
											assign node456 = (inp[2]) ? 3'b101 : 3'b011;
								assign node459 = (inp[0]) ? node461 : 3'b111;
									assign node461 = (inp[5]) ? 3'b011 : 3'b111;
							assign node464 = (inp[2]) ? node478 : node465;
								assign node465 = (inp[5]) ? node473 : node466;
									assign node466 = (inp[1]) ? node468 : 3'b011;
										assign node468 = (inp[11]) ? node470 : 3'b011;
											assign node470 = (inp[0]) ? 3'b011 : 3'b111;
									assign node473 = (inp[11]) ? node475 : 3'b110;
										assign node475 = (inp[0]) ? 3'b101 : 3'b011;
								assign node478 = (inp[1]) ? node484 : node479;
									assign node479 = (inp[0]) ? 3'b110 : node480;
										assign node480 = (inp[5]) ? 3'b001 : 3'b111;
									assign node484 = (inp[11]) ? node486 : 3'b101;
										assign node486 = (inp[8]) ? 3'b101 : node487;
											assign node487 = (inp[5]) ? 3'b101 : 3'b011;
						assign node491 = (inp[7]) ? node519 : node492;
							assign node492 = (inp[0]) ? node510 : node493;
								assign node493 = (inp[11]) ? node503 : node494;
									assign node494 = (inp[1]) ? node496 : 3'b011;
										assign node496 = (inp[5]) ? node500 : node497;
											assign node497 = (inp[8]) ? 3'b001 : 3'b101;
											assign node500 = (inp[8]) ? 3'b110 : 3'b101;
									assign node503 = (inp[2]) ? node507 : node504;
										assign node504 = (inp[8]) ? 3'b011 : 3'b111;
										assign node507 = (inp[8]) ? 3'b101 : 3'b011;
								assign node510 = (inp[8]) ? node516 : node511;
									assign node511 = (inp[11]) ? 3'b101 : node512;
										assign node512 = (inp[5]) ? 3'b001 : 3'b101;
									assign node516 = (inp[5]) ? 3'b110 : 3'b001;
							assign node519 = (inp[0]) ? node533 : node520;
								assign node520 = (inp[2]) ? node524 : node521;
									assign node521 = (inp[8]) ? 3'b110 : 3'b101;
									assign node524 = (inp[5]) ? node530 : node525;
										assign node525 = (inp[1]) ? node527 : 3'b001;
											assign node527 = (inp[8]) ? 3'b001 : 3'b101;
										assign node530 = (inp[8]) ? 3'b110 : 3'b001;
								assign node533 = (inp[11]) ? 3'b110 : node534;
									assign node534 = (inp[5]) ? 3'b010 : node535;
										assign node535 = (inp[8]) ? 3'b010 : 3'b110;
			assign node540 = (inp[3]) ? node772 : node541;
				assign node541 = (inp[10]) ? node659 : node542;
					assign node542 = (inp[7]) ? node590 : node543;
						assign node543 = (inp[4]) ? node563 : node544;
							assign node544 = (inp[0]) ? node560 : node545;
								assign node545 = (inp[8]) ? node553 : node546;
									assign node546 = (inp[11]) ? node550 : node547;
										assign node547 = (inp[1]) ? 3'b001 : 3'b101;
										assign node550 = (inp[1]) ? 3'b101 : 3'b011;
									assign node553 = (inp[11]) ? node555 : 3'b110;
										assign node555 = (inp[5]) ? 3'b101 : node556;
											assign node556 = (inp[1]) ? 3'b101 : 3'b011;
								assign node560 = (inp[8]) ? 3'b001 : 3'b101;
							assign node563 = (inp[0]) ? node577 : node564;
								assign node564 = (inp[1]) ? node570 : node565;
									assign node565 = (inp[2]) ? 3'b001 : node566;
										assign node566 = (inp[11]) ? 3'b101 : 3'b001;
									assign node570 = (inp[11]) ? node574 : node571;
										assign node571 = (inp[5]) ? 3'b010 : 3'b110;
										assign node574 = (inp[5]) ? 3'b010 : 3'b001;
								assign node577 = (inp[5]) ? node585 : node578;
									assign node578 = (inp[1]) ? 3'b110 : node579;
										assign node579 = (inp[8]) ? node581 : 3'b001;
											assign node581 = (inp[2]) ? 3'b110 : 3'b010;
									assign node585 = (inp[8]) ? 3'b010 : node586;
										assign node586 = (inp[11]) ? 3'b110 : 3'b010;
						assign node590 = (inp[4]) ? node624 : node591;
							assign node591 = (inp[0]) ? node609 : node592;
								assign node592 = (inp[5]) ? node598 : node593;
									assign node593 = (inp[8]) ? 3'b001 : node594;
										assign node594 = (inp[11]) ? 3'b101 : 3'b001;
									assign node598 = (inp[1]) ? node604 : node599;
										assign node599 = (inp[11]) ? 3'b110 : node600;
											assign node600 = (inp[2]) ? 3'b110 : 3'b010;
										assign node604 = (inp[8]) ? node606 : 3'b001;
											assign node606 = (inp[2]) ? 3'b100 : 3'b110;
								assign node609 = (inp[11]) ? node619 : node610;
									assign node610 = (inp[2]) ? node612 : 3'b010;
										assign node612 = (inp[8]) ? node616 : node613;
											assign node613 = (inp[5]) ? 3'b010 : 3'b110;
											assign node616 = (inp[5]) ? 3'b100 : 3'b010;
									assign node619 = (inp[5]) ? node621 : 3'b110;
										assign node621 = (inp[8]) ? 3'b010 : 3'b110;
							assign node624 = (inp[8]) ? node648 : node625;
								assign node625 = (inp[5]) ? node639 : node626;
									assign node626 = (inp[2]) ? node632 : node627;
										assign node627 = (inp[1]) ? node629 : 3'b010;
											assign node629 = (inp[11]) ? 3'b010 : 3'b100;
										assign node632 = (inp[11]) ? node634 : 3'b010;
											assign node634 = (inp[0]) ? 3'b010 : node635;
												assign node635 = (inp[1]) ? 3'b010 : 3'b110;
									assign node639 = (inp[0]) ? node645 : node640;
										assign node640 = (inp[11]) ? 3'b010 : node641;
											assign node641 = (inp[1]) ? 3'b000 : 3'b100;
										assign node645 = (inp[11]) ? 3'b100 : 3'b000;
								assign node648 = (inp[0]) ? node654 : node649;
									assign node649 = (inp[5]) ? 3'b100 : node650;
										assign node650 = (inp[1]) ? 3'b000 : 3'b100;
									assign node654 = (inp[1]) ? node656 : 3'b000;
										assign node656 = (inp[11]) ? 3'b100 : 3'b000;
					assign node659 = (inp[11]) ? node723 : node660;
						assign node660 = (inp[7]) ? node684 : node661;
							assign node661 = (inp[4]) ? node667 : node662;
								assign node662 = (inp[8]) ? node664 : 3'b111;
									assign node664 = (inp[2]) ? 3'b011 : 3'b111;
								assign node667 = (inp[0]) ? node679 : node668;
									assign node668 = (inp[2]) ? node674 : node669;
										assign node669 = (inp[5]) ? 3'b101 : node670;
											assign node670 = (inp[8]) ? 3'b101 : 3'b011;
										assign node674 = (inp[8]) ? node676 : 3'b101;
											assign node676 = (inp[5]) ? 3'b001 : 3'b101;
									assign node679 = (inp[8]) ? 3'b110 : node680;
										assign node680 = (inp[5]) ? 3'b001 : 3'b101;
							assign node684 = (inp[4]) ? node698 : node685;
								assign node685 = (inp[1]) ? node691 : node686;
									assign node686 = (inp[5]) ? node688 : 3'b101;
										assign node688 = (inp[8]) ? 3'b001 : 3'b101;
									assign node691 = (inp[5]) ? node695 : node692;
										assign node692 = (inp[8]) ? 3'b001 : 3'b011;
										assign node695 = (inp[8]) ? 3'b110 : 3'b101;
								assign node698 = (inp[1]) ? node708 : node699;
									assign node699 = (inp[2]) ? node701 : 3'b110;
										assign node701 = (inp[8]) ? 3'b010 : node702;
											assign node702 = (inp[0]) ? node704 : 3'b110;
												assign node704 = (inp[5]) ? 3'b010 : 3'b110;
									assign node708 = (inp[0]) ? node716 : node709;
										assign node709 = (inp[8]) ? node713 : node710;
											assign node710 = (inp[5]) ? 3'b110 : 3'b001;
											assign node713 = (inp[2]) ? 3'b110 : 3'b010;
										assign node716 = (inp[2]) ? 3'b010 : node717;
											assign node717 = (inp[8]) ? 3'b100 : node718;
												assign node718 = (inp[5]) ? 3'b010 : 3'b110;
						assign node723 = (inp[7]) ? node745 : node724;
							assign node724 = (inp[4]) ? node730 : node725;
								assign node725 = (inp[0]) ? node727 : 3'b111;
									assign node727 = (inp[5]) ? 3'b011 : 3'b111;
								assign node730 = (inp[0]) ? node738 : node731;
									assign node731 = (inp[5]) ? node735 : node732;
										assign node732 = (inp[8]) ? 3'b011 : 3'b111;
										assign node735 = (inp[8]) ? 3'b101 : 3'b011;
									assign node738 = (inp[8]) ? node740 : 3'b101;
										assign node740 = (inp[1]) ? node742 : 3'b011;
											assign node742 = (inp[5]) ? 3'b001 : 3'b101;
							assign node745 = (inp[4]) ? node761 : node746;
								assign node746 = (inp[0]) ? node754 : node747;
									assign node747 = (inp[5]) ? node751 : node748;
										assign node748 = (inp[8]) ? 3'b011 : 3'b111;
										assign node751 = (inp[8]) ? 3'b101 : 3'b011;
									assign node754 = (inp[1]) ? node756 : 3'b101;
										assign node756 = (inp[8]) ? node758 : 3'b101;
											assign node758 = (inp[5]) ? 3'b001 : 3'b101;
								assign node761 = (inp[5]) ? node767 : node762;
									assign node762 = (inp[8]) ? 3'b001 : node763;
										assign node763 = (inp[1]) ? 3'b001 : 3'b101;
									assign node767 = (inp[1]) ? node769 : 3'b001;
										assign node769 = (inp[2]) ? 3'b010 : 3'b110;
				assign node772 = (inp[10]) ? node812 : node773;
					assign node773 = (inp[11]) ? node785 : node774;
						assign node774 = (inp[8]) ? 3'b000 : node775;
							assign node775 = (inp[0]) ? 3'b000 : node776;
								assign node776 = (inp[5]) ? node780 : node777;
									assign node777 = (inp[7]) ? 3'b000 : 3'b010;
									assign node780 = (inp[4]) ? 3'b000 : 3'b100;
						assign node785 = (inp[4]) ? node805 : node786;
							assign node786 = (inp[7]) ? node800 : node787;
								assign node787 = (inp[8]) ? node793 : node788;
									assign node788 = (inp[1]) ? node790 : 3'b010;
										assign node790 = (inp[5]) ? 3'b100 : 3'b010;
									assign node793 = (inp[2]) ? 3'b100 : node794;
										assign node794 = (inp[1]) ? 3'b010 : node795;
											assign node795 = (inp[0]) ? 3'b000 : 3'b100;
								assign node800 = (inp[0]) ? 3'b000 : node801;
									assign node801 = (inp[8]) ? 3'b000 : 3'b100;
							assign node805 = (inp[8]) ? 3'b000 : node806;
								assign node806 = (inp[0]) ? 3'b000 : node807;
									assign node807 = (inp[2]) ? 3'b000 : 3'b100;
					assign node812 = (inp[4]) ? node864 : node813;
						assign node813 = (inp[7]) ? node841 : node814;
							assign node814 = (inp[8]) ? node826 : node815;
								assign node815 = (inp[0]) ? node823 : node816;
									assign node816 = (inp[1]) ? node818 : 3'b001;
										assign node818 = (inp[11]) ? node820 : 3'b001;
											assign node820 = (inp[5]) ? 3'b001 : 3'b101;
									assign node823 = (inp[2]) ? 3'b001 : 3'b110;
								assign node826 = (inp[1]) ? node834 : node827;
									assign node827 = (inp[5]) ? node831 : node828;
										assign node828 = (inp[11]) ? 3'b001 : 3'b010;
										assign node831 = (inp[11]) ? 3'b110 : 3'b100;
									assign node834 = (inp[5]) ? node836 : 3'b110;
										assign node836 = (inp[0]) ? 3'b010 : node837;
											assign node837 = (inp[2]) ? 3'b010 : 3'b110;
							assign node841 = (inp[11]) ? node857 : node842;
								assign node842 = (inp[8]) ? node852 : node843;
									assign node843 = (inp[5]) ? node847 : node844;
										assign node844 = (inp[0]) ? 3'b100 : 3'b010;
										assign node847 = (inp[2]) ? node849 : 3'b100;
											assign node849 = (inp[1]) ? 3'b000 : 3'b100;
									assign node852 = (inp[5]) ? 3'b000 : node853;
										assign node853 = (inp[1]) ? 3'b000 : 3'b100;
								assign node857 = (inp[5]) ? node861 : node858;
									assign node858 = (inp[8]) ? 3'b010 : 3'b110;
									assign node861 = (inp[8]) ? 3'b100 : 3'b010;
						assign node864 = (inp[11]) ? node872 : node865;
							assign node865 = (inp[7]) ? 3'b000 : node866;
								assign node866 = (inp[8]) ? 3'b000 : node867;
									assign node867 = (inp[0]) ? 3'b000 : 3'b100;
							assign node872 = (inp[7]) ? node882 : node873;
								assign node873 = (inp[8]) ? node877 : node874;
									assign node874 = (inp[5]) ? 3'b010 : 3'b110;
									assign node877 = (inp[5]) ? 3'b100 : node878;
										assign node878 = (inp[0]) ? 3'b100 : 3'b010;
								assign node882 = (inp[5]) ? 3'b000 : node883;
									assign node883 = (inp[8]) ? 3'b000 : node884;
										assign node884 = (inp[0]) ? 3'b000 : 3'b100;

endmodule