module dtc_split66_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node580;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node798;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node938;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node956;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node963;

	assign outp = (inp[3]) ? node756 : node1;
		assign node1 = (inp[4]) ? node493 : node2;
			assign node2 = (inp[0]) ? node350 : node3;
				assign node3 = (inp[6]) ? node207 : node4;
					assign node4 = (inp[9]) ? node96 : node5;
						assign node5 = (inp[1]) ? node47 : node6;
							assign node6 = (inp[5]) ? node28 : node7;
								assign node7 = (inp[7]) ? node19 : node8;
									assign node8 = (inp[11]) ? node14 : node9;
										assign node9 = (inp[8]) ? node11 : 3'b000;
											assign node11 = (inp[10]) ? 3'b000 : 3'b000;
										assign node14 = (inp[8]) ? 3'b000 : node15;
											assign node15 = (inp[10]) ? 3'b000 : 3'b000;
									assign node19 = (inp[11]) ? node21 : 3'b100;
										assign node21 = (inp[8]) ? node25 : node22;
											assign node22 = (inp[2]) ? 3'b010 : 3'b000;
											assign node25 = (inp[10]) ? 3'b010 : 3'b010;
								assign node28 = (inp[2]) ? node36 : node29;
									assign node29 = (inp[10]) ? node31 : 3'b000;
										assign node31 = (inp[7]) ? 3'b000 : node32;
											assign node32 = (inp[11]) ? 3'b100 : 3'b000;
									assign node36 = (inp[10]) ? node42 : node37;
										assign node37 = (inp[7]) ? node39 : 3'b100;
											assign node39 = (inp[11]) ? 3'b100 : 3'b000;
										assign node42 = (inp[7]) ? node44 : 3'b000;
											assign node44 = (inp[11]) ? 3'b100 : 3'b000;
							assign node47 = (inp[2]) ? node71 : node48;
								assign node48 = (inp[10]) ? node62 : node49;
									assign node49 = (inp[11]) ? node55 : node50;
										assign node50 = (inp[5]) ? 3'b000 : node51;
											assign node51 = (inp[7]) ? 3'b010 : 3'b000;
										assign node55 = (inp[5]) ? node59 : node56;
											assign node56 = (inp[8]) ? 3'b000 : 3'b000;
											assign node59 = (inp[7]) ? 3'b100 : 3'b000;
									assign node62 = (inp[7]) ? node68 : node63;
										assign node63 = (inp[5]) ? 3'b100 : node64;
											assign node64 = (inp[11]) ? 3'b010 : 3'b010;
										assign node68 = (inp[5]) ? 3'b010 : 3'b011;
								assign node71 = (inp[8]) ? node85 : node72;
									assign node72 = (inp[11]) ? node80 : node73;
										assign node73 = (inp[10]) ? node77 : node74;
											assign node74 = (inp[7]) ? 3'b110 : 3'b010;
											assign node77 = (inp[7]) ? 3'b100 : 3'b110;
										assign node80 = (inp[7]) ? node82 : 3'b010;
											assign node82 = (inp[10]) ? 3'b110 : 3'b010;
									assign node85 = (inp[5]) ? node91 : node86;
										assign node86 = (inp[7]) ? 3'b101 : node87;
											assign node87 = (inp[11]) ? 3'b001 : 3'b010;
										assign node91 = (inp[10]) ? node93 : 3'b100;
											assign node93 = (inp[7]) ? 3'b110 : 3'b010;
						assign node96 = (inp[1]) ? node154 : node97;
							assign node97 = (inp[5]) ? node127 : node98;
								assign node98 = (inp[2]) ? node114 : node99;
									assign node99 = (inp[7]) ? node107 : node100;
										assign node100 = (inp[11]) ? node104 : node101;
											assign node101 = (inp[8]) ? 3'b010 : 3'b010;
											assign node104 = (inp[8]) ? 3'b010 : 3'b110;
										assign node107 = (inp[8]) ? node111 : node108;
											assign node108 = (inp[10]) ? 3'b110 : 3'b010;
											assign node111 = (inp[11]) ? 3'b000 : 3'b010;
									assign node114 = (inp[10]) ? node122 : node115;
										assign node115 = (inp[11]) ? node119 : node116;
											assign node116 = (inp[7]) ? 3'b110 : 3'b010;
											assign node119 = (inp[7]) ? 3'b110 : 3'b110;
										assign node122 = (inp[7]) ? 3'b101 : node123;
											assign node123 = (inp[8]) ? 3'b001 : 3'b110;
								assign node127 = (inp[10]) ? node141 : node128;
									assign node128 = (inp[11]) ? node134 : node129;
										assign node129 = (inp[8]) ? 3'b100 : node130;
											assign node130 = (inp[7]) ? 3'b000 : 3'b000;
										assign node134 = (inp[2]) ? node138 : node135;
											assign node135 = (inp[7]) ? 3'b100 : 3'b000;
											assign node138 = (inp[7]) ? 3'b010 : 3'b100;
									assign node141 = (inp[7]) ? node149 : node142;
										assign node142 = (inp[2]) ? node146 : node143;
											assign node143 = (inp[8]) ? 3'b100 : 3'b000;
											assign node146 = (inp[11]) ? 3'b010 : 3'b000;
										assign node149 = (inp[2]) ? node151 : 3'b010;
											assign node151 = (inp[11]) ? 3'b110 : 3'b000;
							assign node154 = (inp[5]) ? node182 : node155;
								assign node155 = (inp[7]) ? node169 : node156;
									assign node156 = (inp[10]) ? node162 : node157;
										assign node157 = (inp[2]) ? 3'b101 : node158;
											assign node158 = (inp[8]) ? 3'b000 : 3'b110;
										assign node162 = (inp[2]) ? node166 : node163;
											assign node163 = (inp[8]) ? 3'b101 : 3'b001;
											assign node166 = (inp[8]) ? 3'b011 : 3'b101;
									assign node169 = (inp[2]) ? node177 : node170;
										assign node170 = (inp[8]) ? node174 : node171;
											assign node171 = (inp[10]) ? 3'b101 : 3'b001;
											assign node174 = (inp[10]) ? 3'b011 : 3'b101;
										assign node177 = (inp[8]) ? 3'b011 : node178;
											assign node178 = (inp[11]) ? 3'b011 : 3'b001;
								assign node182 = (inp[10]) ? node196 : node183;
									assign node183 = (inp[2]) ? node189 : node184;
										assign node184 = (inp[7]) ? node186 : 3'b010;
											assign node186 = (inp[11]) ? 3'b110 : 3'b010;
										assign node189 = (inp[7]) ? node193 : node190;
											assign node190 = (inp[8]) ? 3'b110 : 3'b010;
											assign node193 = (inp[11]) ? 3'b001 : 3'b100;
									assign node196 = (inp[2]) ? node202 : node197;
										assign node197 = (inp[7]) ? node199 : 3'b110;
											assign node199 = (inp[11]) ? 3'b001 : 3'b100;
										assign node202 = (inp[7]) ? 3'b101 : node203;
											assign node203 = (inp[8]) ? 3'b001 : 3'b001;
					assign node207 = (inp[9]) ? node259 : node208;
						assign node208 = (inp[1]) ? node250 : node209;
							assign node209 = (inp[5]) ? node229 : node210;
								assign node210 = (inp[7]) ? node222 : node211;
									assign node211 = (inp[2]) ? node217 : node212;
										assign node212 = (inp[11]) ? 3'b010 : node213;
											assign node213 = (inp[10]) ? 3'b010 : 3'b011;
										assign node217 = (inp[8]) ? 3'b011 : node218;
											assign node218 = (inp[11]) ? 3'b011 : 3'b010;
									assign node222 = (inp[8]) ? 3'b011 : node223;
										assign node223 = (inp[2]) ? 3'b011 : node224;
											assign node224 = (inp[10]) ? 3'b011 : 3'b010;
								assign node229 = (inp[10]) ? node243 : node230;
									assign node230 = (inp[7]) ? node238 : node231;
										assign node231 = (inp[11]) ? node235 : node232;
											assign node232 = (inp[2]) ? 3'b011 : 3'b010;
											assign node235 = (inp[8]) ? 3'b010 : 3'b010;
										assign node238 = (inp[2]) ? 3'b010 : node239;
											assign node239 = (inp[8]) ? 3'b010 : 3'b011;
									assign node243 = (inp[8]) ? node245 : 3'b010;
										assign node245 = (inp[7]) ? 3'b011 : node246;
											assign node246 = (inp[11]) ? 3'b010 : 3'b010;
							assign node250 = (inp[7]) ? 3'b011 : node251;
								assign node251 = (inp[5]) ? node253 : 3'b011;
									assign node253 = (inp[10]) ? 3'b011 : node254;
										assign node254 = (inp[2]) ? 3'b011 : 3'b010;
						assign node259 = (inp[5]) ? node301 : node260;
							assign node260 = (inp[1]) ? node282 : node261;
								assign node261 = (inp[11]) ? node269 : node262;
									assign node262 = (inp[2]) ? node264 : 3'b011;
										assign node264 = (inp[7]) ? 3'b111 : node265;
											assign node265 = (inp[10]) ? 3'b111 : 3'b011;
									assign node269 = (inp[7]) ? node275 : node270;
										assign node270 = (inp[10]) ? node272 : 3'b111;
											assign node272 = (inp[8]) ? 3'b111 : 3'b011;
										assign node275 = (inp[10]) ? node279 : node276;
											assign node276 = (inp[2]) ? 3'b011 : 3'b111;
											assign node279 = (inp[2]) ? 3'b111 : 3'b011;
								assign node282 = (inp[10]) ? node294 : node283;
									assign node283 = (inp[2]) ? node289 : node284;
										assign node284 = (inp[8]) ? 3'b011 : node285;
											assign node285 = (inp[7]) ? 3'b011 : 3'b101;
										assign node289 = (inp[8]) ? 3'b111 : node290;
											assign node290 = (inp[11]) ? 3'b111 : 3'b011;
									assign node294 = (inp[8]) ? 3'b111 : node295;
										assign node295 = (inp[7]) ? 3'b111 : node296;
											assign node296 = (inp[2]) ? 3'b111 : 3'b011;
							assign node301 = (inp[7]) ? node331 : node302;
								assign node302 = (inp[11]) ? node318 : node303;
									assign node303 = (inp[10]) ? node311 : node304;
										assign node304 = (inp[2]) ? node308 : node305;
											assign node305 = (inp[8]) ? 3'b101 : 3'b111;
											assign node308 = (inp[8]) ? 3'b101 : 3'b001;
										assign node311 = (inp[2]) ? node315 : node312;
											assign node312 = (inp[1]) ? 3'b101 : 3'b001;
											assign node315 = (inp[1]) ? 3'b011 : 3'b111;
									assign node318 = (inp[8]) ? node326 : node319;
										assign node319 = (inp[1]) ? node323 : node320;
											assign node320 = (inp[10]) ? 3'b001 : 3'b011;
											assign node323 = (inp[2]) ? 3'b001 : 3'b011;
										assign node326 = (inp[1]) ? node328 : 3'b111;
											assign node328 = (inp[10]) ? 3'b011 : 3'b001;
								assign node331 = (inp[8]) ? node343 : node332;
									assign node332 = (inp[10]) ? node340 : node333;
										assign node333 = (inp[2]) ? node337 : node334;
											assign node334 = (inp[1]) ? 3'b111 : 3'b011;
											assign node337 = (inp[1]) ? 3'b011 : 3'b111;
										assign node340 = (inp[2]) ? 3'b111 : 3'b011;
									assign node343 = (inp[11]) ? node345 : 3'b011;
										assign node345 = (inp[10]) ? 3'b111 : node346;
											assign node346 = (inp[1]) ? 3'b011 : 3'b011;
				assign node350 = (inp[6]) ? 3'b111 : node351;
					assign node351 = (inp[1]) ? node443 : node352;
						assign node352 = (inp[7]) ? node404 : node353;
							assign node353 = (inp[9]) ? node381 : node354;
								assign node354 = (inp[5]) ? node368 : node355;
									assign node355 = (inp[10]) ? node361 : node356;
										assign node356 = (inp[11]) ? 3'b101 : node357;
											assign node357 = (inp[2]) ? 3'b011 : 3'b010;
										assign node361 = (inp[11]) ? node365 : node362;
											assign node362 = (inp[8]) ? 3'b001 : 3'b101;
											assign node365 = (inp[2]) ? 3'b011 : 3'b101;
									assign node368 = (inp[2]) ? node376 : node369;
										assign node369 = (inp[11]) ? node373 : node370;
											assign node370 = (inp[10]) ? 3'b010 : 3'b110;
											assign node373 = (inp[10]) ? 3'b110 : 3'b010;
										assign node376 = (inp[11]) ? 3'b110 : node377;
											assign node377 = (inp[10]) ? 3'b010 : 3'b010;
								assign node381 = (inp[5]) ? node395 : node382;
									assign node382 = (inp[8]) ? node390 : node383;
										assign node383 = (inp[11]) ? node387 : node384;
											assign node384 = (inp[10]) ? 3'b011 : 3'b001;
											assign node387 = (inp[10]) ? 3'b111 : 3'b011;
										assign node390 = (inp[11]) ? 3'b111 : node391;
											assign node391 = (inp[2]) ? 3'b111 : 3'b011;
									assign node395 = (inp[2]) ? node399 : node396;
										assign node396 = (inp[10]) ? 3'b101 : 3'b001;
										assign node399 = (inp[11]) ? node401 : 3'b011;
											assign node401 = (inp[8]) ? 3'b111 : 3'b011;
							assign node404 = (inp[9]) ? node430 : node405;
								assign node405 = (inp[2]) ? node417 : node406;
									assign node406 = (inp[11]) ? node412 : node407;
										assign node407 = (inp[8]) ? node409 : 3'b001;
											assign node409 = (inp[10]) ? 3'b001 : 3'b001;
										assign node412 = (inp[10]) ? 3'b011 : node413;
											assign node413 = (inp[5]) ? 3'b111 : 3'b101;
									assign node417 = (inp[5]) ? node423 : node418;
										assign node418 = (inp[10]) ? 3'b111 : node419;
											assign node419 = (inp[11]) ? 3'b011 : 3'b101;
										assign node423 = (inp[10]) ? node427 : node424;
											assign node424 = (inp[8]) ? 3'b101 : 3'b111;
											assign node427 = (inp[8]) ? 3'b101 : 3'b101;
								assign node430 = (inp[5]) ? node432 : 3'b111;
									assign node432 = (inp[2]) ? node438 : node433;
										assign node433 = (inp[10]) ? 3'b011 : node434;
											assign node434 = (inp[11]) ? 3'b011 : 3'b001;
										assign node438 = (inp[11]) ? node440 : 3'b011;
											assign node440 = (inp[10]) ? 3'b111 : 3'b011;
						assign node443 = (inp[9]) ? 3'b111 : node444;
							assign node444 = (inp[5]) ? node464 : node445;
								assign node445 = (inp[10]) ? node457 : node446;
									assign node446 = (inp[7]) ? node452 : node447;
										assign node447 = (inp[2]) ? node449 : 3'b011;
											assign node449 = (inp[8]) ? 3'b111 : 3'b011;
										assign node452 = (inp[8]) ? 3'b111 : node453;
											assign node453 = (inp[2]) ? 3'b111 : 3'b011;
									assign node457 = (inp[11]) ? 3'b111 : node458;
										assign node458 = (inp[7]) ? 3'b111 : node459;
											assign node459 = (inp[2]) ? 3'b111 : 3'b011;
								assign node464 = (inp[7]) ? node478 : node465;
									assign node465 = (inp[10]) ? node473 : node466;
										assign node466 = (inp[8]) ? node470 : node467;
											assign node467 = (inp[11]) ? 3'b001 : 3'b101;
											assign node470 = (inp[11]) ? 3'b001 : 3'b001;
										assign node473 = (inp[11]) ? 3'b011 : node474;
											assign node474 = (inp[2]) ? 3'b011 : 3'b101;
									assign node478 = (inp[10]) ? node486 : node479;
										assign node479 = (inp[2]) ? node483 : node480;
											assign node480 = (inp[8]) ? 3'b011 : 3'b111;
											assign node483 = (inp[8]) ? 3'b011 : 3'b011;
										assign node486 = (inp[11]) ? 3'b111 : node487;
											assign node487 = (inp[2]) ? 3'b011 : 3'b011;
			assign node493 = (inp[0]) ? node587 : node494;
				assign node494 = (inp[9]) ? node496 : 3'b000;
					assign node496 = (inp[6]) ? node562 : node497;
						assign node497 = (inp[7]) ? node527 : node498;
							assign node498 = (inp[1]) ? node508 : node499;
								assign node499 = (inp[5]) ? 3'b000 : node500;
									assign node500 = (inp[2]) ? node502 : 3'b000;
										assign node502 = (inp[8]) ? node504 : 3'b000;
											assign node504 = (inp[10]) ? 3'b100 : 3'b000;
								assign node508 = (inp[5]) ? node522 : node509;
									assign node509 = (inp[8]) ? node515 : node510;
										assign node510 = (inp[2]) ? node512 : 3'b100;
											assign node512 = (inp[10]) ? 3'b010 : 3'b100;
										assign node515 = (inp[10]) ? node519 : node516;
											assign node516 = (inp[2]) ? 3'b010 : 3'b100;
											assign node519 = (inp[11]) ? 3'b010 : 3'b010;
									assign node522 = (inp[11]) ? node524 : 3'b000;
										assign node524 = (inp[8]) ? 3'b000 : 3'b100;
							assign node527 = (inp[5]) ? node555 : node528;
								assign node528 = (inp[1]) ? node540 : node529;
									assign node529 = (inp[8]) ? node535 : node530;
										assign node530 = (inp[10]) ? node532 : 3'b100;
											assign node532 = (inp[11]) ? 3'b000 : 3'b000;
										assign node535 = (inp[2]) ? 3'b010 : node536;
											assign node536 = (inp[10]) ? 3'b100 : 3'b000;
									assign node540 = (inp[10]) ? node548 : node541;
										assign node541 = (inp[2]) ? node545 : node542;
											assign node542 = (inp[11]) ? 3'b100 : 3'b000;
											assign node545 = (inp[8]) ? 3'b110 : 3'b010;
										assign node548 = (inp[11]) ? node552 : node549;
											assign node549 = (inp[2]) ? 3'b010 : 3'b010;
											assign node552 = (inp[2]) ? 3'b110 : 3'b010;
								assign node555 = (inp[2]) ? node557 : 3'b100;
									assign node557 = (inp[11]) ? node559 : 3'b100;
										assign node559 = (inp[1]) ? 3'b010 : 3'b000;
						assign node562 = (inp[1]) ? node564 : 3'b000;
							assign node564 = (inp[7]) ? node578 : node565;
								assign node565 = (inp[5]) ? 3'b000 : node566;
									assign node566 = (inp[2]) ? node572 : node567;
										assign node567 = (inp[8]) ? node569 : 3'b000;
											assign node569 = (inp[11]) ? 3'b000 : 3'b000;
										assign node572 = (inp[11]) ? node574 : 3'b001;
											assign node574 = (inp[8]) ? 3'b000 : 3'b000;
								assign node578 = (inp[5]) ? node580 : 3'b001;
									assign node580 = (inp[2]) ? node582 : 3'b000;
										assign node582 = (inp[8]) ? 3'b001 : node583;
											assign node583 = (inp[11]) ? 3'b001 : 3'b000;
				assign node587 = (inp[9]) ? node665 : node588;
					assign node588 = (inp[6]) ? 3'b000 : node589;
						assign node589 = (inp[7]) ? node637 : node590;
							assign node590 = (inp[1]) ? node608 : node591;
								assign node591 = (inp[8]) ? node601 : node592;
									assign node592 = (inp[10]) ? node594 : 3'b100;
										assign node594 = (inp[11]) ? node598 : node595;
											assign node595 = (inp[5]) ? 3'b000 : 3'b010;
											assign node598 = (inp[2]) ? 3'b100 : 3'b000;
									assign node601 = (inp[5]) ? 3'b000 : node602;
										assign node602 = (inp[10]) ? 3'b010 : node603;
											assign node603 = (inp[2]) ? 3'b000 : 3'b100;
								assign node608 = (inp[5]) ? node622 : node609;
									assign node609 = (inp[10]) ? node615 : node610;
										assign node610 = (inp[2]) ? node612 : 3'b010;
											assign node612 = (inp[11]) ? 3'b110 : 3'b110;
										assign node615 = (inp[8]) ? node619 : node616;
											assign node616 = (inp[2]) ? 3'b101 : 3'b110;
											assign node619 = (inp[2]) ? 3'b101 : 3'b001;
									assign node622 = (inp[2]) ? node630 : node623;
										assign node623 = (inp[8]) ? node627 : node624;
											assign node624 = (inp[11]) ? 3'b100 : 3'b000;
											assign node627 = (inp[10]) ? 3'b000 : 3'b100;
										assign node630 = (inp[10]) ? node634 : node631;
											assign node631 = (inp[8]) ? 3'b010 : 3'b000;
											assign node634 = (inp[8]) ? 3'b110 : 3'b010;
							assign node637 = (inp[1]) ? node647 : node638;
								assign node638 = (inp[2]) ? node640 : 3'b110;
									assign node640 = (inp[8]) ? node642 : 3'b110;
										assign node642 = (inp[11]) ? 3'b110 : node643;
											assign node643 = (inp[10]) ? 3'b110 : 3'b110;
								assign node647 = (inp[5]) ? node657 : node648;
									assign node648 = (inp[8]) ? node650 : 3'b111;
										assign node650 = (inp[10]) ? node654 : node651;
											assign node651 = (inp[11]) ? 3'b110 : 3'b110;
											assign node654 = (inp[11]) ? 3'b110 : 3'b111;
									assign node657 = (inp[11]) ? node659 : 3'b110;
										assign node659 = (inp[2]) ? node661 : 3'b110;
											assign node661 = (inp[10]) ? 3'b111 : 3'b110;
					assign node665 = (inp[6]) ? node751 : node666;
						assign node666 = (inp[1]) ? node712 : node667;
							assign node667 = (inp[7]) ? node693 : node668;
								assign node668 = (inp[10]) ? node680 : node669;
									assign node669 = (inp[5]) ? node675 : node670;
										assign node670 = (inp[2]) ? 3'b110 : node671;
											assign node671 = (inp[11]) ? 3'b010 : 3'b010;
										assign node675 = (inp[2]) ? 3'b010 : node676;
											assign node676 = (inp[8]) ? 3'b100 : 3'b000;
									assign node680 = (inp[5]) ? node688 : node681;
										assign node681 = (inp[2]) ? node685 : node682;
											assign node682 = (inp[8]) ? 3'b001 : 3'b110;
											assign node685 = (inp[11]) ? 3'b101 : 3'b001;
										assign node688 = (inp[2]) ? 3'b110 : node689;
											assign node689 = (inp[11]) ? 3'b010 : 3'b000;
								assign node693 = (inp[2]) ? node701 : node694;
									assign node694 = (inp[5]) ? node696 : 3'b101;
										assign node696 = (inp[10]) ? node698 : 3'b100;
											assign node698 = (inp[8]) ? 3'b110 : 3'b100;
									assign node701 = (inp[11]) ? node707 : node702;
										assign node702 = (inp[5]) ? node704 : 3'b101;
											assign node704 = (inp[8]) ? 3'b111 : 3'b100;
										assign node707 = (inp[10]) ? node709 : 3'b011;
											assign node709 = (inp[5]) ? 3'b001 : 3'b011;
							assign node712 = (inp[5]) ? node726 : node713;
								assign node713 = (inp[7]) ? 3'b111 : node714;
									assign node714 = (inp[10]) ? node720 : node715;
										assign node715 = (inp[2]) ? node717 : 3'b101;
											assign node717 = (inp[11]) ? 3'b011 : 3'b101;
										assign node720 = (inp[11]) ? 3'b111 : node721;
											assign node721 = (inp[8]) ? 3'b011 : 3'b011;
								assign node726 = (inp[7]) ? node740 : node727;
									assign node727 = (inp[10]) ? node735 : node728;
										assign node728 = (inp[11]) ? node732 : node729;
											assign node729 = (inp[2]) ? 3'b100 : 3'b010;
											assign node732 = (inp[2]) ? 3'b001 : 3'b110;
										assign node735 = (inp[8]) ? 3'b101 : node736;
											assign node736 = (inp[2]) ? 3'b101 : 3'b001;
									assign node740 = (inp[8]) ? node744 : node741;
										assign node741 = (inp[10]) ? 3'b101 : 3'b001;
										assign node744 = (inp[11]) ? node748 : node745;
											assign node745 = (inp[10]) ? 3'b001 : 3'b001;
											assign node748 = (inp[2]) ? 3'b101 : 3'b011;
						assign node751 = (inp[10]) ? 3'b111 : node752;
							assign node752 = (inp[7]) ? 3'b111 : 3'b011;
		assign node756 = (inp[0]) ? node770 : node757;
			assign node757 = (inp[8]) ? node759 : 3'b000;
				assign node759 = (inp[11]) ? node761 : 3'b000;
					assign node761 = (inp[6]) ? 3'b000 : node762;
						assign node762 = (inp[7]) ? node764 : 3'b000;
							assign node764 = (inp[4]) ? 3'b000 : node765;
								assign node765 = (inp[9]) ? 3'b100 : 3'b000;
			assign node770 = (inp[4]) ? node922 : node771;
				assign node771 = (inp[9]) ? node791 : node772;
					assign node772 = (inp[6]) ? 3'b000 : node773;
						assign node773 = (inp[7]) ? 3'b100 : node774;
							assign node774 = (inp[5]) ? 3'b000 : node775;
								assign node775 = (inp[1]) ? node777 : 3'b000;
									assign node777 = (inp[2]) ? node783 : node778;
										assign node778 = (inp[8]) ? node780 : 3'b000;
											assign node780 = (inp[10]) ? 3'b100 : 3'b000;
										assign node783 = (inp[8]) ? node785 : 3'b100;
											assign node785 = (inp[11]) ? 3'b000 : 3'b100;
					assign node791 = (inp[6]) ? node877 : node792;
						assign node792 = (inp[1]) ? node822 : node793;
							assign node793 = (inp[5]) ? node815 : node794;
								assign node794 = (inp[11]) ? node802 : node795;
									assign node795 = (inp[2]) ? 3'b100 : node796;
										assign node796 = (inp[7]) ? node798 : 3'b000;
											assign node798 = (inp[8]) ? 3'b100 : 3'b000;
									assign node802 = (inp[7]) ? node808 : node803;
										assign node803 = (inp[2]) ? node805 : 3'b000;
											assign node805 = (inp[10]) ? 3'b000 : 3'b000;
										assign node808 = (inp[2]) ? node812 : node809;
											assign node809 = (inp[8]) ? 3'b000 : 3'b000;
											assign node812 = (inp[10]) ? 3'b110 : 3'b010;
								assign node815 = (inp[7]) ? node817 : 3'b000;
									assign node817 = (inp[2]) ? node819 : 3'b000;
										assign node819 = (inp[11]) ? 3'b100 : 3'b000;
							assign node822 = (inp[2]) ? node850 : node823;
								assign node823 = (inp[10]) ? node837 : node824;
									assign node824 = (inp[11]) ? node832 : node825;
										assign node825 = (inp[7]) ? node829 : node826;
											assign node826 = (inp[5]) ? 3'b000 : 3'b000;
											assign node829 = (inp[5]) ? 3'b000 : 3'b010;
										assign node832 = (inp[8]) ? node834 : 3'b100;
											assign node834 = (inp[5]) ? 3'b000 : 3'b000;
									assign node837 = (inp[11]) ? node845 : node838;
										assign node838 = (inp[5]) ? node842 : node839;
											assign node839 = (inp[7]) ? 3'b011 : 3'b010;
											assign node842 = (inp[7]) ? 3'b010 : 3'b000;
										assign node845 = (inp[8]) ? node847 : 3'b100;
											assign node847 = (inp[5]) ? 3'b010 : 3'b001;
								assign node850 = (inp[7]) ? node866 : node851;
									assign node851 = (inp[5]) ? node859 : node852;
										assign node852 = (inp[11]) ? node856 : node853;
											assign node853 = (inp[8]) ? 3'b010 : 3'b110;
											assign node856 = (inp[8]) ? 3'b001 : 3'b010;
										assign node859 = (inp[10]) ? node863 : node860;
											assign node860 = (inp[8]) ? 3'b100 : 3'b000;
											assign node863 = (inp[11]) ? 3'b010 : 3'b000;
									assign node866 = (inp[11]) ? node870 : node867;
										assign node867 = (inp[5]) ? 3'b100 : 3'b110;
										assign node870 = (inp[5]) ? node874 : node871;
											assign node871 = (inp[10]) ? 3'b101 : 3'b110;
											assign node874 = (inp[10]) ? 3'b110 : 3'b010;
						assign node877 = (inp[7]) ? node911 : node878;
							assign node878 = (inp[1]) ? node898 : node879;
								assign node879 = (inp[10]) ? node891 : node880;
									assign node880 = (inp[5]) ? node886 : node881;
										assign node881 = (inp[2]) ? node883 : 3'b010;
											assign node883 = (inp[11]) ? 3'b011 : 3'b010;
										assign node886 = (inp[8]) ? node888 : 3'b011;
											assign node888 = (inp[11]) ? 3'b010 : 3'b010;
									assign node891 = (inp[5]) ? node893 : 3'b011;
										assign node893 = (inp[2]) ? 3'b010 : node894;
											assign node894 = (inp[11]) ? 3'b010 : 3'b011;
								assign node898 = (inp[5]) ? node902 : node899;
									assign node899 = (inp[2]) ? 3'b011 : 3'b001;
									assign node902 = (inp[2]) ? node908 : node903;
										assign node903 = (inp[10]) ? 3'b011 : node904;
											assign node904 = (inp[8]) ? 3'b010 : 3'b010;
										assign node908 = (inp[11]) ? 3'b001 : 3'b011;
							assign node911 = (inp[1]) ? 3'b101 : node912;
								assign node912 = (inp[5]) ? node914 : 3'b101;
									assign node914 = (inp[10]) ? node916 : 3'b100;
										assign node916 = (inp[11]) ? 3'b101 : node917;
											assign node917 = (inp[8]) ? 3'b100 : 3'b101;
				assign node922 = (inp[1]) ? node924 : 3'b000;
					assign node924 = (inp[9]) ? node926 : 3'b000;
						assign node926 = (inp[6]) ? node942 : node927;
							assign node927 = (inp[5]) ? 3'b000 : node928;
								assign node928 = (inp[2]) ? node934 : node929;
									assign node929 = (inp[10]) ? node931 : 3'b000;
										assign node931 = (inp[8]) ? 3'b100 : 3'b000;
									assign node934 = (inp[7]) ? node938 : node935;
										assign node935 = (inp[11]) ? 3'b100 : 3'b000;
										assign node938 = (inp[11]) ? 3'b010 : 3'b100;
							assign node942 = (inp[7]) ? node956 : node943;
								assign node943 = (inp[8]) ? node947 : node944;
									assign node944 = (inp[11]) ? 3'b100 : 3'b000;
									assign node947 = (inp[11]) ? node951 : node948;
										assign node948 = (inp[5]) ? 3'b000 : 3'b100;
										assign node951 = (inp[5]) ? 3'b000 : node952;
											assign node952 = (inp[2]) ? 3'b000 : 3'b000;
								assign node956 = (inp[5]) ? node958 : 3'b110;
									assign node958 = (inp[2]) ? node962 : node959;
										assign node959 = (inp[8]) ? 3'b100 : 3'b000;
										assign node962 = (inp[11]) ? 3'b010 : node963;
											assign node963 = (inp[8]) ? 3'b010 : 3'b100;

endmodule