module dtc_split25_bm23 (
	input  wire [12-1:0] inp,
	output wire [12-1:0] outp
);

	wire [12-1:0] node1;
	wire [12-1:0] node2;
	wire [12-1:0] node3;
	wire [12-1:0] node4;
	wire [12-1:0] node5;
	wire [12-1:0] node6;
	wire [12-1:0] node7;
	wire [12-1:0] node8;
	wire [12-1:0] node9;
	wire [12-1:0] node13;
	wire [12-1:0] node14;
	wire [12-1:0] node16;
	wire [12-1:0] node19;
	wire [12-1:0] node22;
	wire [12-1:0] node23;
	wire [12-1:0] node24;
	wire [12-1:0] node28;
	wire [12-1:0] node29;
	wire [12-1:0] node31;
	wire [12-1:0] node32;
	wire [12-1:0] node37;
	wire [12-1:0] node38;
	wire [12-1:0] node39;
	wire [12-1:0] node40;
	wire [12-1:0] node41;
	wire [12-1:0] node45;
	wire [12-1:0] node48;
	wire [12-1:0] node49;
	wire [12-1:0] node53;
	wire [12-1:0] node54;
	wire [12-1:0] node56;
	wire [12-1:0] node58;
	wire [12-1:0] node61;
	wire [12-1:0] node62;
	wire [12-1:0] node66;
	wire [12-1:0] node67;
	wire [12-1:0] node68;
	wire [12-1:0] node69;
	wire [12-1:0] node71;
	wire [12-1:0] node74;
	wire [12-1:0] node75;
	wire [12-1:0] node79;
	wire [12-1:0] node80;
	wire [12-1:0] node81;
	wire [12-1:0] node83;
	wire [12-1:0] node87;
	wire [12-1:0] node90;
	wire [12-1:0] node91;
	wire [12-1:0] node92;
	wire [12-1:0] node94;
	wire [12-1:0] node96;
	wire [12-1:0] node99;
	wire [12-1:0] node100;
	wire [12-1:0] node104;
	wire [12-1:0] node106;
	wire [12-1:0] node109;
	wire [12-1:0] node110;
	wire [12-1:0] node111;
	wire [12-1:0] node112;
	wire [12-1:0] node113;
	wire [12-1:0] node114;
	wire [12-1:0] node115;
	wire [12-1:0] node118;
	wire [12-1:0] node119;
	wire [12-1:0] node124;
	wire [12-1:0] node127;
	wire [12-1:0] node128;
	wire [12-1:0] node129;
	wire [12-1:0] node133;
	wire [12-1:0] node136;
	wire [12-1:0] node137;
	wire [12-1:0] node138;
	wire [12-1:0] node139;
	wire [12-1:0] node143;
	wire [12-1:0] node144;
	wire [12-1:0] node147;
	wire [12-1:0] node150;
	wire [12-1:0] node152;
	wire [12-1:0] node153;
	wire [12-1:0] node157;
	wire [12-1:0] node158;
	wire [12-1:0] node159;
	wire [12-1:0] node160;
	wire [12-1:0] node162;
	wire [12-1:0] node166;
	wire [12-1:0] node167;
	wire [12-1:0] node168;
	wire [12-1:0] node172;
	wire [12-1:0] node173;
	wire [12-1:0] node177;
	wire [12-1:0] node178;
	wire [12-1:0] node179;
	wire [12-1:0] node181;
	wire [12-1:0] node182;
	wire [12-1:0] node184;
	wire [12-1:0] node188;
	wire [12-1:0] node190;
	wire [12-1:0] node193;
	wire [12-1:0] node194;
	wire [12-1:0] node198;
	wire [12-1:0] node199;
	wire [12-1:0] node200;
	wire [12-1:0] node201;
	wire [12-1:0] node202;
	wire [12-1:0] node203;
	wire [12-1:0] node204;
	wire [12-1:0] node208;
	wire [12-1:0] node209;
	wire [12-1:0] node213;
	wire [12-1:0] node214;
	wire [12-1:0] node215;
	wire [12-1:0] node219;
	wire [12-1:0] node220;
	wire [12-1:0] node222;
	wire [12-1:0] node226;
	wire [12-1:0] node227;
	wire [12-1:0] node228;
	wire [12-1:0] node229;
	wire [12-1:0] node233;
	wire [12-1:0] node235;
	wire [12-1:0] node238;
	wire [12-1:0] node239;
	wire [12-1:0] node241;
	wire [12-1:0] node244;
	wire [12-1:0] node246;
	wire [12-1:0] node247;
	wire [12-1:0] node248;
	wire [12-1:0] node253;
	wire [12-1:0] node254;
	wire [12-1:0] node255;
	wire [12-1:0] node256;
	wire [12-1:0] node257;
	wire [12-1:0] node258;
	wire [12-1:0] node263;
	wire [12-1:0] node264;
	wire [12-1:0] node265;
	wire [12-1:0] node267;
	wire [12-1:0] node271;
	wire [12-1:0] node274;
	wire [12-1:0] node275;
	wire [12-1:0] node276;
	wire [12-1:0] node280;
	wire [12-1:0] node283;
	wire [12-1:0] node284;
	wire [12-1:0] node286;
	wire [12-1:0] node287;
	wire [12-1:0] node291;
	wire [12-1:0] node293;
	wire [12-1:0] node294;
	wire [12-1:0] node296;
	wire [12-1:0] node298;
	wire [12-1:0] node301;
	wire [12-1:0] node304;
	wire [12-1:0] node305;
	wire [12-1:0] node306;
	wire [12-1:0] node307;
	wire [12-1:0] node308;
	wire [12-1:0] node311;
	wire [12-1:0] node314;
	wire [12-1:0] node315;
	wire [12-1:0] node317;
	wire [12-1:0] node318;
	wire [12-1:0] node322;
	wire [12-1:0] node323;
	wire [12-1:0] node325;
	wire [12-1:0] node326;
	wire [12-1:0] node330;
	wire [12-1:0] node333;
	wire [12-1:0] node334;
	wire [12-1:0] node335;
	wire [12-1:0] node338;
	wire [12-1:0] node339;
	wire [12-1:0] node343;
	wire [12-1:0] node344;
	wire [12-1:0] node345;
	wire [12-1:0] node348;
	wire [12-1:0] node350;
	wire [12-1:0] node353;
	wire [12-1:0] node354;
	wire [12-1:0] node358;
	wire [12-1:0] node359;
	wire [12-1:0] node360;
	wire [12-1:0] node361;
	wire [12-1:0] node363;
	wire [12-1:0] node364;
	wire [12-1:0] node366;
	wire [12-1:0] node370;
	wire [12-1:0] node371;
	wire [12-1:0] node372;
	wire [12-1:0] node376;
	wire [12-1:0] node379;
	wire [12-1:0] node380;
	wire [12-1:0] node382;
	wire [12-1:0] node385;
	wire [12-1:0] node386;
	wire [12-1:0] node390;
	wire [12-1:0] node391;
	wire [12-1:0] node392;
	wire [12-1:0] node394;
	wire [12-1:0] node398;
	wire [12-1:0] node399;
	wire [12-1:0] node400;
	wire [12-1:0] node401;
	wire [12-1:0] node405;
	wire [12-1:0] node408;
	wire [12-1:0] node410;
	wire [12-1:0] node413;
	wire [12-1:0] node414;
	wire [12-1:0] node415;
	wire [12-1:0] node416;
	wire [12-1:0] node417;
	wire [12-1:0] node418;
	wire [12-1:0] node419;
	wire [12-1:0] node420;
	wire [12-1:0] node421;
	wire [12-1:0] node426;
	wire [12-1:0] node429;
	wire [12-1:0] node431;
	wire [12-1:0] node432;
	wire [12-1:0] node436;
	wire [12-1:0] node437;
	wire [12-1:0] node438;
	wire [12-1:0] node439;
	wire [12-1:0] node442;
	wire [12-1:0] node446;
	wire [12-1:0] node447;
	wire [12-1:0] node448;
	wire [12-1:0] node452;
	wire [12-1:0] node453;
	wire [12-1:0] node455;
	wire [12-1:0] node459;
	wire [12-1:0] node460;
	wire [12-1:0] node461;
	wire [12-1:0] node462;
	wire [12-1:0] node463;
	wire [12-1:0] node467;
	wire [12-1:0] node468;
	wire [12-1:0] node470;
	wire [12-1:0] node471;
	wire [12-1:0] node475;
	wire [12-1:0] node478;
	wire [12-1:0] node479;
	wire [12-1:0] node480;
	wire [12-1:0] node481;
	wire [12-1:0] node483;
	wire [12-1:0] node488;
	wire [12-1:0] node491;
	wire [12-1:0] node492;
	wire [12-1:0] node493;
	wire [12-1:0] node497;
	wire [12-1:0] node498;
	wire [12-1:0] node500;
	wire [12-1:0] node503;
	wire [12-1:0] node506;
	wire [12-1:0] node507;
	wire [12-1:0] node508;
	wire [12-1:0] node509;
	wire [12-1:0] node511;
	wire [12-1:0] node514;
	wire [12-1:0] node515;
	wire [12-1:0] node517;
	wire [12-1:0] node520;
	wire [12-1:0] node521;
	wire [12-1:0] node522;
	wire [12-1:0] node526;
	wire [12-1:0] node529;
	wire [12-1:0] node530;
	wire [12-1:0] node533;
	wire [12-1:0] node535;
	wire [12-1:0] node536;
	wire [12-1:0] node538;
	wire [12-1:0] node542;
	wire [12-1:0] node543;
	wire [12-1:0] node544;
	wire [12-1:0] node545;
	wire [12-1:0] node548;
	wire [12-1:0] node549;
	wire [12-1:0] node551;
	wire [12-1:0] node552;
	wire [12-1:0] node556;
	wire [12-1:0] node559;
	wire [12-1:0] node561;
	wire [12-1:0] node562;
	wire [12-1:0] node563;
	wire [12-1:0] node568;
	wire [12-1:0] node569;
	wire [12-1:0] node570;
	wire [12-1:0] node572;
	wire [12-1:0] node574;
	wire [12-1:0] node575;
	wire [12-1:0] node579;
	wire [12-1:0] node582;
	wire [12-1:0] node583;
	wire [12-1:0] node586;
	wire [12-1:0] node587;
	wire [12-1:0] node588;
	wire [12-1:0] node592;
	wire [12-1:0] node595;
	wire [12-1:0] node596;
	wire [12-1:0] node597;
	wire [12-1:0] node598;
	wire [12-1:0] node599;
	wire [12-1:0] node600;
	wire [12-1:0] node601;
	wire [12-1:0] node605;
	wire [12-1:0] node607;
	wire [12-1:0] node610;
	wire [12-1:0] node611;
	wire [12-1:0] node612;
	wire [12-1:0] node616;
	wire [12-1:0] node617;
	wire [12-1:0] node619;
	wire [12-1:0] node622;
	wire [12-1:0] node625;
	wire [12-1:0] node626;
	wire [12-1:0] node627;
	wire [12-1:0] node628;
	wire [12-1:0] node633;
	wire [12-1:0] node634;
	wire [12-1:0] node635;
	wire [12-1:0] node638;
	wire [12-1:0] node642;
	wire [12-1:0] node643;
	wire [12-1:0] node644;
	wire [12-1:0] node645;
	wire [12-1:0] node646;
	wire [12-1:0] node648;
	wire [12-1:0] node651;
	wire [12-1:0] node654;
	wire [12-1:0] node655;
	wire [12-1:0] node659;
	wire [12-1:0] node660;
	wire [12-1:0] node661;
	wire [12-1:0] node664;
	wire [12-1:0] node667;
	wire [12-1:0] node670;
	wire [12-1:0] node671;
	wire [12-1:0] node672;
	wire [12-1:0] node673;
	wire [12-1:0] node676;
	wire [12-1:0] node679;
	wire [12-1:0] node682;
	wire [12-1:0] node683;
	wire [12-1:0] node684;
	wire [12-1:0] node687;
	wire [12-1:0] node688;
	wire [12-1:0] node692;
	wire [12-1:0] node695;
	wire [12-1:0] node696;
	wire [12-1:0] node697;
	wire [12-1:0] node698;
	wire [12-1:0] node699;
	wire [12-1:0] node700;
	wire [12-1:0] node704;
	wire [12-1:0] node705;
	wire [12-1:0] node707;
	wire [12-1:0] node710;
	wire [12-1:0] node712;
	wire [12-1:0] node715;
	wire [12-1:0] node717;
	wire [12-1:0] node720;
	wire [12-1:0] node721;
	wire [12-1:0] node722;
	wire [12-1:0] node725;
	wire [12-1:0] node726;
	wire [12-1:0] node730;
	wire [12-1:0] node732;
	wire [12-1:0] node733;
	wire [12-1:0] node737;
	wire [12-1:0] node738;
	wire [12-1:0] node739;
	wire [12-1:0] node740;
	wire [12-1:0] node741;
	wire [12-1:0] node742;
	wire [12-1:0] node746;
	wire [12-1:0] node749;
	wire [12-1:0] node752;
	wire [12-1:0] node753;
	wire [12-1:0] node755;
	wire [12-1:0] node758;
	wire [12-1:0] node759;
	wire [12-1:0] node763;
	wire [12-1:0] node764;
	wire [12-1:0] node765;
	wire [12-1:0] node767;
	wire [12-1:0] node769;
	wire [12-1:0] node771;
	wire [12-1:0] node774;
	wire [12-1:0] node776;
	wire [12-1:0] node779;
	wire [12-1:0] node781;
	wire [12-1:0] node782;
	wire [12-1:0] node784;
	wire [12-1:0] node787;
	wire [12-1:0] node790;
	wire [12-1:0] node791;
	wire [12-1:0] node792;
	wire [12-1:0] node793;
	wire [12-1:0] node794;
	wire [12-1:0] node795;
	wire [12-1:0] node796;
	wire [12-1:0] node797;
	wire [12-1:0] node799;
	wire [12-1:0] node800;
	wire [12-1:0] node804;
	wire [12-1:0] node807;
	wire [12-1:0] node808;
	wire [12-1:0] node812;
	wire [12-1:0] node813;
	wire [12-1:0] node814;
	wire [12-1:0] node816;
	wire [12-1:0] node819;
	wire [12-1:0] node821;
	wire [12-1:0] node822;
	wire [12-1:0] node823;
	wire [12-1:0] node828;
	wire [12-1:0] node829;
	wire [12-1:0] node831;
	wire [12-1:0] node833;
	wire [12-1:0] node836;
	wire [12-1:0] node837;
	wire [12-1:0] node840;
	wire [12-1:0] node843;
	wire [12-1:0] node844;
	wire [12-1:0] node845;
	wire [12-1:0] node846;
	wire [12-1:0] node849;
	wire [12-1:0] node852;
	wire [12-1:0] node853;
	wire [12-1:0] node855;
	wire [12-1:0] node858;
	wire [12-1:0] node860;
	wire [12-1:0] node863;
	wire [12-1:0] node864;
	wire [12-1:0] node865;
	wire [12-1:0] node869;
	wire [12-1:0] node871;
	wire [12-1:0] node872;
	wire [12-1:0] node876;
	wire [12-1:0] node877;
	wire [12-1:0] node878;
	wire [12-1:0] node879;
	wire [12-1:0] node881;
	wire [12-1:0] node883;
	wire [12-1:0] node886;
	wire [12-1:0] node887;
	wire [12-1:0] node889;
	wire [12-1:0] node892;
	wire [12-1:0] node894;
	wire [12-1:0] node897;
	wire [12-1:0] node898;
	wire [12-1:0] node899;
	wire [12-1:0] node900;
	wire [12-1:0] node904;
	wire [12-1:0] node906;
	wire [12-1:0] node909;
	wire [12-1:0] node910;
	wire [12-1:0] node912;
	wire [12-1:0] node914;
	wire [12-1:0] node915;
	wire [12-1:0] node920;
	wire [12-1:0] node921;
	wire [12-1:0] node922;
	wire [12-1:0] node923;
	wire [12-1:0] node925;
	wire [12-1:0] node926;
	wire [12-1:0] node931;
	wire [12-1:0] node932;
	wire [12-1:0] node934;
	wire [12-1:0] node935;
	wire [12-1:0] node939;
	wire [12-1:0] node941;
	wire [12-1:0] node942;
	wire [12-1:0] node946;
	wire [12-1:0] node947;
	wire [12-1:0] node948;
	wire [12-1:0] node950;
	wire [12-1:0] node953;
	wire [12-1:0] node955;
	wire [12-1:0] node958;
	wire [12-1:0] node961;
	wire [12-1:0] node962;
	wire [12-1:0] node963;
	wire [12-1:0] node964;
	wire [12-1:0] node965;
	wire [12-1:0] node967;
	wire [12-1:0] node968;
	wire [12-1:0] node971;
	wire [12-1:0] node974;
	wire [12-1:0] node975;
	wire [12-1:0] node976;
	wire [12-1:0] node977;
	wire [12-1:0] node983;
	wire [12-1:0] node984;
	wire [12-1:0] node985;
	wire [12-1:0] node986;
	wire [12-1:0] node990;
	wire [12-1:0] node991;
	wire [12-1:0] node994;
	wire [12-1:0] node996;
	wire [12-1:0] node997;
	wire [12-1:0] node1001;
	wire [12-1:0] node1002;
	wire [12-1:0] node1004;
	wire [12-1:0] node1007;
	wire [12-1:0] node1010;
	wire [12-1:0] node1011;
	wire [12-1:0] node1012;
	wire [12-1:0] node1014;
	wire [12-1:0] node1015;
	wire [12-1:0] node1018;
	wire [12-1:0] node1021;
	wire [12-1:0] node1023;
	wire [12-1:0] node1024;
	wire [12-1:0] node1028;
	wire [12-1:0] node1029;
	wire [12-1:0] node1031;
	wire [12-1:0] node1032;
	wire [12-1:0] node1036;
	wire [12-1:0] node1037;
	wire [12-1:0] node1038;
	wire [12-1:0] node1041;
	wire [12-1:0] node1043;
	wire [12-1:0] node1046;
	wire [12-1:0] node1049;
	wire [12-1:0] node1050;
	wire [12-1:0] node1051;
	wire [12-1:0] node1052;
	wire [12-1:0] node1054;
	wire [12-1:0] node1057;
	wire [12-1:0] node1058;
	wire [12-1:0] node1059;
	wire [12-1:0] node1061;
	wire [12-1:0] node1064;
	wire [12-1:0] node1067;
	wire [12-1:0] node1068;
	wire [12-1:0] node1072;
	wire [12-1:0] node1073;
	wire [12-1:0] node1075;
	wire [12-1:0] node1076;
	wire [12-1:0] node1077;
	wire [12-1:0] node1078;
	wire [12-1:0] node1083;
	wire [12-1:0] node1086;
	wire [12-1:0] node1087;
	wire [12-1:0] node1089;
	wire [12-1:0] node1092;
	wire [12-1:0] node1095;
	wire [12-1:0] node1096;
	wire [12-1:0] node1097;
	wire [12-1:0] node1099;
	wire [12-1:0] node1102;
	wire [12-1:0] node1103;
	wire [12-1:0] node1106;
	wire [12-1:0] node1107;
	wire [12-1:0] node1108;
	wire [12-1:0] node1112;
	wire [12-1:0] node1115;
	wire [12-1:0] node1116;
	wire [12-1:0] node1117;
	wire [12-1:0] node1119;
	wire [12-1:0] node1122;
	wire [12-1:0] node1123;
	wire [12-1:0] node1124;
	wire [12-1:0] node1128;
	wire [12-1:0] node1130;
	wire [12-1:0] node1133;
	wire [12-1:0] node1134;
	wire [12-1:0] node1135;
	wire [12-1:0] node1138;
	wire [12-1:0] node1141;
	wire [12-1:0] node1142;
	wire [12-1:0] node1145;
	wire [12-1:0] node1147;
	wire [12-1:0] node1149;
	wire [12-1:0] node1152;
	wire [12-1:0] node1153;
	wire [12-1:0] node1154;
	wire [12-1:0] node1155;
	wire [12-1:0] node1156;
	wire [12-1:0] node1157;
	wire [12-1:0] node1158;
	wire [12-1:0] node1159;
	wire [12-1:0] node1160;
	wire [12-1:0] node1165;
	wire [12-1:0] node1166;
	wire [12-1:0] node1170;
	wire [12-1:0] node1171;
	wire [12-1:0] node1172;
	wire [12-1:0] node1173;
	wire [12-1:0] node1178;
	wire [12-1:0] node1179;
	wire [12-1:0] node1182;
	wire [12-1:0] node1185;
	wire [12-1:0] node1186;
	wire [12-1:0] node1187;
	wire [12-1:0] node1188;
	wire [12-1:0] node1193;
	wire [12-1:0] node1194;
	wire [12-1:0] node1195;
	wire [12-1:0] node1198;
	wire [12-1:0] node1201;
	wire [12-1:0] node1204;
	wire [12-1:0] node1205;
	wire [12-1:0] node1206;
	wire [12-1:0] node1208;
	wire [12-1:0] node1209;
	wire [12-1:0] node1210;
	wire [12-1:0] node1215;
	wire [12-1:0] node1216;
	wire [12-1:0] node1217;
	wire [12-1:0] node1220;
	wire [12-1:0] node1223;
	wire [12-1:0] node1224;
	wire [12-1:0] node1227;
	wire [12-1:0] node1229;
	wire [12-1:0] node1232;
	wire [12-1:0] node1233;
	wire [12-1:0] node1234;
	wire [12-1:0] node1236;
	wire [12-1:0] node1238;
	wire [12-1:0] node1241;
	wire [12-1:0] node1243;
	wire [12-1:0] node1244;
	wire [12-1:0] node1248;
	wire [12-1:0] node1250;
	wire [12-1:0] node1252;
	wire [12-1:0] node1255;
	wire [12-1:0] node1256;
	wire [12-1:0] node1257;
	wire [12-1:0] node1258;
	wire [12-1:0] node1259;
	wire [12-1:0] node1261;
	wire [12-1:0] node1264;
	wire [12-1:0] node1265;
	wire [12-1:0] node1268;
	wire [12-1:0] node1269;
	wire [12-1:0] node1273;
	wire [12-1:0] node1274;
	wire [12-1:0] node1278;
	wire [12-1:0] node1279;
	wire [12-1:0] node1281;
	wire [12-1:0] node1283;
	wire [12-1:0] node1286;
	wire [12-1:0] node1287;
	wire [12-1:0] node1289;
	wire [12-1:0] node1292;
	wire [12-1:0] node1294;
	wire [12-1:0] node1297;
	wire [12-1:0] node1298;
	wire [12-1:0] node1299;
	wire [12-1:0] node1302;
	wire [12-1:0] node1304;
	wire [12-1:0] node1306;
	wire [12-1:0] node1309;
	wire [12-1:0] node1310;
	wire [12-1:0] node1311;
	wire [12-1:0] node1313;
	wire [12-1:0] node1315;
	wire [12-1:0] node1318;
	wire [12-1:0] node1321;
	wire [12-1:0] node1322;
	wire [12-1:0] node1323;
	wire [12-1:0] node1326;
	wire [12-1:0] node1329;
	wire [12-1:0] node1330;
	wire [12-1:0] node1333;
	wire [12-1:0] node1335;
	wire [12-1:0] node1338;
	wire [12-1:0] node1339;
	wire [12-1:0] node1340;
	wire [12-1:0] node1341;
	wire [12-1:0] node1342;
	wire [12-1:0] node1344;
	wire [12-1:0] node1347;
	wire [12-1:0] node1348;
	wire [12-1:0] node1351;
	wire [12-1:0] node1352;
	wire [12-1:0] node1353;
	wire [12-1:0] node1357;
	wire [12-1:0] node1360;
	wire [12-1:0] node1361;
	wire [12-1:0] node1362;
	wire [12-1:0] node1364;
	wire [12-1:0] node1368;
	wire [12-1:0] node1369;
	wire [12-1:0] node1370;
	wire [12-1:0] node1372;
	wire [12-1:0] node1375;
	wire [12-1:0] node1376;
	wire [12-1:0] node1381;
	wire [12-1:0] node1382;
	wire [12-1:0] node1383;
	wire [12-1:0] node1384;
	wire [12-1:0] node1385;
	wire [12-1:0] node1389;
	wire [12-1:0] node1390;
	wire [12-1:0] node1394;
	wire [12-1:0] node1395;
	wire [12-1:0] node1396;
	wire [12-1:0] node1400;
	wire [12-1:0] node1401;
	wire [12-1:0] node1403;
	wire [12-1:0] node1407;
	wire [12-1:0] node1408;
	wire [12-1:0] node1409;
	wire [12-1:0] node1411;
	wire [12-1:0] node1412;
	wire [12-1:0] node1417;
	wire [12-1:0] node1418;
	wire [12-1:0] node1419;
	wire [12-1:0] node1422;
	wire [12-1:0] node1424;
	wire [12-1:0] node1427;
	wire [12-1:0] node1428;
	wire [12-1:0] node1431;
	wire [12-1:0] node1432;
	wire [12-1:0] node1436;
	wire [12-1:0] node1437;
	wire [12-1:0] node1438;
	wire [12-1:0] node1439;
	wire [12-1:0] node1441;
	wire [12-1:0] node1444;
	wire [12-1:0] node1445;
	wire [12-1:0] node1446;
	wire [12-1:0] node1450;
	wire [12-1:0] node1451;
	wire [12-1:0] node1455;
	wire [12-1:0] node1456;
	wire [12-1:0] node1457;
	wire [12-1:0] node1460;
	wire [12-1:0] node1463;
	wire [12-1:0] node1464;
	wire [12-1:0] node1466;
	wire [12-1:0] node1468;
	wire [12-1:0] node1471;
	wire [12-1:0] node1474;
	wire [12-1:0] node1475;
	wire [12-1:0] node1476;
	wire [12-1:0] node1477;
	wire [12-1:0] node1478;
	wire [12-1:0] node1481;
	wire [12-1:0] node1484;
	wire [12-1:0] node1485;
	wire [12-1:0] node1488;
	wire [12-1:0] node1491;
	wire [12-1:0] node1492;
	wire [12-1:0] node1493;
	wire [12-1:0] node1494;
	wire [12-1:0] node1498;
	wire [12-1:0] node1499;
	wire [12-1:0] node1503;
	wire [12-1:0] node1504;
	wire [12-1:0] node1507;
	wire [12-1:0] node1510;
	wire [12-1:0] node1511;
	wire [12-1:0] node1512;
	wire [12-1:0] node1513;
	wire [12-1:0] node1516;
	wire [12-1:0] node1519;
	wire [12-1:0] node1520;
	wire [12-1:0] node1522;
	wire [12-1:0] node1524;
	wire [12-1:0] node1527;
	wire [12-1:0] node1530;
	wire [12-1:0] node1531;
	wire [12-1:0] node1532;
	wire [12-1:0] node1533;
	wire [12-1:0] node1537;
	wire [12-1:0] node1540;
	wire [12-1:0] node1542;

	assign outp = (inp[10]) ? node790 : node1;
		assign node1 = (inp[6]) ? node413 : node2;
			assign node2 = (inp[0]) ? node198 : node3;
				assign node3 = (inp[4]) ? node109 : node4;
					assign node4 = (inp[8]) ? node66 : node5;
						assign node5 = (inp[2]) ? node37 : node6;
							assign node6 = (inp[11]) ? node22 : node7;
								assign node7 = (inp[3]) ? node13 : node8;
									assign node8 = (inp[9]) ? 12'b001111111111 : node9;
										assign node9 = (inp[5]) ? 12'b011111111111 : 12'b111111111111;
									assign node13 = (inp[1]) ? node19 : node14;
										assign node14 = (inp[7]) ? node16 : 12'b001111111111;
											assign node16 = (inp[9]) ? 12'b000111111111 : 12'b001111111111;
										assign node19 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
								assign node22 = (inp[3]) ? node28 : node23;
									assign node23 = (inp[7]) ? 12'b000111111111 : node24;
										assign node24 = (inp[9]) ? 12'b000111111111 : 12'b001111111111;
									assign node28 = (inp[7]) ? 12'b000011111111 : node29;
										assign node29 = (inp[1]) ? node31 : 12'b000111111111;
											assign node31 = (inp[5]) ? 12'b000011111111 : node32;
												assign node32 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
							assign node37 = (inp[9]) ? node53 : node38;
								assign node38 = (inp[3]) ? node48 : node39;
									assign node39 = (inp[11]) ? node45 : node40;
										assign node40 = (inp[5]) ? 12'b000111111111 : node41;
											assign node41 = (inp[7]) ? 12'b001111111111 : 12'b011111111111;
										assign node45 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
									assign node48 = (inp[11]) ? 12'b000011111111 : node49;
										assign node49 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
								assign node53 = (inp[11]) ? node61 : node54;
									assign node54 = (inp[7]) ? node56 : 12'b000111111111;
										assign node56 = (inp[3]) ? node58 : 12'b000011111111;
											assign node58 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
									assign node61 = (inp[5]) ? 12'b000001111111 : node62;
										assign node62 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
						assign node66 = (inp[5]) ? node90 : node67;
							assign node67 = (inp[11]) ? node79 : node68;
								assign node68 = (inp[2]) ? node74 : node69;
									assign node69 = (inp[7]) ? node71 : 12'b011111111111;
										assign node71 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
									assign node74 = (inp[7]) ? 12'b000011111111 : node75;
										assign node75 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
								assign node79 = (inp[1]) ? node87 : node80;
									assign node80 = (inp[2]) ? 12'b000011111111 : node81;
										assign node81 = (inp[9]) ? node83 : 12'b000111111111;
											assign node83 = (inp[3]) ? 12'b000011111111 : 12'b000111111111;
									assign node87 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
							assign node90 = (inp[1]) ? node104 : node91;
								assign node91 = (inp[7]) ? node99 : node92;
									assign node92 = (inp[2]) ? node94 : 12'b001111111111;
										assign node94 = (inp[3]) ? node96 : 12'b000011111111;
											assign node96 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node99 = (inp[9]) ? 12'b000001111111 : node100;
										assign node100 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
								assign node104 = (inp[2]) ? node106 : 12'b000001111111;
									assign node106 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
					assign node109 = (inp[1]) ? node157 : node110;
						assign node110 = (inp[2]) ? node136 : node111;
							assign node111 = (inp[7]) ? node127 : node112;
								assign node112 = (inp[9]) ? node124 : node113;
									assign node113 = (inp[11]) ? 12'b000111111111 : node114;
										assign node114 = (inp[8]) ? node118 : node115;
											assign node115 = (inp[3]) ? 12'b001111111111 : 12'b011111111111;
											assign node118 = (inp[3]) ? 12'b000111111111 : node119;
												assign node119 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
									assign node124 = (inp[3]) ? 12'b000011111111 : 12'b001111111111;
								assign node127 = (inp[8]) ? node133 : node128;
									assign node128 = (inp[9]) ? 12'b000011111111 : node129;
										assign node129 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node133 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
							assign node136 = (inp[7]) ? node150 : node137;
								assign node137 = (inp[9]) ? node143 : node138;
									assign node138 = (inp[8]) ? 12'b000011111111 : node139;
										assign node139 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node143 = (inp[8]) ? node147 : node144;
										assign node144 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node147 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node150 = (inp[8]) ? node152 : 12'b000001111111;
									assign node152 = (inp[11]) ? 12'b000000011111 : node153;
										assign node153 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
						assign node157 = (inp[3]) ? node177 : node158;
							assign node158 = (inp[8]) ? node166 : node159;
								assign node159 = (inp[11]) ? 12'b000001111111 : node160;
									assign node160 = (inp[2]) ? node162 : 12'b000011111111;
										assign node162 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node166 = (inp[2]) ? node172 : node167;
									assign node167 = (inp[7]) ? 12'b000001111111 : node168;
										assign node168 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node172 = (inp[9]) ? 12'b000000011111 : node173;
										assign node173 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
							assign node177 = (inp[8]) ? node193 : node178;
								assign node178 = (inp[5]) ? node188 : node179;
									assign node179 = (inp[2]) ? node181 : 12'b000011111111;
										assign node181 = (inp[7]) ? 12'b000000111111 : node182;
											assign node182 = (inp[9]) ? node184 : 12'b000001111111;
												assign node184 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node188 = (inp[11]) ? node190 : 12'b000000111111;
										assign node190 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
								assign node193 = (inp[2]) ? 12'b000000011111 : node194;
									assign node194 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
				assign node198 = (inp[8]) ? node304 : node199;
					assign node199 = (inp[9]) ? node253 : node200;
						assign node200 = (inp[3]) ? node226 : node201;
							assign node201 = (inp[11]) ? node213 : node202;
								assign node202 = (inp[4]) ? node208 : node203;
									assign node203 = (inp[7]) ? 12'b000111111111 : node204;
										assign node204 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
									assign node208 = (inp[1]) ? 12'b000011111111 : node209;
										assign node209 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
								assign node213 = (inp[5]) ? node219 : node214;
									assign node214 = (inp[4]) ? 12'b000011111111 : node215;
										assign node215 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
									assign node219 = (inp[1]) ? 12'b000001111111 : node220;
										assign node220 = (inp[7]) ? node222 : 12'b000011111111;
											assign node222 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
							assign node226 = (inp[1]) ? node238 : node227;
								assign node227 = (inp[11]) ? node233 : node228;
									assign node228 = (inp[7]) ? 12'b000011111111 : node229;
										assign node229 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node233 = (inp[2]) ? node235 : 12'b000011111111;
										assign node235 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
								assign node238 = (inp[5]) ? node244 : node239;
									assign node239 = (inp[2]) ? node241 : 12'b000011111111;
										assign node241 = (inp[11]) ? 12'b000000011111 : 12'b000001111111;
									assign node244 = (inp[7]) ? node246 : 12'b000001111111;
										assign node246 = (inp[11]) ? 12'b000000111111 : node247;
											assign node247 = (inp[2]) ? 12'b000000111111 : node248;
												assign node248 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
						assign node253 = (inp[11]) ? node283 : node254;
							assign node254 = (inp[4]) ? node274 : node255;
								assign node255 = (inp[3]) ? node263 : node256;
									assign node256 = (inp[1]) ? 12'b000001111111 : node257;
										assign node257 = (inp[7]) ? 12'b000011111111 : node258;
											assign node258 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
									assign node263 = (inp[2]) ? node271 : node264;
										assign node264 = (inp[7]) ? 12'b000001111111 : node265;
											assign node265 = (inp[5]) ? node267 : 12'b000011111111;
												assign node267 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
										assign node271 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node274 = (inp[3]) ? node280 : node275;
									assign node275 = (inp[5]) ? 12'b000000111111 : node276;
										assign node276 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
									assign node280 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
							assign node283 = (inp[5]) ? node291 : node284;
								assign node284 = (inp[3]) ? node286 : 12'b000001111111;
									assign node286 = (inp[2]) ? 12'b000000011111 : node287;
										assign node287 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node291 = (inp[1]) ? node293 : 12'b000000111111;
									assign node293 = (inp[4]) ? node301 : node294;
										assign node294 = (inp[7]) ? node296 : 12'b000000111111;
											assign node296 = (inp[2]) ? node298 : 12'b000000011111;
												assign node298 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
										assign node301 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
					assign node304 = (inp[4]) ? node358 : node305;
						assign node305 = (inp[3]) ? node333 : node306;
							assign node306 = (inp[1]) ? node314 : node307;
								assign node307 = (inp[2]) ? node311 : node308;
									assign node308 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node311 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node314 = (inp[11]) ? node322 : node315;
									assign node315 = (inp[9]) ? node317 : 12'b000011111111;
										assign node317 = (inp[5]) ? 12'b000001111111 : node318;
											assign node318 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
									assign node322 = (inp[7]) ? node330 : node323;
										assign node323 = (inp[5]) ? node325 : 12'b000001111111;
											assign node325 = (inp[2]) ? 12'b000000111111 : node326;
												assign node326 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node330 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
							assign node333 = (inp[5]) ? node343 : node334;
								assign node334 = (inp[7]) ? node338 : node335;
									assign node335 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
									assign node338 = (inp[11]) ? 12'b000000011111 : node339;
										assign node339 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node343 = (inp[7]) ? node353 : node344;
									assign node344 = (inp[1]) ? node348 : node345;
										assign node345 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node348 = (inp[9]) ? node350 : 12'b000000111111;
											assign node350 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node353 = (inp[11]) ? 12'b000000011111 : node354;
										assign node354 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
						assign node358 = (inp[2]) ? node390 : node359;
							assign node359 = (inp[5]) ? node379 : node360;
								assign node360 = (inp[1]) ? node370 : node361;
									assign node361 = (inp[9]) ? node363 : 12'b000001111111;
										assign node363 = (inp[3]) ? 12'b000000111111 : node364;
											assign node364 = (inp[7]) ? node366 : 12'b000001111111;
												assign node366 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node370 = (inp[3]) ? node376 : node371;
										assign node371 = (inp[9]) ? 12'b000000111111 : node372;
											assign node372 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
										assign node376 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node379 = (inp[9]) ? node385 : node380;
									assign node380 = (inp[1]) ? node382 : 12'b000001111111;
										assign node382 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node385 = (inp[3]) ? 12'b000000011111 : node386;
										assign node386 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node390 = (inp[11]) ? node398 : node391;
								assign node391 = (inp[9]) ? 12'b000000011111 : node392;
									assign node392 = (inp[1]) ? node394 : 12'b000000111111;
										assign node394 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
								assign node398 = (inp[9]) ? node408 : node399;
									assign node399 = (inp[1]) ? node405 : node400;
										assign node400 = (inp[5]) ? 12'b000000011111 : node401;
											assign node401 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
										assign node405 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
									assign node408 = (inp[7]) ? node410 : 12'b000000001111;
										assign node410 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
			assign node413 = (inp[9]) ? node595 : node414;
				assign node414 = (inp[5]) ? node506 : node415;
					assign node415 = (inp[7]) ? node459 : node416;
						assign node416 = (inp[1]) ? node436 : node417;
							assign node417 = (inp[4]) ? node429 : node418;
								assign node418 = (inp[2]) ? node426 : node419;
									assign node419 = (inp[11]) ? 12'b000111111111 : node420;
										assign node420 = (inp[0]) ? 12'b000111111111 : node421;
											assign node421 = (inp[8]) ? 12'b001111111111 : 12'b011111111111;
									assign node426 = (inp[3]) ? 12'b000001111111 : 12'b000111111111;
								assign node429 = (inp[8]) ? node431 : 12'b000011111111;
									assign node431 = (inp[3]) ? 12'b000001111111 : node432;
										assign node432 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
							assign node436 = (inp[2]) ? node446 : node437;
								assign node437 = (inp[11]) ? 12'b000001111111 : node438;
									assign node438 = (inp[3]) ? node442 : node439;
										assign node439 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
										assign node442 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node446 = (inp[8]) ? node452 : node447;
									assign node447 = (inp[4]) ? 12'b000001111111 : node448;
										assign node448 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
									assign node452 = (inp[0]) ? 12'b000000111111 : node453;
										assign node453 = (inp[3]) ? node455 : 12'b000001111111;
											assign node455 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
						assign node459 = (inp[1]) ? node491 : node460;
							assign node460 = (inp[3]) ? node478 : node461;
								assign node461 = (inp[0]) ? node467 : node462;
									assign node462 = (inp[11]) ? 12'b000011111111 : node463;
										assign node463 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
									assign node467 = (inp[4]) ? node475 : node468;
										assign node468 = (inp[8]) ? node470 : 12'b000011111111;
											assign node470 = (inp[11]) ? 12'b000001111111 : node471;
												assign node471 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node475 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
								assign node478 = (inp[8]) ? node488 : node479;
									assign node479 = (inp[0]) ? 12'b000000111111 : node480;
										assign node480 = (inp[2]) ? 12'b000000111111 : node481;
											assign node481 = (inp[11]) ? node483 : 12'b000011111111;
												assign node483 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node488 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
							assign node491 = (inp[8]) ? node497 : node492;
								assign node492 = (inp[2]) ? 12'b000000111111 : node493;
									assign node493 = (inp[3]) ? 12'b000001111111 : 12'b000000111111;
								assign node497 = (inp[2]) ? node503 : node498;
									assign node498 = (inp[0]) ? node500 : 12'b000000011111;
										assign node500 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
									assign node503 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
					assign node506 = (inp[11]) ? node542 : node507;
						assign node507 = (inp[4]) ? node529 : node508;
							assign node508 = (inp[0]) ? node514 : node509;
								assign node509 = (inp[3]) ? node511 : 12'b000011111111;
									assign node511 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
								assign node514 = (inp[2]) ? node520 : node515;
									assign node515 = (inp[3]) ? node517 : 12'b000011111111;
										assign node517 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node520 = (inp[7]) ? node526 : node521;
										assign node521 = (inp[8]) ? 12'b000000111111 : node522;
											assign node522 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
										assign node526 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
							assign node529 = (inp[2]) ? node533 : node530;
								assign node530 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node533 = (inp[7]) ? node535 : 12'b000000111111;
									assign node535 = (inp[1]) ? 12'b000000011111 : node536;
										assign node536 = (inp[8]) ? node538 : 12'b000000111111;
											assign node538 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
						assign node542 = (inp[3]) ? node568 : node543;
							assign node543 = (inp[0]) ? node559 : node544;
								assign node544 = (inp[1]) ? node548 : node545;
									assign node545 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
									assign node548 = (inp[8]) ? node556 : node549;
										assign node549 = (inp[7]) ? node551 : 12'b000001111111;
											assign node551 = (inp[4]) ? 12'b000000111111 : node552;
												assign node552 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node556 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
								assign node559 = (inp[7]) ? node561 : 12'b000000111111;
									assign node561 = (inp[4]) ? 12'b000000000111 : node562;
										assign node562 = (inp[8]) ? 12'b000000011111 : node563;
											assign node563 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
							assign node568 = (inp[8]) ? node582 : node569;
								assign node569 = (inp[4]) ? node579 : node570;
									assign node570 = (inp[1]) ? node572 : 12'b000000111111;
										assign node572 = (inp[2]) ? node574 : 12'b000000111111;
											assign node574 = (inp[7]) ? 12'b000000011111 : node575;
												assign node575 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node579 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
								assign node582 = (inp[1]) ? node586 : node583;
									assign node583 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
									assign node586 = (inp[0]) ? node592 : node587;
										assign node587 = (inp[7]) ? 12'b000000001111 : node588;
											assign node588 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node592 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
				assign node595 = (inp[11]) ? node695 : node596;
					assign node596 = (inp[4]) ? node642 : node597;
						assign node597 = (inp[0]) ? node625 : node598;
							assign node598 = (inp[7]) ? node610 : node599;
								assign node599 = (inp[1]) ? node605 : node600;
									assign node600 = (inp[8]) ? 12'b000011111111 : node601;
										assign node601 = (inp[3]) ? 12'b000011111111 : 12'b000111111111;
									assign node605 = (inp[2]) ? node607 : 12'b000001111111;
										assign node607 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
								assign node610 = (inp[5]) ? node616 : node611;
									assign node611 = (inp[2]) ? 12'b000001111111 : node612;
										assign node612 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
									assign node616 = (inp[1]) ? node622 : node617;
										assign node617 = (inp[8]) ? node619 : 12'b000001111111;
											assign node619 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node622 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
							assign node625 = (inp[2]) ? node633 : node626;
								assign node626 = (inp[3]) ? 12'b000000111111 : node627;
									assign node627 = (inp[7]) ? 12'b000000111111 : node628;
										assign node628 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
								assign node633 = (inp[5]) ? 12'b000000001111 : node634;
									assign node634 = (inp[3]) ? node638 : node635;
										assign node635 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
										assign node638 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
						assign node642 = (inp[8]) ? node670 : node643;
							assign node643 = (inp[0]) ? node659 : node644;
								assign node644 = (inp[1]) ? node654 : node645;
									assign node645 = (inp[7]) ? node651 : node646;
										assign node646 = (inp[5]) ? node648 : 12'b000011111111;
											assign node648 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node651 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
									assign node654 = (inp[7]) ? 12'b000000111111 : node655;
										assign node655 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
								assign node659 = (inp[3]) ? node667 : node660;
									assign node660 = (inp[1]) ? node664 : node661;
										assign node661 = (inp[2]) ? 12'b000000111111 : 12'b000011111111;
										assign node664 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node667 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
							assign node670 = (inp[1]) ? node682 : node671;
								assign node671 = (inp[3]) ? node679 : node672;
									assign node672 = (inp[7]) ? node676 : node673;
										assign node673 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node676 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node679 = (inp[2]) ? 12'b000000011111 : 12'b000000001111;
								assign node682 = (inp[3]) ? node692 : node683;
									assign node683 = (inp[5]) ? node687 : node684;
										assign node684 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node687 = (inp[0]) ? 12'b000000001111 : node688;
											assign node688 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node692 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
					assign node695 = (inp[2]) ? node737 : node696;
						assign node696 = (inp[7]) ? node720 : node697;
							assign node697 = (inp[3]) ? node715 : node698;
								assign node698 = (inp[0]) ? node704 : node699;
									assign node699 = (inp[1]) ? 12'b000001111111 : node700;
										assign node700 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
									assign node704 = (inp[4]) ? node710 : node705;
										assign node705 = (inp[5]) ? node707 : 12'b000001111111;
											assign node707 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node710 = (inp[8]) ? node712 : 12'b000000111111;
											assign node712 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
								assign node715 = (inp[0]) ? node717 : 12'b000000111111;
									assign node717 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
							assign node720 = (inp[4]) ? node730 : node721;
								assign node721 = (inp[5]) ? node725 : node722;
									assign node722 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node725 = (inp[8]) ? 12'b000000011111 : node726;
										assign node726 = (inp[3]) ? 12'b000000011111 : 12'b000001111111;
								assign node730 = (inp[5]) ? node732 : 12'b000000011111;
									assign node732 = (inp[1]) ? 12'b000000001111 : node733;
										assign node733 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
						assign node737 = (inp[8]) ? node763 : node738;
							assign node738 = (inp[4]) ? node752 : node739;
								assign node739 = (inp[3]) ? node749 : node740;
									assign node740 = (inp[0]) ? node746 : node741;
										assign node741 = (inp[5]) ? 12'b000000111111 : node742;
											assign node742 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
										assign node746 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node749 = (inp[1]) ? 12'b000000011111 : 12'b000000001111;
								assign node752 = (inp[5]) ? node758 : node753;
									assign node753 = (inp[1]) ? node755 : 12'b000000011111;
										assign node755 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node758 = (inp[3]) ? 12'b000000000111 : node759;
										assign node759 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
							assign node763 = (inp[4]) ? node779 : node764;
								assign node764 = (inp[0]) ? node774 : node765;
									assign node765 = (inp[1]) ? node767 : 12'b000000011111;
										assign node767 = (inp[3]) ? node769 : 12'b000000011111;
											assign node769 = (inp[7]) ? node771 : 12'b000000001111;
												assign node771 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
									assign node774 = (inp[7]) ? node776 : 12'b000000001111;
										assign node776 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
								assign node779 = (inp[1]) ? node781 : 12'b000000001111;
									assign node781 = (inp[7]) ? node787 : node782;
										assign node782 = (inp[0]) ? node784 : 12'b000000000111;
											assign node784 = (inp[3]) ? 12'b000000000011 : 12'b000000000111;
										assign node787 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
		assign node790 = (inp[8]) ? node1152 : node791;
			assign node791 = (inp[2]) ? node961 : node792;
				assign node792 = (inp[6]) ? node876 : node793;
					assign node793 = (inp[7]) ? node843 : node794;
						assign node794 = (inp[3]) ? node812 : node795;
							assign node795 = (inp[4]) ? node807 : node796;
								assign node796 = (inp[11]) ? node804 : node797;
									assign node797 = (inp[9]) ? node799 : 12'b001111111111;
										assign node799 = (inp[0]) ? 12'b000111111111 : node800;
											assign node800 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
									assign node804 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
								assign node807 = (inp[5]) ? 12'b000001111111 : node808;
									assign node808 = (inp[1]) ? 12'b000001111111 : 12'b000111111111;
							assign node812 = (inp[1]) ? node828 : node813;
								assign node813 = (inp[0]) ? node819 : node814;
									assign node814 = (inp[4]) ? node816 : 12'b000011111111;
										assign node816 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node819 = (inp[5]) ? node821 : 12'b000111111111;
										assign node821 = (inp[11]) ? 12'b000001111111 : node822;
											assign node822 = (inp[4]) ? 12'b000001111111 : node823;
												assign node823 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node828 = (inp[11]) ? node836 : node829;
									assign node829 = (inp[5]) ? node831 : 12'b000011111111;
										assign node831 = (inp[0]) ? node833 : 12'b000011111111;
											assign node833 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
									assign node836 = (inp[4]) ? node840 : node837;
										assign node837 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node840 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
						assign node843 = (inp[1]) ? node863 : node844;
							assign node844 = (inp[3]) ? node852 : node845;
								assign node845 = (inp[4]) ? node849 : node846;
									assign node846 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node849 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
								assign node852 = (inp[4]) ? node858 : node853;
									assign node853 = (inp[9]) ? node855 : 12'b000001111111;
										assign node855 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
									assign node858 = (inp[9]) ? node860 : 12'b000000111111;
										assign node860 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node863 = (inp[3]) ? node869 : node864;
								assign node864 = (inp[4]) ? 12'b000000111111 : node865;
									assign node865 = (inp[0]) ? 12'b000001111111 : 12'b000000111111;
								assign node869 = (inp[0]) ? node871 : 12'b000000111111;
									assign node871 = (inp[5]) ? 12'b000000011111 : node872;
										assign node872 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
					assign node876 = (inp[5]) ? node920 : node877;
						assign node877 = (inp[1]) ? node897 : node878;
							assign node878 = (inp[9]) ? node886 : node879;
								assign node879 = (inp[4]) ? node881 : 12'b000011111111;
									assign node881 = (inp[7]) ? node883 : 12'b000011111111;
										assign node883 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node886 = (inp[7]) ? node892 : node887;
									assign node887 = (inp[4]) ? node889 : 12'b000011111111;
										assign node889 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
									assign node892 = (inp[11]) ? node894 : 12'b000000111111;
										assign node894 = (inp[0]) ? 12'b000000111111 : 12'b000000011111;
							assign node897 = (inp[7]) ? node909 : node898;
								assign node898 = (inp[9]) ? node904 : node899;
									assign node899 = (inp[0]) ? 12'b000001111111 : node900;
										assign node900 = (inp[4]) ? 12'b000000111111 : 12'b000011111111;
									assign node904 = (inp[3]) ? node906 : 12'b000000111111;
										assign node906 = (inp[4]) ? 12'b000000011111 : 12'b000001111111;
								assign node909 = (inp[9]) ? 12'b000000011111 : node910;
									assign node910 = (inp[0]) ? node912 : 12'b000001111111;
										assign node912 = (inp[3]) ? node914 : 12'b000000111111;
											assign node914 = (inp[11]) ? 12'b000000011111 : node915;
												assign node915 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
						assign node920 = (inp[9]) ? node946 : node921;
							assign node921 = (inp[11]) ? node931 : node922;
								assign node922 = (inp[1]) ? 12'b000000111111 : node923;
									assign node923 = (inp[7]) ? node925 : 12'b000001111111;
										assign node925 = (inp[0]) ? 12'b000000111111 : node926;
											assign node926 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
								assign node931 = (inp[0]) ? node939 : node932;
									assign node932 = (inp[7]) ? node934 : 12'b000000111111;
										assign node934 = (inp[4]) ? 12'b000000011111 : node935;
											assign node935 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node939 = (inp[1]) ? node941 : 12'b000000111111;
										assign node941 = (inp[7]) ? 12'b000000001111 : node942;
											assign node942 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
							assign node946 = (inp[3]) ? node958 : node947;
								assign node947 = (inp[1]) ? node953 : node948;
									assign node948 = (inp[0]) ? node950 : 12'b000000111111;
										assign node950 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node953 = (inp[0]) ? node955 : 12'b000000011111;
										assign node955 = (inp[7]) ? 12'b000000000111 : 12'b000000011111;
								assign node958 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
				assign node961 = (inp[9]) ? node1049 : node962;
					assign node962 = (inp[1]) ? node1010 : node963;
						assign node963 = (inp[3]) ? node983 : node964;
							assign node964 = (inp[6]) ? node974 : node965;
								assign node965 = (inp[11]) ? node967 : 12'b000011111111;
									assign node967 = (inp[0]) ? node971 : node968;
										assign node968 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node971 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
								assign node974 = (inp[11]) ? 12'b000000111111 : node975;
									assign node975 = (inp[0]) ? 12'b000000111111 : node976;
										assign node976 = (inp[5]) ? 12'b000001111111 : node977;
											assign node977 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
							assign node983 = (inp[7]) ? node1001 : node984;
								assign node984 = (inp[5]) ? node990 : node985;
									assign node985 = (inp[11]) ? 12'b000000011111 : node986;
										assign node986 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
									assign node990 = (inp[6]) ? node994 : node991;
										assign node991 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node994 = (inp[0]) ? node996 : 12'b000000111111;
											assign node996 = (inp[4]) ? 12'b000000011111 : node997;
												assign node997 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node1001 = (inp[0]) ? node1007 : node1002;
									assign node1002 = (inp[5]) ? node1004 : 12'b000000111111;
										assign node1004 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node1007 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
						assign node1010 = (inp[3]) ? node1028 : node1011;
							assign node1011 = (inp[6]) ? node1021 : node1012;
								assign node1012 = (inp[7]) ? node1014 : 12'b000001111111;
									assign node1014 = (inp[5]) ? node1018 : node1015;
										assign node1015 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1018 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node1021 = (inp[4]) ? node1023 : 12'b000000111111;
									assign node1023 = (inp[5]) ? 12'b000000011111 : node1024;
										assign node1024 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
							assign node1028 = (inp[4]) ? node1036 : node1029;
								assign node1029 = (inp[0]) ? node1031 : 12'b000001111111;
									assign node1031 = (inp[11]) ? 12'b000000011111 : node1032;
										assign node1032 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
								assign node1036 = (inp[7]) ? node1046 : node1037;
									assign node1037 = (inp[0]) ? node1041 : node1038;
										assign node1038 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node1041 = (inp[6]) ? node1043 : 12'b000000011111;
											assign node1043 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
									assign node1046 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
					assign node1049 = (inp[4]) ? node1095 : node1050;
						assign node1050 = (inp[6]) ? node1072 : node1051;
							assign node1051 = (inp[1]) ? node1057 : node1052;
								assign node1052 = (inp[5]) ? node1054 : 12'b000001111111;
									assign node1054 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node1057 = (inp[11]) ? node1067 : node1058;
									assign node1058 = (inp[7]) ? node1064 : node1059;
										assign node1059 = (inp[0]) ? node1061 : 12'b000001111111;
											assign node1061 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
										assign node1064 = (inp[0]) ? 12'b000000111111 : 12'b000000011111;
									assign node1067 = (inp[3]) ? 12'b000000011111 : node1068;
										assign node1068 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
							assign node1072 = (inp[0]) ? node1086 : node1073;
								assign node1073 = (inp[3]) ? node1075 : 12'b000000111111;
									assign node1075 = (inp[1]) ? node1083 : node1076;
										assign node1076 = (inp[7]) ? 12'b000000011111 : node1077;
											assign node1077 = (inp[11]) ? 12'b000000011111 : node1078;
												assign node1078 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node1083 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
								assign node1086 = (inp[3]) ? node1092 : node1087;
									assign node1087 = (inp[5]) ? node1089 : 12'b000000111111;
										assign node1089 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
									assign node1092 = (inp[5]) ? 12'b000000000011 : 12'b000000000111;
						assign node1095 = (inp[1]) ? node1115 : node1096;
							assign node1096 = (inp[11]) ? node1102 : node1097;
								assign node1097 = (inp[7]) ? node1099 : 12'b000000111111;
									assign node1099 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
								assign node1102 = (inp[6]) ? node1106 : node1103;
									assign node1103 = (inp[5]) ? 12'b000000111111 : 12'b000000011111;
									assign node1106 = (inp[5]) ? node1112 : node1107;
										assign node1107 = (inp[7]) ? 12'b000000001111 : node1108;
											assign node1108 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
										assign node1112 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
							assign node1115 = (inp[0]) ? node1133 : node1116;
								assign node1116 = (inp[7]) ? node1122 : node1117;
									assign node1117 = (inp[11]) ? node1119 : 12'b000000011111;
										assign node1119 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
									assign node1122 = (inp[3]) ? node1128 : node1123;
										assign node1123 = (inp[11]) ? 12'b000000001111 : node1124;
											assign node1124 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
										assign node1128 = (inp[6]) ? node1130 : 12'b000000001111;
											assign node1130 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
								assign node1133 = (inp[5]) ? node1141 : node1134;
									assign node1134 = (inp[3]) ? node1138 : node1135;
										assign node1135 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
										assign node1138 = (inp[6]) ? 12'b000000000111 : 12'b000000001111;
									assign node1141 = (inp[3]) ? node1145 : node1142;
										assign node1142 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
										assign node1145 = (inp[11]) ? node1147 : 12'b000000000111;
											assign node1147 = (inp[6]) ? node1149 : 12'b000000000011;
												assign node1149 = (inp[7]) ? 12'b000000000001 : 12'b000000000011;
			assign node1152 = (inp[5]) ? node1338 : node1153;
				assign node1153 = (inp[2]) ? node1255 : node1154;
					assign node1154 = (inp[1]) ? node1204 : node1155;
						assign node1155 = (inp[4]) ? node1185 : node1156;
							assign node1156 = (inp[3]) ? node1170 : node1157;
								assign node1157 = (inp[11]) ? node1165 : node1158;
									assign node1158 = (inp[9]) ? 12'b000011111111 : node1159;
										assign node1159 = (inp[0]) ? 12'b000011111111 : node1160;
											assign node1160 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
									assign node1165 = (inp[0]) ? 12'b000001111111 : node1166;
										assign node1166 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
								assign node1170 = (inp[6]) ? node1178 : node1171;
									assign node1171 = (inp[0]) ? 12'b000001111111 : node1172;
										assign node1172 = (inp[11]) ? 12'b000001111111 : node1173;
											assign node1173 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
									assign node1178 = (inp[11]) ? node1182 : node1179;
										assign node1179 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node1182 = (inp[0]) ? 12'b000000001111 : 12'b000000111111;
							assign node1185 = (inp[9]) ? node1193 : node1186;
								assign node1186 = (inp[3]) ? 12'b000000111111 : node1187;
									assign node1187 = (inp[6]) ? 12'b000001111111 : node1188;
										assign node1188 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node1193 = (inp[11]) ? node1201 : node1194;
									assign node1194 = (inp[6]) ? node1198 : node1195;
										assign node1195 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node1198 = (inp[7]) ? 12'b000000111111 : 12'b000000011111;
									assign node1201 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
						assign node1204 = (inp[7]) ? node1232 : node1205;
							assign node1205 = (inp[9]) ? node1215 : node1206;
								assign node1206 = (inp[0]) ? node1208 : 12'b000001111111;
									assign node1208 = (inp[11]) ? 12'b000000111111 : node1209;
										assign node1209 = (inp[3]) ? 12'b000000111111 : node1210;
											assign node1210 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
								assign node1215 = (inp[6]) ? node1223 : node1216;
									assign node1216 = (inp[0]) ? node1220 : node1217;
										assign node1217 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1220 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node1223 = (inp[11]) ? node1227 : node1224;
										assign node1224 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
										assign node1227 = (inp[4]) ? node1229 : 12'b000000011111;
											assign node1229 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
							assign node1232 = (inp[11]) ? node1248 : node1233;
								assign node1233 = (inp[0]) ? node1241 : node1234;
									assign node1234 = (inp[4]) ? node1236 : 12'b000001111111;
										assign node1236 = (inp[9]) ? node1238 : 12'b000000111111;
											assign node1238 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
									assign node1241 = (inp[6]) ? node1243 : 12'b000000011111;
										assign node1243 = (inp[3]) ? 12'b000000001111 : node1244;
											assign node1244 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node1248 = (inp[4]) ? node1250 : 12'b000000001111;
									assign node1250 = (inp[9]) ? node1252 : 12'b000000001111;
										assign node1252 = (inp[0]) ? 12'b000000000011 : 12'b000000001111;
					assign node1255 = (inp[3]) ? node1297 : node1256;
						assign node1256 = (inp[1]) ? node1278 : node1257;
							assign node1257 = (inp[7]) ? node1273 : node1258;
								assign node1258 = (inp[9]) ? node1264 : node1259;
									assign node1259 = (inp[4]) ? node1261 : 12'b000011111111;
										assign node1261 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node1264 = (inp[0]) ? node1268 : node1265;
										assign node1265 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1268 = (inp[6]) ? 12'b000000011111 : node1269;
											assign node1269 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
								assign node1273 = (inp[4]) ? 12'b000000001111 : node1274;
									assign node1274 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node1278 = (inp[6]) ? node1286 : node1279;
								assign node1279 = (inp[11]) ? node1281 : 12'b000000111111;
									assign node1281 = (inp[7]) ? node1283 : 12'b000000011111;
										assign node1283 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
								assign node1286 = (inp[11]) ? node1292 : node1287;
									assign node1287 = (inp[7]) ? node1289 : 12'b000000011111;
										assign node1289 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node1292 = (inp[4]) ? node1294 : 12'b000000001111;
										assign node1294 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
						assign node1297 = (inp[0]) ? node1309 : node1298;
							assign node1298 = (inp[6]) ? node1302 : node1299;
								assign node1299 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
								assign node1302 = (inp[4]) ? node1304 : 12'b000000011111;
									assign node1304 = (inp[7]) ? node1306 : 12'b000000001111;
										assign node1306 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
							assign node1309 = (inp[7]) ? node1321 : node1310;
								assign node1310 = (inp[9]) ? node1318 : node1311;
									assign node1311 = (inp[1]) ? node1313 : 12'b000000011111;
										assign node1313 = (inp[6]) ? node1315 : 12'b000000011111;
											assign node1315 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1318 = (inp[6]) ? 12'b000000000111 : 12'b000000001111;
								assign node1321 = (inp[11]) ? node1329 : node1322;
									assign node1322 = (inp[6]) ? node1326 : node1323;
										assign node1323 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
										assign node1326 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
									assign node1329 = (inp[1]) ? node1333 : node1330;
										assign node1330 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
										assign node1333 = (inp[9]) ? node1335 : 12'b000000000111;
											assign node1335 = (inp[4]) ? 12'b000000000001 : 12'b000000000011;
				assign node1338 = (inp[9]) ? node1436 : node1339;
					assign node1339 = (inp[3]) ? node1381 : node1340;
						assign node1340 = (inp[7]) ? node1360 : node1341;
							assign node1341 = (inp[6]) ? node1347 : node1342;
								assign node1342 = (inp[4]) ? node1344 : 12'b000001111111;
									assign node1344 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node1347 = (inp[2]) ? node1351 : node1348;
									assign node1348 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node1351 = (inp[4]) ? node1357 : node1352;
										assign node1352 = (inp[11]) ? 12'b000000011111 : node1353;
											assign node1353 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node1357 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
							assign node1360 = (inp[1]) ? node1368 : node1361;
								assign node1361 = (inp[11]) ? 12'b000000011111 : node1362;
									assign node1362 = (inp[6]) ? node1364 : 12'b000000111111;
										assign node1364 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
								assign node1368 = (inp[2]) ? 12'b000000001111 : node1369;
									assign node1369 = (inp[6]) ? node1375 : node1370;
										assign node1370 = (inp[4]) ? node1372 : 12'b000000011111;
											assign node1372 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node1375 = (inp[11]) ? 12'b000000011111 : node1376;
											assign node1376 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
						assign node1381 = (inp[6]) ? node1407 : node1382;
							assign node1382 = (inp[0]) ? node1394 : node1383;
								assign node1383 = (inp[11]) ? node1389 : node1384;
									assign node1384 = (inp[7]) ? 12'b000000111111 : node1385;
										assign node1385 = (inp[2]) ? 12'b000000111111 : 12'b000011111111;
									assign node1389 = (inp[1]) ? 12'b000000000111 : node1390;
										assign node1390 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
								assign node1394 = (inp[4]) ? node1400 : node1395;
									assign node1395 = (inp[1]) ? 12'b000000011111 : node1396;
										assign node1396 = (inp[11]) ? 12'b000000011111 : 12'b000001111111;
									assign node1400 = (inp[2]) ? 12'b000000001111 : node1401;
										assign node1401 = (inp[1]) ? node1403 : 12'b000000011111;
											assign node1403 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
							assign node1407 = (inp[1]) ? node1417 : node1408;
								assign node1408 = (inp[4]) ? 12'b000000001111 : node1409;
									assign node1409 = (inp[2]) ? node1411 : 12'b000000011111;
										assign node1411 = (inp[7]) ? 12'b000000001111 : node1412;
											assign node1412 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
								assign node1417 = (inp[0]) ? node1427 : node1418;
									assign node1418 = (inp[11]) ? node1422 : node1419;
										assign node1419 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node1422 = (inp[4]) ? node1424 : 12'b000000001111;
											assign node1424 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
									assign node1427 = (inp[7]) ? node1431 : node1428;
										assign node1428 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
										assign node1431 = (inp[2]) ? 12'b000000000011 : node1432;
											assign node1432 = (inp[11]) ? 12'b000000000011 : 12'b000000000111;
					assign node1436 = (inp[11]) ? node1474 : node1437;
						assign node1437 = (inp[0]) ? node1455 : node1438;
							assign node1438 = (inp[7]) ? node1444 : node1439;
								assign node1439 = (inp[6]) ? node1441 : 12'b000000111111;
									assign node1441 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
								assign node1444 = (inp[4]) ? node1450 : node1445;
									assign node1445 = (inp[2]) ? 12'b000000011111 : node1446;
										assign node1446 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node1450 = (inp[3]) ? 12'b000000000111 : node1451;
										assign node1451 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
							assign node1455 = (inp[2]) ? node1463 : node1456;
								assign node1456 = (inp[3]) ? node1460 : node1457;
									assign node1457 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
									assign node1460 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node1463 = (inp[6]) ? node1471 : node1464;
									assign node1464 = (inp[7]) ? node1466 : 12'b000000001111;
										assign node1466 = (inp[4]) ? node1468 : 12'b000000001111;
											assign node1468 = (inp[3]) ? 12'b000000000011 : 12'b000000001111;
									assign node1471 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
						assign node1474 = (inp[6]) ? node1510 : node1475;
							assign node1475 = (inp[3]) ? node1491 : node1476;
								assign node1476 = (inp[0]) ? node1484 : node1477;
									assign node1477 = (inp[1]) ? node1481 : node1478;
										assign node1478 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node1481 = (inp[4]) ? 12'b000000011111 : 12'b000000001111;
									assign node1484 = (inp[7]) ? node1488 : node1485;
										assign node1485 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node1488 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
								assign node1491 = (inp[7]) ? node1503 : node1492;
									assign node1492 = (inp[1]) ? node1498 : node1493;
										assign node1493 = (inp[2]) ? 12'b000000001111 : node1494;
											assign node1494 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node1498 = (inp[4]) ? 12'b000000000111 : node1499;
											assign node1499 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
									assign node1503 = (inp[0]) ? node1507 : node1504;
										assign node1504 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
										assign node1507 = (inp[1]) ? 12'b000000000011 : 12'b000000000111;
							assign node1510 = (inp[1]) ? node1530 : node1511;
								assign node1511 = (inp[4]) ? node1519 : node1512;
									assign node1512 = (inp[7]) ? node1516 : node1513;
										assign node1513 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
										assign node1516 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
									assign node1519 = (inp[0]) ? node1527 : node1520;
										assign node1520 = (inp[7]) ? node1522 : 12'b000000000111;
											assign node1522 = (inp[2]) ? node1524 : 12'b000000000111;
												assign node1524 = (inp[3]) ? 12'b000000000011 : 12'b000000000111;
										assign node1527 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
								assign node1530 = (inp[2]) ? node1540 : node1531;
									assign node1531 = (inp[4]) ? node1537 : node1532;
										assign node1532 = (inp[3]) ? 12'b000000000111 : node1533;
											assign node1533 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
										assign node1537 = (inp[0]) ? 12'b000000000011 : 12'b000000000111;
									assign node1540 = (inp[3]) ? node1542 : 12'b000000001111;
										assign node1542 = (inp[7]) ? 12'b000000000001 : 12'b000000000011;

endmodule