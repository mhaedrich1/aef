module dtc_split33_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node729;
	wire [3-1:0] node730;

	assign outp = (inp[6]) ? node196 : node1;
		assign node1 = (inp[9]) ? node175 : node2;
			assign node2 = (inp[0]) ? node116 : node3;
				assign node3 = (inp[10]) ? node75 : node4;
					assign node4 = (inp[7]) ? node44 : node5;
						assign node5 = (inp[1]) ? node27 : node6;
							assign node6 = (inp[11]) ? node14 : node7;
								assign node7 = (inp[3]) ? node9 : 3'b110;
									assign node9 = (inp[8]) ? node11 : 3'b110;
										assign node11 = (inp[5]) ? 3'b010 : 3'b110;
								assign node14 = (inp[8]) ? node20 : node15;
									assign node15 = (inp[3]) ? node17 : 3'b100;
										assign node17 = (inp[2]) ? 3'b000 : 3'b100;
									assign node20 = (inp[2]) ? 3'b010 : node21;
										assign node21 = (inp[4]) ? 3'b010 : node22;
											assign node22 = (inp[3]) ? 3'b010 : 3'b110;
							assign node27 = (inp[2]) ? node35 : node28;
								assign node28 = (inp[11]) ? node32 : node29;
									assign node29 = (inp[8]) ? 3'b010 : 3'b100;
									assign node32 = (inp[4]) ? 3'b000 : 3'b100;
								assign node35 = (inp[4]) ? node37 : 3'b100;
									assign node37 = (inp[3]) ? node39 : 3'b000;
										assign node39 = (inp[8]) ? node41 : 3'b000;
											assign node41 = (inp[11]) ? 3'b000 : 3'b100;
						assign node44 = (inp[1]) ? node58 : node45;
							assign node45 = (inp[4]) ? node51 : node46;
								assign node46 = (inp[11]) ? 3'b001 : node47;
									assign node47 = (inp[8]) ? 3'b101 : 3'b001;
								assign node51 = (inp[8]) ? node55 : node52;
									assign node52 = (inp[5]) ? 3'b110 : 3'b001;
									assign node55 = (inp[3]) ? 3'b001 : 3'b101;
							assign node58 = (inp[2]) ? node66 : node59;
								assign node59 = (inp[11]) ? node63 : node60;
									assign node60 = (inp[8]) ? 3'b001 : 3'b110;
									assign node63 = (inp[8]) ? 3'b110 : 3'b010;
								assign node66 = (inp[4]) ? node72 : node67;
									assign node67 = (inp[8]) ? node69 : 3'b010;
										assign node69 = (inp[5]) ? 3'b010 : 3'b110;
									assign node72 = (inp[3]) ? 3'b100 : 3'b110;
					assign node75 = (inp[7]) ? node83 : node76;
						assign node76 = (inp[11]) ? 3'b000 : node77;
							assign node77 = (inp[8]) ? node79 : 3'b000;
								assign node79 = (inp[1]) ? 3'b000 : 3'b100;
						assign node83 = (inp[1]) ? node101 : node84;
							assign node84 = (inp[8]) ? node94 : node85;
								assign node85 = (inp[11]) ? 3'b100 : node86;
									assign node86 = (inp[5]) ? node88 : 3'b010;
										assign node88 = (inp[4]) ? node90 : 3'b010;
											assign node90 = (inp[2]) ? 3'b100 : 3'b010;
								assign node94 = (inp[11]) ? node96 : 3'b110;
									assign node96 = (inp[5]) ? 3'b010 : node97;
										assign node97 = (inp[2]) ? 3'b010 : 3'b110;
							assign node101 = (inp[8]) ? node109 : node102;
								assign node102 = (inp[11]) ? 3'b000 : node103;
									assign node103 = (inp[2]) ? node105 : 3'b100;
										assign node105 = (inp[4]) ? 3'b100 : 3'b000;
								assign node109 = (inp[4]) ? 3'b100 : node110;
									assign node110 = (inp[2]) ? node112 : 3'b010;
										assign node112 = (inp[11]) ? 3'b100 : 3'b010;
				assign node116 = (inp[10]) ? node162 : node117;
					assign node117 = (inp[7]) ? node127 : node118;
						assign node118 = (inp[11]) ? 3'b000 : node119;
							assign node119 = (inp[2]) ? 3'b000 : node120;
								assign node120 = (inp[1]) ? 3'b000 : node121;
									assign node121 = (inp[8]) ? 3'b100 : 3'b000;
						assign node127 = (inp[1]) ? node143 : node128;
							assign node128 = (inp[11]) ? node136 : node129;
								assign node129 = (inp[8]) ? node133 : node130;
									assign node130 = (inp[2]) ? 3'b100 : 3'b010;
									assign node133 = (inp[2]) ? 3'b010 : 3'b110;
								assign node136 = (inp[8]) ? node140 : node137;
									assign node137 = (inp[2]) ? 3'b000 : 3'b100;
									assign node140 = (inp[2]) ? 3'b100 : 3'b010;
							assign node143 = (inp[2]) ? node157 : node144;
								assign node144 = (inp[8]) ? node150 : node145;
									assign node145 = (inp[3]) ? 3'b000 : node146;
										assign node146 = (inp[11]) ? 3'b000 : 3'b100;
									assign node150 = (inp[4]) ? node152 : 3'b100;
										assign node152 = (inp[3]) ? 3'b100 : node153;
											assign node153 = (inp[11]) ? 3'b100 : 3'b010;
								assign node157 = (inp[11]) ? 3'b000 : node158;
									assign node158 = (inp[8]) ? 3'b100 : 3'b000;
					assign node162 = (inp[1]) ? 3'b000 : node163;
						assign node163 = (inp[11]) ? 3'b000 : node164;
							assign node164 = (inp[8]) ? node166 : 3'b000;
								assign node166 = (inp[7]) ? node168 : 3'b000;
									assign node168 = (inp[4]) ? node170 : 3'b100;
										assign node170 = (inp[2]) ? 3'b000 : 3'b100;
			assign node175 = (inp[0]) ? 3'b000 : node176;
				assign node176 = (inp[7]) ? node178 : 3'b000;
					assign node178 = (inp[10]) ? 3'b000 : node179;
						assign node179 = (inp[1]) ? 3'b000 : node180;
							assign node180 = (inp[11]) ? 3'b000 : node181;
								assign node181 = (inp[2]) ? node189 : node182;
									assign node182 = (inp[8]) ? node184 : 3'b100;
										assign node184 = (inp[3]) ? node186 : 3'b010;
											assign node186 = (inp[5]) ? 3'b100 : 3'b010;
									assign node189 = (inp[8]) ? 3'b100 : 3'b000;
		assign node196 = (inp[9]) ? node496 : node197;
			assign node197 = (inp[0]) ? node325 : node198;
				assign node198 = (inp[7]) ? node278 : node199;
					assign node199 = (inp[10]) ? node239 : node200;
						assign node200 = (inp[8]) ? node220 : node201;
							assign node201 = (inp[1]) ? node213 : node202;
								assign node202 = (inp[11]) ? node208 : node203;
									assign node203 = (inp[3]) ? 3'b011 : node204;
										assign node204 = (inp[2]) ? 3'b011 : 3'b111;
									assign node208 = (inp[2]) ? 3'b101 : node209;
										assign node209 = (inp[3]) ? 3'b101 : 3'b011;
								assign node213 = (inp[11]) ? node215 : 3'b101;
									assign node215 = (inp[2]) ? 3'b001 : node216;
										assign node216 = (inp[4]) ? 3'b001 : 3'b101;
							assign node220 = (inp[11]) ? node230 : node221;
								assign node221 = (inp[1]) ? node223 : 3'b111;
									assign node223 = (inp[2]) ? 3'b011 : node224;
										assign node224 = (inp[4]) ? 3'b011 : node225;
											assign node225 = (inp[5]) ? 3'b111 : 3'b011;
								assign node230 = (inp[1]) ? 3'b101 : node231;
									assign node231 = (inp[5]) ? node233 : 3'b111;
										assign node233 = (inp[3]) ? 3'b011 : node234;
											assign node234 = (inp[2]) ? 3'b011 : 3'b111;
						assign node239 = (inp[1]) ? node251 : node240;
							assign node240 = (inp[8]) ? node246 : node241;
								assign node241 = (inp[11]) ? 3'b110 : node242;
									assign node242 = (inp[2]) ? 3'b001 : 3'b101;
								assign node246 = (inp[2]) ? node248 : 3'b011;
									assign node248 = (inp[11]) ? 3'b001 : 3'b101;
							assign node251 = (inp[8]) ? node265 : node252;
								assign node252 = (inp[4]) ? node258 : node253;
									assign node253 = (inp[11]) ? node255 : 3'b110;
										assign node255 = (inp[2]) ? 3'b010 : 3'b110;
									assign node258 = (inp[11]) ? 3'b010 : node259;
										assign node259 = (inp[3]) ? node261 : 3'b110;
											assign node261 = (inp[2]) ? 3'b010 : 3'b110;
								assign node265 = (inp[11]) ? node275 : node266;
									assign node266 = (inp[3]) ? node270 : node267;
										assign node267 = (inp[2]) ? 3'b001 : 3'b101;
										assign node270 = (inp[5]) ? node272 : 3'b001;
											assign node272 = (inp[2]) ? 3'b110 : 3'b001;
									assign node275 = (inp[2]) ? 3'b110 : 3'b001;
					assign node278 = (inp[10]) ? node294 : node279;
						assign node279 = (inp[8]) ? 3'b111 : node280;
							assign node280 = (inp[1]) ? node282 : 3'b111;
								assign node282 = (inp[2]) ? node284 : 3'b111;
									assign node284 = (inp[5]) ? node288 : node285;
										assign node285 = (inp[11]) ? 3'b011 : 3'b111;
										assign node288 = (inp[11]) ? 3'b101 : node289;
											assign node289 = (inp[3]) ? 3'b011 : 3'b111;
						assign node294 = (inp[11]) ? node312 : node295;
							assign node295 = (inp[2]) ? node305 : node296;
								assign node296 = (inp[3]) ? node302 : node297;
									assign node297 = (inp[8]) ? 3'b111 : node298;
										assign node298 = (inp[5]) ? 3'b011 : 3'b111;
									assign node302 = (inp[1]) ? 3'b101 : 3'b111;
								assign node305 = (inp[5]) ? node307 : 3'b111;
									assign node307 = (inp[3]) ? node309 : 3'b011;
										assign node309 = (inp[1]) ? 3'b011 : 3'b111;
							assign node312 = (inp[8]) ? node320 : node313;
								assign node313 = (inp[1]) ? node315 : 3'b101;
									assign node315 = (inp[3]) ? 3'b001 : node316;
										assign node316 = (inp[2]) ? 3'b001 : 3'b101;
								assign node320 = (inp[1]) ? 3'b101 : node321;
									assign node321 = (inp[3]) ? 3'b011 : 3'b111;
				assign node325 = (inp[7]) ? node397 : node326;
					assign node326 = (inp[10]) ? node364 : node327;
						assign node327 = (inp[8]) ? node343 : node328;
							assign node328 = (inp[5]) ? node336 : node329;
								assign node329 = (inp[2]) ? node333 : node330;
									assign node330 = (inp[3]) ? 3'b110 : 3'b010;
									assign node333 = (inp[1]) ? 3'b100 : 3'b110;
								assign node336 = (inp[2]) ? 3'b010 : node337;
									assign node337 = (inp[11]) ? node339 : 3'b001;
										assign node339 = (inp[1]) ? 3'b100 : 3'b110;
							assign node343 = (inp[1]) ? node353 : node344;
								assign node344 = (inp[11]) ? node348 : node345;
									assign node345 = (inp[2]) ? 3'b001 : 3'b101;
									assign node348 = (inp[2]) ? node350 : 3'b001;
										assign node350 = (inp[3]) ? 3'b110 : 3'b001;
								assign node353 = (inp[11]) ? node361 : node354;
									assign node354 = (inp[2]) ? 3'b110 : node355;
										assign node355 = (inp[3]) ? node357 : 3'b001;
											assign node357 = (inp[4]) ? 3'b110 : 3'b001;
									assign node361 = (inp[2]) ? 3'b010 : 3'b110;
						assign node364 = (inp[8]) ? node378 : node365;
							assign node365 = (inp[11]) ? node371 : node366;
								assign node366 = (inp[1]) ? node368 : 3'b010;
									assign node368 = (inp[2]) ? 3'b000 : 3'b100;
								assign node371 = (inp[1]) ? 3'b000 : node372;
									assign node372 = (inp[2]) ? node374 : 3'b100;
										assign node374 = (inp[3]) ? 3'b000 : 3'b100;
							assign node378 = (inp[2]) ? node390 : node379;
								assign node379 = (inp[1]) ? node387 : node380;
									assign node380 = (inp[11]) ? node382 : 3'b110;
										assign node382 = (inp[5]) ? 3'b010 : node383;
											assign node383 = (inp[4]) ? 3'b010 : 3'b110;
									assign node387 = (inp[11]) ? 3'b100 : 3'b010;
								assign node390 = (inp[1]) ? 3'b100 : node391;
									assign node391 = (inp[11]) ? 3'b100 : node392;
										assign node392 = (inp[3]) ? 3'b010 : 3'b110;
					assign node397 = (inp[10]) ? node441 : node398;
						assign node398 = (inp[8]) ? node414 : node399;
							assign node399 = (inp[1]) ? node405 : node400;
								assign node400 = (inp[11]) ? 3'b101 : node401;
									assign node401 = (inp[4]) ? 3'b101 : 3'b011;
								assign node405 = (inp[11]) ? node411 : node406;
									assign node406 = (inp[4]) ? node408 : 3'b101;
										assign node408 = (inp[2]) ? 3'b001 : 3'b101;
									assign node411 = (inp[2]) ? 3'b110 : 3'b001;
							assign node414 = (inp[1]) ? node428 : node415;
								assign node415 = (inp[11]) ? node421 : node416;
									assign node416 = (inp[3]) ? node418 : 3'b111;
										assign node418 = (inp[2]) ? 3'b011 : 3'b111;
									assign node421 = (inp[2]) ? 3'b011 : node422;
										assign node422 = (inp[3]) ? 3'b011 : node423;
											assign node423 = (inp[5]) ? 3'b111 : 3'b011;
								assign node428 = (inp[11]) ? node432 : node429;
									assign node429 = (inp[5]) ? 3'b101 : 3'b011;
									assign node432 = (inp[2]) ? node434 : 3'b101;
										assign node434 = (inp[3]) ? 3'b001 : node435;
											assign node435 = (inp[4]) ? node437 : 3'b101;
												assign node437 = (inp[5]) ? 3'b001 : 3'b101;
						assign node441 = (inp[11]) ? node469 : node442;
							assign node442 = (inp[8]) ? node452 : node443;
								assign node443 = (inp[1]) ? node449 : node444;
									assign node444 = (inp[2]) ? 3'b110 : node445;
										assign node445 = (inp[4]) ? 3'b001 : 3'b101;
									assign node449 = (inp[2]) ? 3'b010 : 3'b110;
								assign node452 = (inp[2]) ? node460 : node453;
									assign node453 = (inp[1]) ? 3'b001 : node454;
										assign node454 = (inp[3]) ? 3'b101 : node455;
											assign node455 = (inp[4]) ? 3'b101 : 3'b011;
									assign node460 = (inp[1]) ? node464 : node461;
										assign node461 = (inp[5]) ? 3'b101 : 3'b001;
										assign node464 = (inp[3]) ? 3'b110 : node465;
											assign node465 = (inp[5]) ? 3'b110 : 3'b001;
							assign node469 = (inp[4]) ? node481 : node470;
								assign node470 = (inp[8]) ? node478 : node471;
									assign node471 = (inp[1]) ? node473 : 3'b110;
										assign node473 = (inp[5]) ? 3'b010 : node474;
											assign node474 = (inp[2]) ? 3'b100 : 3'b010;
									assign node478 = (inp[1]) ? 3'b110 : 3'b101;
								assign node481 = (inp[8]) ? node489 : node482;
									assign node482 = (inp[1]) ? node486 : node483;
										assign node483 = (inp[3]) ? 3'b010 : 3'b110;
										assign node486 = (inp[2]) ? 3'b100 : 3'b010;
									assign node489 = (inp[1]) ? node493 : node490;
										assign node490 = (inp[3]) ? 3'b001 : 3'b011;
										assign node493 = (inp[2]) ? 3'b010 : 3'b110;
			assign node496 = (inp[0]) ? node666 : node497;
				assign node497 = (inp[7]) ? node571 : node498;
					assign node498 = (inp[10]) ? node546 : node499;
						assign node499 = (inp[8]) ? node517 : node500;
							assign node500 = (inp[1]) ? node508 : node501;
								assign node501 = (inp[2]) ? 3'b100 : node502;
									assign node502 = (inp[5]) ? node504 : 3'b100;
										assign node504 = (inp[11]) ? 3'b010 : 3'b110;
								assign node508 = (inp[11]) ? 3'b000 : node509;
									assign node509 = (inp[4]) ? node513 : node510;
										assign node510 = (inp[2]) ? 3'b100 : 3'b010;
										assign node513 = (inp[2]) ? 3'b000 : 3'b100;
							assign node517 = (inp[2]) ? node533 : node518;
								assign node518 = (inp[11]) ? node524 : node519;
									assign node519 = (inp[1]) ? node521 : 3'b001;
										assign node521 = (inp[3]) ? 3'b010 : 3'b110;
									assign node524 = (inp[3]) ? node526 : 3'b010;
										assign node526 = (inp[1]) ? 3'b100 : node527;
											assign node527 = (inp[5]) ? node529 : 3'b110;
												assign node529 = (inp[4]) ? 3'b010 : 3'b110;
								assign node533 = (inp[5]) ? node541 : node534;
									assign node534 = (inp[1]) ? 3'b010 : node535;
										assign node535 = (inp[11]) ? node537 : 3'b110;
											assign node537 = (inp[4]) ? 3'b010 : 3'b110;
									assign node541 = (inp[1]) ? node543 : 3'b010;
										assign node543 = (inp[11]) ? 3'b100 : 3'b010;
						assign node546 = (inp[2]) ? 3'b000 : node547;
							assign node547 = (inp[5]) ? node553 : node548;
								assign node548 = (inp[11]) ? 3'b000 : node549;
									assign node549 = (inp[3]) ? 3'b000 : 3'b100;
								assign node553 = (inp[11]) ? node567 : node554;
									assign node554 = (inp[3]) ? node560 : node555;
										assign node555 = (inp[1]) ? node557 : 3'b010;
											assign node557 = (inp[8]) ? 3'b100 : 3'b000;
										assign node560 = (inp[1]) ? 3'b000 : node561;
											assign node561 = (inp[8]) ? 3'b100 : node562;
												assign node562 = (inp[4]) ? 3'b000 : 3'b100;
									assign node567 = (inp[1]) ? 3'b000 : 3'b100;
					assign node571 = (inp[10]) ? node623 : node572;
						assign node572 = (inp[1]) ? node592 : node573;
							assign node573 = (inp[8]) ? node585 : node574;
								assign node574 = (inp[5]) ? node576 : 3'b001;
									assign node576 = (inp[2]) ? node582 : node577;
										assign node577 = (inp[3]) ? 3'b001 : node578;
											assign node578 = (inp[11]) ? 3'b001 : 3'b101;
										assign node582 = (inp[4]) ? 3'b001 : 3'b110;
								assign node585 = (inp[2]) ? node589 : node586;
									assign node586 = (inp[11]) ? 3'b101 : 3'b011;
									assign node589 = (inp[11]) ? 3'b001 : 3'b101;
							assign node592 = (inp[2]) ? node608 : node593;
								assign node593 = (inp[3]) ? node599 : node594;
									assign node594 = (inp[8]) ? node596 : 3'b001;
										assign node596 = (inp[11]) ? 3'b001 : 3'b101;
									assign node599 = (inp[11]) ? node605 : node600;
										assign node600 = (inp[8]) ? node602 : 3'b110;
											assign node602 = (inp[4]) ? 3'b001 : 3'b101;
										assign node605 = (inp[4]) ? 3'b110 : 3'b010;
								assign node608 = (inp[4]) ? node616 : node609;
									assign node609 = (inp[3]) ? node611 : 3'b110;
										assign node611 = (inp[11]) ? node613 : 3'b110;
											assign node613 = (inp[8]) ? 3'b110 : 3'b010;
									assign node616 = (inp[3]) ? 3'b110 : node617;
										assign node617 = (inp[11]) ? node619 : 3'b001;
											assign node619 = (inp[8]) ? 3'b110 : 3'b010;
						assign node623 = (inp[1]) ? node651 : node624;
							assign node624 = (inp[3]) ? node636 : node625;
								assign node625 = (inp[11]) ? node631 : node626;
									assign node626 = (inp[8]) ? 3'b001 : node627;
										assign node627 = (inp[4]) ? 3'b010 : 3'b110;
									assign node631 = (inp[8]) ? node633 : 3'b100;
										assign node633 = (inp[5]) ? 3'b010 : 3'b110;
								assign node636 = (inp[11]) ? node644 : node637;
									assign node637 = (inp[2]) ? node641 : node638;
										assign node638 = (inp[8]) ? 3'b001 : 3'b110;
										assign node641 = (inp[8]) ? 3'b110 : 3'b010;
									assign node644 = (inp[4]) ? node646 : 3'b010;
										assign node646 = (inp[5]) ? node648 : 3'b010;
											assign node648 = (inp[8]) ? 3'b110 : 3'b010;
							assign node651 = (inp[8]) ? node661 : node652;
								assign node652 = (inp[4]) ? node654 : 3'b100;
									assign node654 = (inp[3]) ? 3'b000 : node655;
										assign node655 = (inp[2]) ? node657 : 3'b100;
											assign node657 = (inp[11]) ? 3'b000 : 3'b100;
								assign node661 = (inp[2]) ? node663 : 3'b010;
									assign node663 = (inp[11]) ? 3'b100 : 3'b010;
				assign node666 = (inp[10]) ? node720 : node667;
					assign node667 = (inp[7]) ? node679 : node668;
						assign node668 = (inp[8]) ? node670 : 3'b000;
							assign node670 = (inp[1]) ? 3'b000 : node671;
								assign node671 = (inp[11]) ? node673 : 3'b100;
									assign node673 = (inp[2]) ? 3'b000 : node674;
										assign node674 = (inp[3]) ? 3'b000 : 3'b100;
						assign node679 = (inp[3]) ? node699 : node680;
							assign node680 = (inp[8]) ? node690 : node681;
								assign node681 = (inp[1]) ? node687 : node682;
									assign node682 = (inp[2]) ? node684 : 3'b010;
										assign node684 = (inp[11]) ? 3'b100 : 3'b010;
									assign node687 = (inp[11]) ? 3'b000 : 3'b100;
								assign node690 = (inp[1]) ? 3'b010 : node691;
									assign node691 = (inp[5]) ? node695 : node692;
										assign node692 = (inp[11]) ? 3'b110 : 3'b001;
										assign node695 = (inp[11]) ? 3'b010 : 3'b110;
							assign node699 = (inp[1]) ? node709 : node700;
								assign node700 = (inp[11]) ? node702 : 3'b110;
									assign node702 = (inp[8]) ? node704 : 3'b100;
										assign node704 = (inp[2]) ? node706 : 3'b010;
											assign node706 = (inp[4]) ? 3'b100 : 3'b000;
								assign node709 = (inp[11]) ? node715 : node710;
									assign node710 = (inp[2]) ? node712 : 3'b100;
										assign node712 = (inp[8]) ? 3'b100 : 3'b000;
									assign node715 = (inp[8]) ? node717 : 3'b000;
										assign node717 = (inp[2]) ? 3'b000 : 3'b100;
					assign node720 = (inp[1]) ? 3'b000 : node721;
						assign node721 = (inp[7]) ? node723 : 3'b000;
							assign node723 = (inp[8]) ? node725 : 3'b000;
								assign node725 = (inp[11]) ? node729 : node726;
									assign node726 = (inp[3]) ? 3'b100 : 3'b011;
									assign node729 = (inp[2]) ? 3'b000 : node730;
										assign node730 = (inp[3]) ? 3'b000 : 3'b100;

endmodule