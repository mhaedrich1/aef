module dtc_split75_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node430;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node460;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node467;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node678;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node795;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node909;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node979;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node991;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1004;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1035;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1056;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1064;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1071;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1085;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1097;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1114;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1193;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1206;
	wire [3-1:0] node1210;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1224;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1232;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1252;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;

	assign outp = (inp[6]) ? node372 : node1;
		assign node1 = (inp[9]) ? node333 : node2;
			assign node2 = (inp[0]) ? node248 : node3;
				assign node3 = (inp[7]) ? node103 : node4;
					assign node4 = (inp[10]) ? node78 : node5;
						assign node5 = (inp[1]) ? node53 : node6;
							assign node6 = (inp[8]) ? node30 : node7;
								assign node7 = (inp[2]) ? node19 : node8;
									assign node8 = (inp[11]) ? node14 : node9;
										assign node9 = (inp[4]) ? 3'b110 : node10;
											assign node10 = (inp[5]) ? 3'b110 : 3'b100;
										assign node14 = (inp[3]) ? 3'b100 : node15;
											assign node15 = (inp[4]) ? 3'b100 : 3'b110;
									assign node19 = (inp[3]) ? 3'b000 : node20;
										assign node20 = (inp[11]) ? node24 : node21;
											assign node21 = (inp[5]) ? 3'b010 : 3'b110;
											assign node24 = (inp[5]) ? node26 : 3'b100;
												assign node26 = (inp[4]) ? 3'b000 : 3'b100;
								assign node30 = (inp[11]) ? node46 : node31;
									assign node31 = (inp[2]) ? node39 : node32;
										assign node32 = (inp[4]) ? 3'b110 : node33;
											assign node33 = (inp[3]) ? 3'b110 : node34;
												assign node34 = (inp[5]) ? 3'b110 : 3'b010;
										assign node39 = (inp[3]) ? node41 : 3'b110;
											assign node41 = (inp[4]) ? 3'b010 : node42;
												assign node42 = (inp[5]) ? 3'b010 : 3'b110;
									assign node46 = (inp[4]) ? 3'b010 : node47;
										assign node47 = (inp[3]) ? 3'b010 : node48;
											assign node48 = (inp[2]) ? 3'b010 : 3'b110;
							assign node53 = (inp[11]) ? node69 : node54;
								assign node54 = (inp[8]) ? node60 : node55;
									assign node55 = (inp[2]) ? node57 : 3'b100;
										assign node57 = (inp[3]) ? 3'b000 : 3'b100;
									assign node60 = (inp[2]) ? node62 : 3'b010;
										assign node62 = (inp[3]) ? 3'b100 : node63;
											assign node63 = (inp[5]) ? node65 : 3'b010;
												assign node65 = (inp[4]) ? 3'b100 : 3'b010;
								assign node69 = (inp[8]) ? node71 : 3'b000;
									assign node71 = (inp[2]) ? node73 : 3'b100;
										assign node73 = (inp[3]) ? 3'b000 : node74;
											assign node74 = (inp[5]) ? 3'b000 : 3'b100;
						assign node78 = (inp[8]) ? node80 : 3'b000;
							assign node80 = (inp[1]) ? 3'b000 : node81;
								assign node81 = (inp[11]) ? node97 : node82;
									assign node82 = (inp[2]) ? node90 : node83;
										assign node83 = (inp[3]) ? 3'b100 : node84;
											assign node84 = (inp[5]) ? node86 : 3'b000;
												assign node86 = (inp[4]) ? 3'b100 : 3'b000;
										assign node90 = (inp[3]) ? node92 : 3'b100;
											assign node92 = (inp[4]) ? node94 : 3'b100;
												assign node94 = (inp[5]) ? 3'b000 : 3'b100;
									assign node97 = (inp[3]) ? 3'b000 : node98;
										assign node98 = (inp[4]) ? 3'b000 : 3'b100;
					assign node103 = (inp[10]) ? node171 : node104;
						assign node104 = (inp[1]) ? node138 : node105;
							assign node105 = (inp[8]) ? node131 : node106;
								assign node106 = (inp[11]) ? node118 : node107;
									assign node107 = (inp[3]) ? node113 : node108;
										assign node108 = (inp[2]) ? 3'b001 : node109;
											assign node109 = (inp[4]) ? 3'b001 : 3'b101;
										assign node113 = (inp[2]) ? node115 : 3'b001;
											assign node115 = (inp[4]) ? 3'b110 : 3'b001;
									assign node118 = (inp[2]) ? node126 : node119;
										assign node119 = (inp[3]) ? 3'b110 : node120;
											assign node120 = (inp[5]) ? node122 : 3'b001;
												assign node122 = (inp[4]) ? 3'b110 : 3'b001;
										assign node126 = (inp[3]) ? node128 : 3'b110;
											assign node128 = (inp[4]) ? 3'b010 : 3'b110;
								assign node131 = (inp[11]) ? node133 : 3'b101;
									assign node133 = (inp[2]) ? 3'b001 : node134;
										assign node134 = (inp[3]) ? 3'b001 : 3'b101;
							assign node138 = (inp[8]) ? node154 : node139;
								assign node139 = (inp[11]) ? node149 : node140;
									assign node140 = (inp[2]) ? node142 : 3'b110;
										assign node142 = (inp[3]) ? 3'b010 : node143;
											assign node143 = (inp[5]) ? node145 : 3'b110;
												assign node145 = (inp[4]) ? 3'b010 : 3'b110;
									assign node149 = (inp[2]) ? node151 : 3'b010;
										assign node151 = (inp[3]) ? 3'b100 : 3'b010;
								assign node154 = (inp[11]) ? node160 : node155;
									assign node155 = (inp[3]) ? node157 : 3'b001;
										assign node157 = (inp[2]) ? 3'b110 : 3'b001;
									assign node160 = (inp[2]) ? node166 : node161;
										assign node161 = (inp[5]) ? 3'b110 : node162;
											assign node162 = (inp[3]) ? 3'b110 : 3'b001;
										assign node166 = (inp[3]) ? node168 : 3'b110;
											assign node168 = (inp[4]) ? 3'b010 : 3'b110;
						assign node171 = (inp[1]) ? node207 : node172;
							assign node172 = (inp[8]) ? node196 : node173;
								assign node173 = (inp[11]) ? node185 : node174;
									assign node174 = (inp[2]) ? node180 : node175;
										assign node175 = (inp[3]) ? 3'b010 : node176;
											assign node176 = (inp[4]) ? 3'b010 : 3'b110;
										assign node180 = (inp[3]) ? node182 : 3'b010;
											assign node182 = (inp[4]) ? 3'b100 : 3'b010;
									assign node185 = (inp[3]) ? node189 : node186;
										assign node186 = (inp[2]) ? 3'b100 : 3'b010;
										assign node189 = (inp[4]) ? node191 : 3'b100;
											assign node191 = (inp[5]) ? node193 : 3'b100;
												assign node193 = (inp[2]) ? 3'b000 : 3'b100;
								assign node196 = (inp[11]) ? node202 : node197;
									assign node197 = (inp[3]) ? 3'b110 : node198;
										assign node198 = (inp[2]) ? 3'b110 : 3'b001;
									assign node202 = (inp[3]) ? 3'b010 : node203;
										assign node203 = (inp[2]) ? 3'b010 : 3'b110;
							assign node207 = (inp[8]) ? node219 : node208;
								assign node208 = (inp[11]) ? node214 : node209;
									assign node209 = (inp[2]) ? node211 : 3'b100;
										assign node211 = (inp[3]) ? 3'b000 : 3'b100;
									assign node214 = (inp[3]) ? 3'b000 : node215;
										assign node215 = (inp[4]) ? 3'b000 : 3'b100;
								assign node219 = (inp[11]) ? node235 : node220;
									assign node220 = (inp[3]) ? node228 : node221;
										assign node221 = (inp[5]) ? 3'b010 : node222;
											assign node222 = (inp[4]) ? 3'b010 : node223;
												assign node223 = (inp[2]) ? 3'b010 : 3'b110;
										assign node228 = (inp[2]) ? node230 : 3'b010;
											assign node230 = (inp[5]) ? 3'b100 : node231;
												assign node231 = (inp[4]) ? 3'b100 : 3'b010;
									assign node235 = (inp[3]) ? node241 : node236;
										assign node236 = (inp[2]) ? 3'b100 : node237;
											assign node237 = (inp[4]) ? 3'b100 : 3'b010;
										assign node241 = (inp[2]) ? node243 : 3'b100;
											assign node243 = (inp[4]) ? 3'b000 : node244;
												assign node244 = (inp[5]) ? 3'b000 : 3'b100;
				assign node248 = (inp[7]) ? node264 : node249;
					assign node249 = (inp[10]) ? 3'b000 : node250;
						assign node250 = (inp[8]) ? node252 : 3'b000;
							assign node252 = (inp[2]) ? 3'b000 : node253;
								assign node253 = (inp[11]) ? 3'b000 : node254;
									assign node254 = (inp[1]) ? 3'b000 : node255;
										assign node255 = (inp[3]) ? node257 : 3'b100;
											assign node257 = (inp[4]) ? 3'b000 : 3'b100;
					assign node264 = (inp[10]) ? node318 : node265;
						assign node265 = (inp[1]) ? node295 : node266;
							assign node266 = (inp[8]) ? node280 : node267;
								assign node267 = (inp[11]) ? node275 : node268;
									assign node268 = (inp[2]) ? node270 : 3'b010;
										assign node270 = (inp[4]) ? 3'b100 : node271;
											assign node271 = (inp[3]) ? 3'b100 : 3'b010;
									assign node275 = (inp[2]) ? node277 : 3'b100;
										assign node277 = (inp[4]) ? 3'b000 : 3'b100;
								assign node280 = (inp[11]) ? node288 : node281;
									assign node281 = (inp[2]) ? node283 : 3'b110;
										assign node283 = (inp[3]) ? 3'b010 : node284;
											assign node284 = (inp[5]) ? 3'b010 : 3'b110;
									assign node288 = (inp[2]) ? node290 : 3'b010;
										assign node290 = (inp[3]) ? 3'b100 : node291;
											assign node291 = (inp[4]) ? 3'b100 : 3'b010;
							assign node295 = (inp[8]) ? node303 : node296;
								assign node296 = (inp[3]) ? 3'b000 : node297;
									assign node297 = (inp[2]) ? 3'b000 : node298;
										assign node298 = (inp[11]) ? 3'b000 : 3'b100;
								assign node303 = (inp[11]) ? node313 : node304;
									assign node304 = (inp[2]) ? 3'b100 : node305;
										assign node305 = (inp[3]) ? node307 : 3'b010;
											assign node307 = (inp[4]) ? 3'b100 : node308;
												assign node308 = (inp[5]) ? 3'b100 : 3'b010;
									assign node313 = (inp[2]) ? 3'b000 : node314;
										assign node314 = (inp[3]) ? 3'b000 : 3'b100;
						assign node318 = (inp[11]) ? 3'b000 : node319;
							assign node319 = (inp[8]) ? node321 : 3'b000;
								assign node321 = (inp[2]) ? node325 : node322;
									assign node322 = (inp[1]) ? 3'b000 : 3'b100;
									assign node325 = (inp[3]) ? 3'b000 : node326;
										assign node326 = (inp[1]) ? 3'b000 : node327;
											assign node327 = (inp[4]) ? 3'b000 : 3'b100;
			assign node333 = (inp[7]) ? node335 : 3'b000;
				assign node335 = (inp[0]) ? 3'b000 : node336;
					assign node336 = (inp[10]) ? 3'b000 : node337;
						assign node337 = (inp[1]) ? node359 : node338;
							assign node338 = (inp[11]) ? node352 : node339;
								assign node339 = (inp[8]) ? node345 : node340;
									assign node340 = (inp[3]) ? 3'b000 : node341;
										assign node341 = (inp[2]) ? 3'b000 : 3'b100;
									assign node345 = (inp[2]) ? 3'b100 : node346;
										assign node346 = (inp[3]) ? node348 : 3'b010;
											assign node348 = (inp[5]) ? 3'b100 : 3'b010;
								assign node352 = (inp[2]) ? 3'b000 : node353;
									assign node353 = (inp[3]) ? 3'b000 : node354;
										assign node354 = (inp[8]) ? 3'b100 : 3'b000;
							assign node359 = (inp[4]) ? 3'b000 : node360;
								assign node360 = (inp[11]) ? 3'b000 : node361;
									assign node361 = (inp[3]) ? 3'b000 : node362;
										assign node362 = (inp[2]) ? 3'b000 : node363;
											assign node363 = (inp[8]) ? 3'b100 : 3'b000;
		assign node372 = (inp[9]) ? node900 : node373;
			assign node373 = (inp[0]) ? node593 : node374;
				assign node374 = (inp[7]) ? node518 : node375;
					assign node375 = (inp[10]) ? node439 : node376;
						assign node376 = (inp[1]) ? node400 : node377;
							assign node377 = (inp[8]) ? node389 : node378;
								assign node378 = (inp[11]) ? node384 : node379;
									assign node379 = (inp[3]) ? 3'b011 : node380;
										assign node380 = (inp[2]) ? 3'b011 : 3'b111;
									assign node384 = (inp[3]) ? 3'b101 : node385;
										assign node385 = (inp[2]) ? 3'b101 : 3'b011;
								assign node389 = (inp[11]) ? node391 : 3'b111;
									assign node391 = (inp[2]) ? 3'b011 : node392;
										assign node392 = (inp[3]) ? node394 : 3'b111;
											assign node394 = (inp[4]) ? 3'b011 : node395;
												assign node395 = (inp[5]) ? 3'b011 : 3'b111;
							assign node400 = (inp[8]) ? node416 : node401;
								assign node401 = (inp[11]) ? node407 : node402;
									assign node402 = (inp[2]) ? node404 : 3'b101;
										assign node404 = (inp[3]) ? 3'b001 : 3'b101;
									assign node407 = (inp[2]) ? node413 : node408;
										assign node408 = (inp[3]) ? 3'b001 : node409;
											assign node409 = (inp[4]) ? 3'b001 : 3'b101;
										assign node413 = (inp[4]) ? 3'b110 : 3'b001;
								assign node416 = (inp[11]) ? node426 : node417;
									assign node417 = (inp[5]) ? 3'b011 : node418;
										assign node418 = (inp[3]) ? node422 : node419;
											assign node419 = (inp[2]) ? 3'b011 : 3'b111;
											assign node422 = (inp[2]) ? 3'b101 : 3'b011;
									assign node426 = (inp[3]) ? node434 : node427;
										assign node427 = (inp[2]) ? 3'b101 : node428;
											assign node428 = (inp[4]) ? node430 : 3'b011;
												assign node430 = (inp[5]) ? 3'b101 : 3'b011;
										assign node434 = (inp[5]) ? node436 : 3'b101;
											assign node436 = (inp[4]) ? 3'b001 : 3'b101;
						assign node439 = (inp[1]) ? node471 : node440;
							assign node440 = (inp[11]) ? node456 : node441;
								assign node441 = (inp[8]) ? node449 : node442;
									assign node442 = (inp[2]) ? 3'b001 : node443;
										assign node443 = (inp[3]) ? node445 : 3'b101;
											assign node445 = (inp[5]) ? 3'b001 : 3'b101;
									assign node449 = (inp[2]) ? 3'b101 : node450;
										assign node450 = (inp[3]) ? node452 : 3'b011;
											assign node452 = (inp[4]) ? 3'b101 : 3'b011;
								assign node456 = (inp[8]) ? node464 : node457;
									assign node457 = (inp[2]) ? 3'b110 : node458;
										assign node458 = (inp[3]) ? node460 : 3'b001;
											assign node460 = (inp[5]) ? 3'b110 : 3'b001;
									assign node464 = (inp[2]) ? 3'b001 : node465;
										assign node465 = (inp[3]) ? node467 : 3'b101;
											assign node467 = (inp[4]) ? 3'b001 : 3'b101;
							assign node471 = (inp[8]) ? node495 : node472;
								assign node472 = (inp[11]) ? node482 : node473;
									assign node473 = (inp[2]) ? node477 : node474;
										assign node474 = (inp[4]) ? 3'b110 : 3'b001;
										assign node477 = (inp[4]) ? node479 : 3'b110;
											assign node479 = (inp[5]) ? 3'b110 : 3'b010;
									assign node482 = (inp[2]) ? node490 : node483;
										assign node483 = (inp[3]) ? 3'b010 : node484;
											assign node484 = (inp[4]) ? node486 : 3'b110;
												assign node486 = (inp[5]) ? 3'b010 : 3'b110;
										assign node490 = (inp[4]) ? node492 : 3'b010;
											assign node492 = (inp[3]) ? 3'b100 : 3'b010;
								assign node495 = (inp[11]) ? node509 : node496;
									assign node496 = (inp[5]) ? node502 : node497;
										assign node497 = (inp[3]) ? 3'b001 : node498;
											assign node498 = (inp[2]) ? 3'b001 : 3'b101;
										assign node502 = (inp[3]) ? node504 : 3'b001;
											assign node504 = (inp[4]) ? node506 : 3'b001;
												assign node506 = (inp[2]) ? 3'b110 : 3'b001;
									assign node509 = (inp[3]) ? node513 : node510;
										assign node510 = (inp[2]) ? 3'b110 : 3'b001;
										assign node513 = (inp[2]) ? node515 : 3'b110;
											assign node515 = (inp[4]) ? 3'b010 : 3'b110;
					assign node518 = (inp[10]) ? node544 : node519;
						assign node519 = (inp[8]) ? 3'b111 : node520;
							assign node520 = (inp[1]) ? node522 : 3'b111;
								assign node522 = (inp[11]) ? node532 : node523;
									assign node523 = (inp[2]) ? node525 : 3'b111;
										assign node525 = (inp[5]) ? node527 : 3'b111;
											assign node527 = (inp[3]) ? node529 : 3'b111;
												assign node529 = (inp[4]) ? 3'b011 : 3'b111;
									assign node532 = (inp[2]) ? node536 : node533;
										assign node533 = (inp[3]) ? 3'b011 : 3'b111;
										assign node536 = (inp[4]) ? node538 : 3'b011;
											assign node538 = (inp[3]) ? node540 : 3'b011;
												assign node540 = (inp[5]) ? 3'b101 : 3'b011;
						assign node544 = (inp[1]) ? node564 : node545;
							assign node545 = (inp[8]) ? node557 : node546;
								assign node546 = (inp[11]) ? node550 : node547;
									assign node547 = (inp[2]) ? 3'b011 : 3'b111;
									assign node550 = (inp[2]) ? node552 : 3'b011;
										assign node552 = (inp[3]) ? 3'b101 : node553;
											assign node553 = (inp[4]) ? 3'b101 : 3'b011;
								assign node557 = (inp[11]) ? node559 : 3'b111;
									assign node559 = (inp[2]) ? node561 : 3'b111;
										assign node561 = (inp[3]) ? 3'b011 : 3'b111;
							assign node564 = (inp[8]) ? node576 : node565;
								assign node565 = (inp[11]) ? node571 : node566;
									assign node566 = (inp[2]) ? 3'b101 : node567;
										assign node567 = (inp[3]) ? 3'b101 : 3'b011;
									assign node571 = (inp[2]) ? 3'b001 : node572;
										assign node572 = (inp[3]) ? 3'b001 : 3'b101;
								assign node576 = (inp[11]) ? node586 : node577;
									assign node577 = (inp[2]) ? 3'b011 : node578;
										assign node578 = (inp[3]) ? node580 : 3'b111;
											assign node580 = (inp[5]) ? 3'b011 : node581;
												assign node581 = (inp[4]) ? 3'b011 : 3'b111;
									assign node586 = (inp[2]) ? 3'b101 : node587;
										assign node587 = (inp[5]) ? 3'b101 : node588;
											assign node588 = (inp[4]) ? 3'b101 : 3'b011;
				assign node593 = (inp[7]) ? node737 : node594;
					assign node594 = (inp[10]) ? node670 : node595;
						assign node595 = (inp[1]) ? node625 : node596;
							assign node596 = (inp[11]) ? node610 : node597;
								assign node597 = (inp[8]) ? node605 : node598;
									assign node598 = (inp[2]) ? node600 : 3'b001;
										assign node600 = (inp[4]) ? 3'b110 : node601;
											assign node601 = (inp[3]) ? 3'b110 : 3'b001;
									assign node605 = (inp[2]) ? node607 : 3'b101;
										assign node607 = (inp[3]) ? 3'b001 : 3'b101;
								assign node610 = (inp[8]) ? node620 : node611;
									assign node611 = (inp[2]) ? node613 : 3'b110;
										assign node613 = (inp[5]) ? node615 : 3'b110;
											assign node615 = (inp[3]) ? 3'b010 : node616;
												assign node616 = (inp[4]) ? 3'b010 : 3'b110;
									assign node620 = (inp[3]) ? node622 : 3'b001;
										assign node622 = (inp[2]) ? 3'b110 : 3'b001;
							assign node625 = (inp[8]) ? node641 : node626;
								assign node626 = (inp[11]) ? node632 : node627;
									assign node627 = (inp[2]) ? 3'b010 : node628;
										assign node628 = (inp[4]) ? 3'b010 : 3'b110;
									assign node632 = (inp[2]) ? 3'b100 : node633;
										assign node633 = (inp[4]) ? node635 : 3'b010;
											assign node635 = (inp[5]) ? node637 : 3'b010;
												assign node637 = (inp[3]) ? 3'b100 : 3'b010;
								assign node641 = (inp[11]) ? node655 : node642;
									assign node642 = (inp[2]) ? node648 : node643;
										assign node643 = (inp[3]) ? node645 : 3'b001;
											assign node645 = (inp[4]) ? 3'b110 : 3'b001;
										assign node648 = (inp[4]) ? 3'b110 : node649;
											assign node649 = (inp[3]) ? 3'b110 : node650;
												assign node650 = (inp[5]) ? 3'b110 : 3'b001;
									assign node655 = (inp[2]) ? node663 : node656;
										assign node656 = (inp[4]) ? node658 : 3'b110;
											assign node658 = (inp[5]) ? node660 : 3'b110;
												assign node660 = (inp[3]) ? 3'b010 : 3'b110;
										assign node663 = (inp[4]) ? 3'b010 : node664;
											assign node664 = (inp[5]) ? 3'b010 : node665;
												assign node665 = (inp[3]) ? 3'b010 : 3'b110;
						assign node670 = (inp[8]) ? node700 : node671;
							assign node671 = (inp[1]) ? node687 : node672;
								assign node672 = (inp[11]) ? node682 : node673;
									assign node673 = (inp[5]) ? node675 : 3'b010;
										assign node675 = (inp[3]) ? 3'b100 : node676;
											assign node676 = (inp[2]) ? node678 : 3'b010;
												assign node678 = (inp[4]) ? 3'b100 : 3'b010;
									assign node682 = (inp[3]) ? node684 : 3'b100;
										assign node684 = (inp[2]) ? 3'b000 : 3'b100;
								assign node687 = (inp[11]) ? 3'b000 : node688;
									assign node688 = (inp[2]) ? node696 : node689;
										assign node689 = (inp[5]) ? node691 : 3'b100;
											assign node691 = (inp[4]) ? node693 : 3'b100;
												assign node693 = (inp[3]) ? 3'b000 : 3'b100;
										assign node696 = (inp[3]) ? 3'b000 : 3'b100;
							assign node700 = (inp[1]) ? node722 : node701;
								assign node701 = (inp[11]) ? node707 : node702;
									assign node702 = (inp[3]) ? node704 : 3'b110;
										assign node704 = (inp[2]) ? 3'b010 : 3'b110;
									assign node707 = (inp[2]) ? node715 : node708;
										assign node708 = (inp[5]) ? 3'b010 : node709;
											assign node709 = (inp[3]) ? 3'b010 : node710;
												assign node710 = (inp[4]) ? 3'b010 : 3'b110;
										assign node715 = (inp[3]) ? node717 : 3'b010;
											assign node717 = (inp[5]) ? 3'b100 : node718;
												assign node718 = (inp[4]) ? 3'b100 : 3'b010;
								assign node722 = (inp[11]) ? node732 : node723;
									assign node723 = (inp[2]) ? node725 : 3'b010;
										assign node725 = (inp[5]) ? 3'b100 : node726;
											assign node726 = (inp[3]) ? 3'b100 : node727;
												assign node727 = (inp[4]) ? 3'b100 : 3'b010;
									assign node732 = (inp[2]) ? node734 : 3'b100;
										assign node734 = (inp[3]) ? 3'b000 : 3'b100;
					assign node737 = (inp[10]) ? node819 : node738;
						assign node738 = (inp[1]) ? node786 : node739;
							assign node739 = (inp[8]) ? node765 : node740;
								assign node740 = (inp[11]) ? node752 : node741;
									assign node741 = (inp[3]) ? node749 : node742;
										assign node742 = (inp[2]) ? 3'b011 : node743;
											assign node743 = (inp[5]) ? 3'b011 : node744;
												assign node744 = (inp[4]) ? 3'b011 : 3'b111;
										assign node749 = (inp[2]) ? 3'b101 : 3'b011;
									assign node752 = (inp[4]) ? 3'b101 : node753;
										assign node753 = (inp[5]) ? node759 : node754;
											assign node754 = (inp[3]) ? 3'b101 : node755;
												assign node755 = (inp[2]) ? 3'b101 : 3'b011;
											assign node759 = (inp[2]) ? node761 : 3'b101;
												assign node761 = (inp[3]) ? 3'b001 : 3'b101;
								assign node765 = (inp[11]) ? node775 : node766;
									assign node766 = (inp[3]) ? node768 : 3'b111;
										assign node768 = (inp[2]) ? node770 : 3'b111;
											assign node770 = (inp[4]) ? 3'b011 : node771;
												assign node771 = (inp[5]) ? 3'b011 : 3'b111;
									assign node775 = (inp[2]) ? node781 : node776;
										assign node776 = (inp[4]) ? 3'b011 : node777;
											assign node777 = (inp[3]) ? 3'b011 : 3'b111;
										assign node781 = (inp[4]) ? node783 : 3'b011;
											assign node783 = (inp[3]) ? 3'b101 : 3'b011;
							assign node786 = (inp[11]) ? node802 : node787;
								assign node787 = (inp[8]) ? node795 : node788;
									assign node788 = (inp[2]) ? node790 : 3'b101;
										assign node790 = (inp[3]) ? 3'b001 : node791;
											assign node791 = (inp[4]) ? 3'b001 : 3'b101;
									assign node795 = (inp[2]) ? node797 : 3'b011;
										assign node797 = (inp[5]) ? node799 : 3'b101;
											assign node799 = (inp[4]) ? 3'b101 : 3'b011;
								assign node802 = (inp[8]) ? node810 : node803;
									assign node803 = (inp[2]) ? node805 : 3'b001;
										assign node805 = (inp[3]) ? 3'b110 : node806;
											assign node806 = (inp[4]) ? 3'b110 : 3'b001;
									assign node810 = (inp[2]) ? node812 : 3'b101;
										assign node812 = (inp[3]) ? 3'b001 : node813;
											assign node813 = (inp[4]) ? node815 : 3'b101;
												assign node815 = (inp[5]) ? 3'b001 : 3'b101;
						assign node819 = (inp[1]) ? node871 : node820;
							assign node820 = (inp[4]) ? node844 : node821;
								assign node821 = (inp[8]) ? node833 : node822;
									assign node822 = (inp[11]) ? node830 : node823;
										assign node823 = (inp[5]) ? 3'b001 : node824;
											assign node824 = (inp[2]) ? 3'b001 : node825;
												assign node825 = (inp[3]) ? 3'b001 : 3'b101;
										assign node830 = (inp[3]) ? 3'b010 : 3'b001;
									assign node833 = (inp[11]) ? node839 : node834;
										assign node834 = (inp[2]) ? 3'b101 : node835;
											assign node835 = (inp[3]) ? 3'b101 : 3'b011;
										assign node839 = (inp[2]) ? 3'b001 : node840;
											assign node840 = (inp[3]) ? 3'b001 : 3'b101;
								assign node844 = (inp[11]) ? node856 : node845;
									assign node845 = (inp[8]) ? node851 : node846;
										assign node846 = (inp[3]) ? node848 : 3'b001;
											assign node848 = (inp[2]) ? 3'b110 : 3'b001;
										assign node851 = (inp[5]) ? 3'b101 : node852;
											assign node852 = (inp[3]) ? 3'b001 : 3'b101;
									assign node856 = (inp[8]) ? node862 : node857;
										assign node857 = (inp[3]) ? node859 : 3'b110;
											assign node859 = (inp[2]) ? 3'b010 : 3'b110;
										assign node862 = (inp[2]) ? node868 : node863;
											assign node863 = (inp[3]) ? 3'b001 : node864;
												assign node864 = (inp[5]) ? 3'b001 : 3'b101;
											assign node868 = (inp[3]) ? 3'b110 : 3'b011;
							assign node871 = (inp[8]) ? node887 : node872;
								assign node872 = (inp[11]) ? node880 : node873;
									assign node873 = (inp[2]) ? node875 : 3'b110;
										assign node875 = (inp[4]) ? 3'b010 : node876;
											assign node876 = (inp[3]) ? 3'b010 : 3'b110;
									assign node880 = (inp[2]) ? node882 : 3'b010;
										assign node882 = (inp[3]) ? 3'b100 : node883;
											assign node883 = (inp[4]) ? 3'b100 : 3'b010;
								assign node887 = (inp[11]) ? node895 : node888;
									assign node888 = (inp[2]) ? node890 : 3'b001;
										assign node890 = (inp[3]) ? 3'b110 : node891;
											assign node891 = (inp[5]) ? 3'b110 : 3'b001;
									assign node895 = (inp[2]) ? node897 : 3'b110;
										assign node897 = (inp[3]) ? 3'b010 : 3'b110;
			assign node900 = (inp[0]) ? node1140 : node901;
				assign node901 = (inp[7]) ? node1009 : node902;
					assign node902 = (inp[10]) ? node962 : node903;
						assign node903 = (inp[1]) ? node939 : node904;
							assign node904 = (inp[8]) ? node920 : node905;
								assign node905 = (inp[11]) ? node913 : node906;
									assign node906 = (inp[2]) ? 3'b010 : node907;
										assign node907 = (inp[4]) ? node909 : 3'b110;
											assign node909 = (inp[3]) ? 3'b010 : 3'b110;
									assign node913 = (inp[2]) ? 3'b100 : node914;
										assign node914 = (inp[4]) ? node916 : 3'b010;
											assign node916 = (inp[3]) ? 3'b100 : 3'b010;
								assign node920 = (inp[2]) ? node930 : node921;
									assign node921 = (inp[11]) ? node923 : 3'b001;
										assign node923 = (inp[3]) ? node925 : 3'b110;
											assign node925 = (inp[5]) ? node927 : 3'b110;
												assign node927 = (inp[4]) ? 3'b010 : 3'b110;
									assign node930 = (inp[11]) ? node932 : 3'b110;
										assign node932 = (inp[3]) ? 3'b010 : node933;
											assign node933 = (inp[5]) ? 3'b010 : node934;
												assign node934 = (inp[4]) ? 3'b010 : 3'b110;
							assign node939 = (inp[11]) ? node951 : node940;
								assign node940 = (inp[8]) ? node946 : node941;
									assign node941 = (inp[2]) ? 3'b100 : node942;
										assign node942 = (inp[3]) ? 3'b100 : 3'b010;
									assign node946 = (inp[2]) ? 3'b010 : node947;
										assign node947 = (inp[3]) ? 3'b010 : 3'b110;
								assign node951 = (inp[8]) ? node957 : node952;
									assign node952 = (inp[3]) ? 3'b000 : node953;
										assign node953 = (inp[2]) ? 3'b000 : 3'b100;
									assign node957 = (inp[2]) ? 3'b100 : node958;
										assign node958 = (inp[3]) ? 3'b100 : 3'b010;
						assign node962 = (inp[1]) ? node998 : node963;
							assign node963 = (inp[8]) ? node975 : node964;
								assign node964 = (inp[11]) ? 3'b000 : node965;
									assign node965 = (inp[2]) ? 3'b000 : node966;
										assign node966 = (inp[4]) ? node968 : 3'b100;
											assign node968 = (inp[3]) ? node970 : 3'b100;
												assign node970 = (inp[5]) ? 3'b000 : 3'b100;
								assign node975 = (inp[11]) ? node991 : node976;
									assign node976 = (inp[2]) ? node984 : node977;
										assign node977 = (inp[4]) ? node979 : 3'b010;
											assign node979 = (inp[3]) ? node981 : 3'b010;
												assign node981 = (inp[5]) ? 3'b100 : 3'b010;
										assign node984 = (inp[4]) ? 3'b100 : node985;
											assign node985 = (inp[3]) ? 3'b100 : node986;
												assign node986 = (inp[5]) ? 3'b100 : 3'b010;
									assign node991 = (inp[2]) ? node993 : 3'b100;
										assign node993 = (inp[3]) ? 3'b000 : node994;
											assign node994 = (inp[4]) ? 3'b000 : 3'b100;
							assign node998 = (inp[2]) ? 3'b000 : node999;
								assign node999 = (inp[8]) ? node1001 : 3'b000;
									assign node1001 = (inp[11]) ? 3'b000 : node1002;
										assign node1002 = (inp[4]) ? node1004 : 3'b100;
											assign node1004 = (inp[3]) ? 3'b000 : 3'b100;
					assign node1009 = (inp[10]) ? node1075 : node1010;
						assign node1010 = (inp[1]) ? node1042 : node1011;
							assign node1011 = (inp[11]) ? node1027 : node1012;
								assign node1012 = (inp[8]) ? node1022 : node1013;
									assign node1013 = (inp[2]) ? node1019 : node1014;
										assign node1014 = (inp[3]) ? node1016 : 3'b101;
											assign node1016 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1019 = (inp[4]) ? 3'b001 : 3'b101;
									assign node1022 = (inp[2]) ? node1024 : 3'b011;
										assign node1024 = (inp[5]) ? 3'b101 : 3'b011;
								assign node1027 = (inp[8]) ? node1035 : node1028;
									assign node1028 = (inp[2]) ? node1030 : 3'b001;
										assign node1030 = (inp[3]) ? 3'b110 : node1031;
											assign node1031 = (inp[4]) ? 3'b110 : 3'b001;
									assign node1035 = (inp[2]) ? node1037 : 3'b101;
										assign node1037 = (inp[4]) ? 3'b001 : node1038;
											assign node1038 = (inp[3]) ? 3'b001 : 3'b101;
							assign node1042 = (inp[8]) ? node1060 : node1043;
								assign node1043 = (inp[11]) ? node1053 : node1044;
									assign node1044 = (inp[2]) ? 3'b110 : node1045;
										assign node1045 = (inp[3]) ? node1047 : 3'b001;
											assign node1047 = (inp[4]) ? 3'b110 : node1048;
												assign node1048 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1053 = (inp[2]) ? 3'b010 : node1054;
										assign node1054 = (inp[3]) ? node1056 : 3'b110;
											assign node1056 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1060 = (inp[11]) ? node1068 : node1061;
									assign node1061 = (inp[2]) ? 3'b001 : node1062;
										assign node1062 = (inp[4]) ? node1064 : 3'b101;
											assign node1064 = (inp[3]) ? 3'b001 : 3'b101;
									assign node1068 = (inp[2]) ? 3'b110 : node1069;
										assign node1069 = (inp[3]) ? node1071 : 3'b001;
											assign node1071 = (inp[4]) ? 3'b110 : 3'b001;
						assign node1075 = (inp[1]) ? node1109 : node1076;
							assign node1076 = (inp[11]) ? node1094 : node1077;
								assign node1077 = (inp[8]) ? node1085 : node1078;
									assign node1078 = (inp[2]) ? node1080 : 3'b110;
										assign node1080 = (inp[4]) ? 3'b010 : node1081;
											assign node1081 = (inp[3]) ? 3'b010 : 3'b110;
									assign node1085 = (inp[2]) ? node1087 : 3'b001;
										assign node1087 = (inp[3]) ? 3'b110 : node1088;
											assign node1088 = (inp[5]) ? node1090 : 3'b001;
												assign node1090 = (inp[4]) ? 3'b110 : 3'b001;
								assign node1094 = (inp[8]) ? node1100 : node1095;
									assign node1095 = (inp[3]) ? node1097 : 3'b010;
										assign node1097 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1100 = (inp[2]) ? node1102 : 3'b110;
										assign node1102 = (inp[3]) ? 3'b010 : node1103;
											assign node1103 = (inp[4]) ? node1105 : 3'b110;
												assign node1105 = (inp[5]) ? 3'b010 : 3'b110;
							assign node1109 = (inp[8]) ? node1125 : node1110;
								assign node1110 = (inp[11]) ? node1118 : node1111;
									assign node1111 = (inp[2]) ? 3'b100 : node1112;
										assign node1112 = (inp[4]) ? node1114 : 3'b010;
											assign node1114 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1118 = (inp[2]) ? 3'b000 : node1119;
										assign node1119 = (inp[3]) ? node1121 : 3'b100;
											assign node1121 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1125 = (inp[11]) ? node1133 : node1126;
									assign node1126 = (inp[2]) ? 3'b010 : node1127;
										assign node1127 = (inp[3]) ? node1129 : 3'b110;
											assign node1129 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1133 = (inp[2]) ? 3'b100 : node1134;
										assign node1134 = (inp[5]) ? node1136 : 3'b010;
											assign node1136 = (inp[3]) ? 3'b100 : 3'b010;
				assign node1140 = (inp[7]) ? node1166 : node1141;
					assign node1141 = (inp[10]) ? 3'b000 : node1142;
						assign node1142 = (inp[8]) ? node1144 : 3'b000;
							assign node1144 = (inp[1]) ? 3'b000 : node1145;
								assign node1145 = (inp[11]) ? node1157 : node1146;
									assign node1146 = (inp[2]) ? node1154 : node1147;
										assign node1147 = (inp[5]) ? 3'b100 : node1148;
											assign node1148 = (inp[4]) ? 3'b100 : node1149;
												assign node1149 = (inp[3]) ? 3'b100 : 3'b010;
										assign node1154 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1157 = (inp[3]) ? 3'b000 : node1158;
										assign node1158 = (inp[4]) ? 3'b000 : node1159;
											assign node1159 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1166 = (inp[10]) ? node1244 : node1167;
						assign node1167 = (inp[1]) ? node1217 : node1168;
							assign node1168 = (inp[11]) ? node1188 : node1169;
								assign node1169 = (inp[8]) ? node1177 : node1170;
									assign node1170 = (inp[4]) ? 3'b010 : node1171;
										assign node1171 = (inp[3]) ? 3'b010 : node1172;
											assign node1172 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1177 = (inp[3]) ? node1185 : node1178;
										assign node1178 = (inp[2]) ? 3'b110 : node1179;
											assign node1179 = (inp[5]) ? node1181 : 3'b001;
												assign node1181 = (inp[4]) ? 3'b110 : 3'b001;
										assign node1185 = (inp[2]) ? 3'b010 : 3'b110;
								assign node1188 = (inp[8]) ? node1202 : node1189;
									assign node1189 = (inp[3]) ? node1197 : node1190;
										assign node1190 = (inp[2]) ? 3'b100 : node1191;
											assign node1191 = (inp[5]) ? node1193 : 3'b010;
												assign node1193 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1197 = (inp[2]) ? node1199 : 3'b100;
											assign node1199 = (inp[4]) ? 3'b000 : 3'b100;
									assign node1202 = (inp[2]) ? node1210 : node1203;
										assign node1203 = (inp[3]) ? 3'b010 : node1204;
											assign node1204 = (inp[5]) ? node1206 : 3'b110;
												assign node1206 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1210 = (inp[3]) ? node1212 : 3'b010;
											assign node1212 = (inp[4]) ? 3'b100 : node1213;
												assign node1213 = (inp[5]) ? 3'b000 : 3'b010;
							assign node1217 = (inp[8]) ? node1229 : node1218;
								assign node1218 = (inp[11]) ? 3'b000 : node1219;
									assign node1219 = (inp[2]) ? node1221 : 3'b100;
										assign node1221 = (inp[3]) ? 3'b000 : node1222;
											assign node1222 = (inp[4]) ? node1224 : 3'b100;
												assign node1224 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1229 = (inp[11]) ? node1235 : node1230;
									assign node1230 = (inp[3]) ? node1232 : 3'b010;
										assign node1232 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1235 = (inp[2]) ? node1241 : node1236;
										assign node1236 = (inp[3]) ? 3'b100 : node1237;
											assign node1237 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1241 = (inp[3]) ? 3'b000 : 3'b100;
						assign node1244 = (inp[8]) ? node1246 : 3'b000;
							assign node1246 = (inp[1]) ? 3'b000 : node1247;
								assign node1247 = (inp[11]) ? node1257 : node1248;
									assign node1248 = (inp[2]) ? 3'b100 : node1249;
										assign node1249 = (inp[3]) ? 3'b100 : node1250;
											assign node1250 = (inp[5]) ? node1252 : 3'b011;
												assign node1252 = (inp[4]) ? 3'b010 : 3'b011;
									assign node1257 = (inp[3]) ? 3'b000 : node1258;
										assign node1258 = (inp[2]) ? 3'b000 : 3'b100;

endmodule