module dtc_split5_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node976;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1128;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1162;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1259;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1327;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1335;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1347;
	wire [3-1:0] node1349;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1357;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1382;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1394;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1409;
	wire [3-1:0] node1411;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1453;
	wire [3-1:0] node1454;
	wire [3-1:0] node1456;
	wire [3-1:0] node1458;
	wire [3-1:0] node1461;
	wire [3-1:0] node1462;
	wire [3-1:0] node1463;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1481;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1498;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1525;
	wire [3-1:0] node1526;
	wire [3-1:0] node1528;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1548;
	wire [3-1:0] node1550;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1559;
	wire [3-1:0] node1560;
	wire [3-1:0] node1564;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1567;
	wire [3-1:0] node1571;
	wire [3-1:0] node1572;
	wire [3-1:0] node1576;
	wire [3-1:0] node1578;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1583;
	wire [3-1:0] node1585;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1594;
	wire [3-1:0] node1596;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1602;
	wire [3-1:0] node1605;
	wire [3-1:0] node1606;
	wire [3-1:0] node1608;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1614;
	wire [3-1:0] node1615;
	wire [3-1:0] node1616;
	wire [3-1:0] node1617;
	wire [3-1:0] node1621;
	wire [3-1:0] node1624;
	wire [3-1:0] node1625;
	wire [3-1:0] node1626;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1634;
	wire [3-1:0] node1637;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1640;
	wire [3-1:0] node1643;
	wire [3-1:0] node1646;
	wire [3-1:0] node1648;
	wire [3-1:0] node1651;
	wire [3-1:0] node1653;
	wire [3-1:0] node1656;
	wire [3-1:0] node1657;
	wire [3-1:0] node1660;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1666;
	wire [3-1:0] node1669;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1678;
	wire [3-1:0] node1681;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1687;
	wire [3-1:0] node1690;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1695;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1705;
	wire [3-1:0] node1706;
	wire [3-1:0] node1710;
	wire [3-1:0] node1711;
	wire [3-1:0] node1712;
	wire [3-1:0] node1713;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1718;
	wire [3-1:0] node1721;
	wire [3-1:0] node1722;
	wire [3-1:0] node1723;
	wire [3-1:0] node1724;
	wire [3-1:0] node1728;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1736;
	wire [3-1:0] node1739;
	wire [3-1:0] node1740;
	wire [3-1:0] node1743;
	wire [3-1:0] node1746;
	wire [3-1:0] node1747;
	wire [3-1:0] node1750;
	wire [3-1:0] node1753;
	wire [3-1:0] node1754;
	wire [3-1:0] node1755;
	wire [3-1:0] node1756;
	wire [3-1:0] node1757;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1767;
	wire [3-1:0] node1768;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1783;
	wire [3-1:0] node1787;
	wire [3-1:0] node1788;
	wire [3-1:0] node1792;
	wire [3-1:0] node1793;

	assign outp = (inp[5]) ? node1028 : node1;
		assign node1 = (inp[8]) ? node631 : node2;
			assign node2 = (inp[6]) ? node326 : node3;
				assign node3 = (inp[4]) ? node165 : node4;
					assign node4 = (inp[0]) ? node92 : node5;
						assign node5 = (inp[9]) ? node45 : node6;
							assign node6 = (inp[7]) ? node20 : node7;
								assign node7 = (inp[10]) ? node11 : node8;
									assign node8 = (inp[3]) ? 3'b010 : 3'b000;
									assign node11 = (inp[3]) ? node17 : node12;
										assign node12 = (inp[2]) ? 3'b011 : node13;
											assign node13 = (inp[11]) ? 3'b011 : 3'b010;
										assign node17 = (inp[11]) ? 3'b000 : 3'b001;
								assign node20 = (inp[11]) ? node32 : node21;
									assign node21 = (inp[10]) ? node27 : node22;
										assign node22 = (inp[1]) ? node24 : 3'b011;
											assign node24 = (inp[2]) ? 3'b010 : 3'b011;
										assign node27 = (inp[2]) ? 3'b011 : node28;
											assign node28 = (inp[3]) ? 3'b000 : 3'b010;
									assign node32 = (inp[2]) ? node38 : node33;
										assign node33 = (inp[3]) ? 3'b011 : node34;
											assign node34 = (inp[1]) ? 3'b011 : 3'b010;
										assign node38 = (inp[1]) ? node42 : node39;
											assign node39 = (inp[10]) ? 3'b000 : 3'b000;
											assign node42 = (inp[3]) ? 3'b001 : 3'b011;
							assign node45 = (inp[7]) ? node73 : node46;
								assign node46 = (inp[1]) ? node58 : node47;
									assign node47 = (inp[11]) ? node53 : node48;
										assign node48 = (inp[10]) ? 3'b011 : node49;
											assign node49 = (inp[3]) ? 3'b011 : 3'b001;
										assign node53 = (inp[10]) ? 3'b000 : node54;
											assign node54 = (inp[3]) ? 3'b011 : 3'b001;
									assign node58 = (inp[11]) ? node66 : node59;
										assign node59 = (inp[2]) ? node63 : node60;
											assign node60 = (inp[3]) ? 3'b011 : 3'b001;
											assign node63 = (inp[3]) ? 3'b010 : 3'b000;
										assign node66 = (inp[2]) ? node70 : node67;
											assign node67 = (inp[10]) ? 3'b010 : 3'b011;
											assign node70 = (inp[3]) ? 3'b001 : 3'b011;
								assign node73 = (inp[11]) ? node81 : node74;
									assign node74 = (inp[2]) ? 3'b001 : node75;
										assign node75 = (inp[1]) ? 3'b001 : node76;
											assign node76 = (inp[10]) ? 3'b000 : 3'b010;
									assign node81 = (inp[3]) ? node89 : node82;
										assign node82 = (inp[10]) ? node86 : node83;
											assign node83 = (inp[2]) ? 3'b010 : 3'b011;
											assign node86 = (inp[1]) ? 3'b000 : 3'b001;
										assign node89 = (inp[10]) ? 3'b010 : 3'b000;
						assign node92 = (inp[11]) ? node132 : node93;
							assign node93 = (inp[9]) ? node113 : node94;
								assign node94 = (inp[2]) ? node100 : node95;
									assign node95 = (inp[3]) ? 3'b000 : node96;
										assign node96 = (inp[10]) ? 3'b011 : 3'b001;
									assign node100 = (inp[1]) ? node108 : node101;
										assign node101 = (inp[3]) ? node105 : node102;
											assign node102 = (inp[10]) ? 3'b011 : 3'b001;
											assign node105 = (inp[10]) ? 3'b000 : 3'b010;
										assign node108 = (inp[3]) ? 3'b001 : node109;
											assign node109 = (inp[10]) ? 3'b010 : 3'b000;
								assign node113 = (inp[3]) ? node121 : node114;
									assign node114 = (inp[10]) ? node116 : 3'b000;
										assign node116 = (inp[2]) ? node118 : 3'b010;
											assign node118 = (inp[1]) ? 3'b011 : 3'b010;
									assign node121 = (inp[10]) ? node127 : node122;
										assign node122 = (inp[2]) ? node124 : 3'b011;
											assign node124 = (inp[1]) ? 3'b010 : 3'b010;
										assign node127 = (inp[2]) ? 3'b001 : node128;
											assign node128 = (inp[7]) ? 3'b001 : 3'b000;
							assign node132 = (inp[2]) ? node148 : node133;
								assign node133 = (inp[3]) ? node139 : node134;
									assign node134 = (inp[1]) ? 3'b010 : node135;
										assign node135 = (inp[10]) ? 3'b000 : 3'b010;
									assign node139 = (inp[7]) ? node143 : node140;
										assign node140 = (inp[10]) ? 3'b000 : 3'b010;
										assign node143 = (inp[10]) ? node145 : 3'b000;
											assign node145 = (inp[9]) ? 3'b011 : 3'b010;
								assign node148 = (inp[7]) ? node156 : node149;
									assign node149 = (inp[10]) ? node153 : node150;
										assign node150 = (inp[3]) ? 3'b011 : 3'b001;
										assign node153 = (inp[3]) ? 3'b000 : 3'b011;
									assign node156 = (inp[1]) ? node160 : node157;
										assign node157 = (inp[9]) ? 3'b000 : 3'b001;
										assign node160 = (inp[9]) ? 3'b010 : node161;
											assign node161 = (inp[3]) ? 3'b000 : 3'b000;
					assign node165 = (inp[3]) ? node249 : node166;
						assign node166 = (inp[7]) ? node216 : node167;
							assign node167 = (inp[1]) ? node193 : node168;
								assign node168 = (inp[9]) ? node178 : node169;
									assign node169 = (inp[0]) ? node171 : 3'b110;
										assign node171 = (inp[2]) ? node175 : node172;
											assign node172 = (inp[10]) ? 3'b111 : 3'b101;
											assign node175 = (inp[11]) ? 3'b100 : 3'b110;
									assign node178 = (inp[11]) ? node186 : node179;
										assign node179 = (inp[10]) ? node183 : node180;
											assign node180 = (inp[2]) ? 3'b100 : 3'b101;
											assign node183 = (inp[2]) ? 3'b110 : 3'b110;
										assign node186 = (inp[10]) ? node190 : node187;
											assign node187 = (inp[0]) ? 3'b111 : 3'b110;
											assign node190 = (inp[2]) ? 3'b100 : 3'b100;
								assign node193 = (inp[2]) ? node205 : node194;
									assign node194 = (inp[0]) ? node202 : node195;
										assign node195 = (inp[9]) ? node199 : node196;
											assign node196 = (inp[11]) ? 3'b100 : 3'b100;
											assign node199 = (inp[11]) ? 3'b100 : 3'b100;
										assign node202 = (inp[9]) ? 3'b111 : 3'b101;
									assign node205 = (inp[0]) ? node211 : node206;
										assign node206 = (inp[11]) ? node208 : 3'b101;
											assign node208 = (inp[10]) ? 3'b101 : 3'b111;
										assign node211 = (inp[9]) ? 3'b100 : node212;
											assign node212 = (inp[10]) ? 3'b110 : 3'b100;
							assign node216 = (inp[2]) ? node228 : node217;
								assign node217 = (inp[0]) ? node223 : node218;
									assign node218 = (inp[10]) ? node220 : 3'b100;
										assign node220 = (inp[11]) ? 3'b100 : 3'b110;
									assign node223 = (inp[10]) ? node225 : 3'b101;
										assign node225 = (inp[11]) ? 3'b101 : 3'b111;
								assign node228 = (inp[0]) ? node242 : node229;
									assign node229 = (inp[9]) ? node235 : node230;
										assign node230 = (inp[10]) ? 3'b101 : node231;
											assign node231 = (inp[11]) ? 3'b110 : 3'b101;
										assign node235 = (inp[10]) ? node239 : node236;
											assign node236 = (inp[11]) ? 3'b111 : 3'b101;
											assign node239 = (inp[11]) ? 3'b101 : 3'b111;
									assign node242 = (inp[10]) ? 3'b100 : node243;
										assign node243 = (inp[1]) ? 3'b111 : node244;
											assign node244 = (inp[11]) ? 3'b110 : 3'b100;
						assign node249 = (inp[7]) ? node287 : node250;
							assign node250 = (inp[11]) ? node270 : node251;
								assign node251 = (inp[10]) ? node261 : node252;
									assign node252 = (inp[2]) ? node254 : 3'b101;
										assign node254 = (inp[0]) ? node258 : node255;
											assign node255 = (inp[1]) ? 3'b100 : 3'b101;
											assign node258 = (inp[1]) ? 3'b101 : 3'b100;
									assign node261 = (inp[0]) ? node263 : 3'b110;
										assign node263 = (inp[1]) ? node267 : node264;
											assign node264 = (inp[2]) ? 3'b110 : 3'b111;
											assign node267 = (inp[2]) ? 3'b111 : 3'b110;
								assign node270 = (inp[10]) ? node284 : node271;
									assign node271 = (inp[2]) ? node279 : node272;
										assign node272 = (inp[9]) ? node276 : node273;
											assign node273 = (inp[1]) ? 3'b110 : 3'b110;
											assign node276 = (inp[0]) ? 3'b110 : 3'b110;
										assign node279 = (inp[1]) ? 3'b111 : node280;
											assign node280 = (inp[0]) ? 3'b110 : 3'b111;
									assign node284 = (inp[1]) ? 3'b101 : 3'b100;
							assign node287 = (inp[9]) ? node305 : node288;
								assign node288 = (inp[11]) ? node298 : node289;
									assign node289 = (inp[10]) ? node293 : node290;
										assign node290 = (inp[1]) ? 3'b101 : 3'b100;
										assign node293 = (inp[1]) ? 3'b110 : node294;
											assign node294 = (inp[0]) ? 3'b110 : 3'b111;
									assign node298 = (inp[10]) ? node300 : 3'b110;
										assign node300 = (inp[2]) ? node302 : 3'b100;
											assign node302 = (inp[0]) ? 3'b100 : 3'b100;
								assign node305 = (inp[1]) ? node315 : node306;
									assign node306 = (inp[11]) ? node312 : node307;
										assign node307 = (inp[10]) ? node309 : 3'b100;
											assign node309 = (inp[2]) ? 3'b111 : 3'b110;
										assign node312 = (inp[0]) ? 3'b101 : 3'b111;
									assign node315 = (inp[10]) ? node321 : node316;
										assign node316 = (inp[11]) ? node318 : 3'b100;
											assign node318 = (inp[0]) ? 3'b110 : 3'b110;
										assign node321 = (inp[0]) ? 3'b110 : node322;
											assign node322 = (inp[2]) ? 3'b111 : 3'b110;
				assign node326 = (inp[11]) ? node472 : node327;
					assign node327 = (inp[10]) ? node399 : node328;
						assign node328 = (inp[4]) ? node368 : node329;
							assign node329 = (inp[7]) ? node351 : node330;
								assign node330 = (inp[3]) ? node344 : node331;
									assign node331 = (inp[1]) ? node337 : node332;
										assign node332 = (inp[2]) ? 3'b101 : node333;
											assign node333 = (inp[0]) ? 3'b101 : 3'b100;
										assign node337 = (inp[9]) ? node341 : node338;
											assign node338 = (inp[0]) ? 3'b100 : 3'b100;
											assign node341 = (inp[2]) ? 3'b100 : 3'b100;
									assign node344 = (inp[9]) ? node346 : 3'b111;
										assign node346 = (inp[1]) ? 3'b110 : node347;
											assign node347 = (inp[0]) ? 3'b110 : 3'b111;
								assign node351 = (inp[3]) ? node361 : node352;
									assign node352 = (inp[2]) ? node356 : node353;
										assign node353 = (inp[9]) ? 3'b110 : 3'b111;
										assign node356 = (inp[9]) ? node358 : 3'b110;
											assign node358 = (inp[1]) ? 3'b111 : 3'b110;
									assign node361 = (inp[9]) ? 3'b101 : node362;
										assign node362 = (inp[0]) ? 3'b100 : node363;
											assign node363 = (inp[2]) ? 3'b100 : 3'b101;
							assign node368 = (inp[2]) ? node380 : node369;
								assign node369 = (inp[0]) ? node371 : 3'b100;
									assign node371 = (inp[1]) ? node373 : 3'b101;
										assign node373 = (inp[3]) ? node377 : node374;
											assign node374 = (inp[7]) ? 3'b101 : 3'b100;
											assign node377 = (inp[7]) ? 3'b100 : 3'b101;
								assign node380 = (inp[0]) ? node390 : node381;
									assign node381 = (inp[1]) ? node383 : 3'b101;
										assign node383 = (inp[9]) ? node387 : node384;
											assign node384 = (inp[3]) ? 3'b101 : 3'b100;
											assign node387 = (inp[7]) ? 3'b100 : 3'b101;
									assign node390 = (inp[1]) ? node392 : 3'b100;
										assign node392 = (inp[3]) ? node396 : node393;
											assign node393 = (inp[7]) ? 3'b100 : 3'b101;
											assign node396 = (inp[7]) ? 3'b101 : 3'b100;
						assign node399 = (inp[4]) ? node439 : node400;
							assign node400 = (inp[2]) ? node420 : node401;
								assign node401 = (inp[3]) ? node409 : node402;
									assign node402 = (inp[7]) ? 3'b101 : node403;
										assign node403 = (inp[9]) ? 3'b111 : node404;
											assign node404 = (inp[0]) ? 3'b111 : 3'b110;
									assign node409 = (inp[7]) ? node415 : node410;
										assign node410 = (inp[0]) ? node412 : 3'b100;
											assign node412 = (inp[1]) ? 3'b100 : 3'b101;
										assign node415 = (inp[1]) ? 3'b110 : node416;
											assign node416 = (inp[9]) ? 3'b110 : 3'b111;
								assign node420 = (inp[3]) ? node428 : node421;
									assign node421 = (inp[7]) ? 3'b100 : node422;
										assign node422 = (inp[1]) ? node424 : 3'b110;
											assign node424 = (inp[9]) ? 3'b111 : 3'b110;
									assign node428 = (inp[7]) ? node434 : node429;
										assign node429 = (inp[1]) ? 3'b101 : node430;
											assign node430 = (inp[0]) ? 3'b100 : 3'b101;
										assign node434 = (inp[0]) ? 3'b111 : node435;
											assign node435 = (inp[1]) ? 3'b110 : 3'b111;
							assign node439 = (inp[9]) ? node459 : node440;
								assign node440 = (inp[3]) ? node450 : node441;
									assign node441 = (inp[7]) ? 3'b110 : node442;
										assign node442 = (inp[0]) ? node446 : node443;
											assign node443 = (inp[2]) ? 3'b111 : 3'b110;
											assign node446 = (inp[2]) ? 3'b110 : 3'b111;
									assign node450 = (inp[2]) ? node456 : node451;
										assign node451 = (inp[0]) ? node453 : 3'b110;
											assign node453 = (inp[1]) ? 3'b111 : 3'b110;
										assign node456 = (inp[0]) ? 3'b110 : 3'b111;
								assign node459 = (inp[3]) ? node461 : 3'b111;
									assign node461 = (inp[2]) ? node467 : node462;
										assign node462 = (inp[7]) ? node464 : 3'b111;
											assign node464 = (inp[0]) ? 3'b111 : 3'b110;
										assign node467 = (inp[1]) ? 3'b110 : node468;
											assign node468 = (inp[0]) ? 3'b111 : 3'b110;
					assign node472 = (inp[10]) ? node550 : node473;
						assign node473 = (inp[3]) ? node513 : node474;
							assign node474 = (inp[4]) ? node494 : node475;
								assign node475 = (inp[0]) ? node485 : node476;
									assign node476 = (inp[1]) ? 3'b100 : node477;
										assign node477 = (inp[9]) ? node481 : node478;
											assign node478 = (inp[7]) ? 3'b101 : 3'b100;
											assign node481 = (inp[7]) ? 3'b100 : 3'b101;
									assign node485 = (inp[7]) ? node491 : node486;
										assign node486 = (inp[9]) ? 3'b100 : node487;
											assign node487 = (inp[2]) ? 3'b101 : 3'b100;
										assign node491 = (inp[9]) ? 3'b101 : 3'b100;
								assign node494 = (inp[9]) ? node502 : node495;
									assign node495 = (inp[2]) ? 3'b110 : node496;
										assign node496 = (inp[0]) ? node498 : 3'b110;
											assign node498 = (inp[7]) ? 3'b110 : 3'b110;
									assign node502 = (inp[2]) ? node508 : node503;
										assign node503 = (inp[7]) ? node505 : 3'b110;
											assign node505 = (inp[1]) ? 3'b110 : 3'b110;
										assign node508 = (inp[7]) ? node510 : 3'b111;
											assign node510 = (inp[1]) ? 3'b110 : 3'b110;
							assign node513 = (inp[7]) ? node535 : node514;
								assign node514 = (inp[4]) ? node528 : node515;
									assign node515 = (inp[2]) ? node521 : node516;
										assign node516 = (inp[1]) ? node518 : 3'b110;
											assign node518 = (inp[9]) ? 3'b110 : 3'b110;
										assign node521 = (inp[1]) ? node525 : node522;
											assign node522 = (inp[0]) ? 3'b111 : 3'b110;
											assign node525 = (inp[0]) ? 3'b110 : 3'b110;
									assign node528 = (inp[2]) ? node532 : node529;
										assign node529 = (inp[0]) ? 3'b111 : 3'b110;
										assign node532 = (inp[0]) ? 3'b110 : 3'b111;
								assign node535 = (inp[0]) ? node543 : node536;
									assign node536 = (inp[9]) ? 3'b111 : node537;
										assign node537 = (inp[1]) ? node539 : 3'b110;
											assign node539 = (inp[2]) ? 3'b110 : 3'b110;
									assign node543 = (inp[9]) ? 3'b110 : node544;
										assign node544 = (inp[4]) ? 3'b110 : node545;
											assign node545 = (inp[1]) ? 3'b110 : 3'b111;
						assign node550 = (inp[3]) ? node590 : node551;
							assign node551 = (inp[4]) ? node575 : node552;
								assign node552 = (inp[7]) ? node566 : node553;
									assign node553 = (inp[1]) ? node559 : node554;
										assign node554 = (inp[9]) ? node556 : 3'b111;
											assign node556 = (inp[2]) ? 3'b111 : 3'b110;
										assign node559 = (inp[2]) ? node563 : node560;
											assign node560 = (inp[9]) ? 3'b110 : 3'b110;
											assign node563 = (inp[9]) ? 3'b110 : 3'b110;
									assign node566 = (inp[9]) ? 3'b111 : node567;
										assign node567 = (inp[0]) ? node571 : node568;
											assign node568 = (inp[2]) ? 3'b111 : 3'b110;
											assign node571 = (inp[1]) ? 3'b111 : 3'b110;
								assign node575 = (inp[0]) ? node583 : node576;
									assign node576 = (inp[2]) ? node578 : 3'b101;
										assign node578 = (inp[1]) ? 3'b101 : node579;
											assign node579 = (inp[7]) ? 3'b100 : 3'b101;
									assign node583 = (inp[1]) ? 3'b100 : node584;
										assign node584 = (inp[2]) ? 3'b100 : node585;
											assign node585 = (inp[7]) ? 3'b100 : 3'b101;
							assign node590 = (inp[4]) ? node610 : node591;
								assign node591 = (inp[0]) ? node601 : node592;
									assign node592 = (inp[2]) ? 3'b100 : node593;
										assign node593 = (inp[9]) ? node597 : node594;
											assign node594 = (inp[1]) ? 3'b101 : 3'b100;
											assign node597 = (inp[1]) ? 3'b100 : 3'b101;
									assign node601 = (inp[9]) ? node605 : node602;
										assign node602 = (inp[1]) ? 3'b100 : 3'b101;
										assign node605 = (inp[1]) ? node607 : 3'b100;
											assign node607 = (inp[7]) ? 3'b100 : 3'b101;
								assign node610 = (inp[1]) ? node624 : node611;
									assign node611 = (inp[7]) ? node619 : node612;
										assign node612 = (inp[2]) ? node616 : node613;
											assign node613 = (inp[0]) ? 3'b101 : 3'b100;
											assign node616 = (inp[0]) ? 3'b100 : 3'b101;
										assign node619 = (inp[0]) ? 3'b100 : node620;
											assign node620 = (inp[2]) ? 3'b101 : 3'b100;
									assign node624 = (inp[0]) ? node628 : node625;
										assign node625 = (inp[2]) ? 3'b101 : 3'b100;
										assign node628 = (inp[2]) ? 3'b100 : 3'b101;
			assign node631 = (inp[4]) ? node887 : node632;
				assign node632 = (inp[6]) ? node780 : node633;
					assign node633 = (inp[11]) ? node707 : node634;
						assign node634 = (inp[7]) ? node668 : node635;
							assign node635 = (inp[3]) ? node655 : node636;
								assign node636 = (inp[0]) ? node650 : node637;
									assign node637 = (inp[10]) ? node643 : node638;
										assign node638 = (inp[9]) ? 3'b101 : node639;
											assign node639 = (inp[1]) ? 3'b101 : 3'b100;
										assign node643 = (inp[9]) ? node647 : node644;
											assign node644 = (inp[1]) ? 3'b101 : 3'b100;
											assign node647 = (inp[1]) ? 3'b100 : 3'b101;
									assign node650 = (inp[9]) ? node652 : 3'b101;
										assign node652 = (inp[1]) ? 3'b100 : 3'b101;
								assign node655 = (inp[9]) ? node661 : node656;
									assign node656 = (inp[2]) ? 3'b111 : node657;
										assign node657 = (inp[1]) ? 3'b111 : 3'b110;
									assign node661 = (inp[0]) ? 3'b110 : node662;
										assign node662 = (inp[2]) ? node664 : 3'b111;
											assign node664 = (inp[10]) ? 3'b110 : 3'b110;
							assign node668 = (inp[3]) ? node684 : node669;
								assign node669 = (inp[1]) ? node679 : node670;
									assign node670 = (inp[9]) ? node674 : node671;
										assign node671 = (inp[10]) ? 3'b111 : 3'b110;
										assign node674 = (inp[10]) ? node676 : 3'b111;
											assign node676 = (inp[2]) ? 3'b110 : 3'b111;
									assign node679 = (inp[10]) ? 3'b110 : node680;
										assign node680 = (inp[9]) ? 3'b110 : 3'b111;
								assign node684 = (inp[10]) ? node696 : node685;
									assign node685 = (inp[9]) ? node691 : node686;
										assign node686 = (inp[2]) ? node688 : 3'b100;
											assign node688 = (inp[1]) ? 3'b101 : 3'b100;
										assign node691 = (inp[2]) ? node693 : 3'b101;
											assign node693 = (inp[1]) ? 3'b100 : 3'b101;
									assign node696 = (inp[2]) ? node702 : node697;
										assign node697 = (inp[9]) ? node699 : 3'b100;
											assign node699 = (inp[1]) ? 3'b100 : 3'b101;
										assign node702 = (inp[0]) ? 3'b100 : node703;
											assign node703 = (inp[9]) ? 3'b100 : 3'b100;
						assign node707 = (inp[7]) ? node749 : node708;
							assign node708 = (inp[3]) ? node730 : node709;
								assign node709 = (inp[9]) ? node719 : node710;
									assign node710 = (inp[1]) ? node714 : node711;
										assign node711 = (inp[10]) ? 3'b101 : 3'b100;
										assign node714 = (inp[10]) ? node716 : 3'b101;
											assign node716 = (inp[2]) ? 3'b101 : 3'b100;
									assign node719 = (inp[1]) ? node725 : node720;
										assign node720 = (inp[2]) ? 3'b101 : node721;
											assign node721 = (inp[10]) ? 3'b100 : 3'b101;
										assign node725 = (inp[2]) ? 3'b100 : node726;
											assign node726 = (inp[10]) ? 3'b101 : 3'b100;
								assign node730 = (inp[0]) ? node740 : node731;
									assign node731 = (inp[2]) ? node733 : 3'b110;
										assign node733 = (inp[10]) ? node737 : node734;
											assign node734 = (inp[1]) ? 3'b111 : 3'b110;
											assign node737 = (inp[9]) ? 3'b110 : 3'b110;
									assign node740 = (inp[1]) ? node744 : node741;
										assign node741 = (inp[9]) ? 3'b111 : 3'b110;
										assign node744 = (inp[9]) ? 3'b110 : node745;
											assign node745 = (inp[10]) ? 3'b110 : 3'b111;
							assign node749 = (inp[3]) ? node759 : node750;
								assign node750 = (inp[2]) ? node752 : 3'b111;
									assign node752 = (inp[9]) ? 3'b110 : node753;
										assign node753 = (inp[10]) ? node755 : 3'b111;
											assign node755 = (inp[1]) ? 3'b111 : 3'b110;
								assign node759 = (inp[1]) ? node771 : node760;
									assign node760 = (inp[9]) ? node766 : node761;
										assign node761 = (inp[10]) ? node763 : 3'b100;
											assign node763 = (inp[2]) ? 3'b100 : 3'b101;
										assign node766 = (inp[10]) ? node768 : 3'b101;
											assign node768 = (inp[2]) ? 3'b101 : 3'b100;
									assign node771 = (inp[9]) ? node777 : node772;
										assign node772 = (inp[10]) ? node774 : 3'b101;
											assign node774 = (inp[2]) ? 3'b101 : 3'b100;
										assign node777 = (inp[2]) ? 3'b100 : 3'b101;
					assign node780 = (inp[9]) ? node834 : node781;
						assign node781 = (inp[10]) ? node811 : node782;
							assign node782 = (inp[7]) ? node798 : node783;
								assign node783 = (inp[2]) ? node791 : node784;
									assign node784 = (inp[11]) ? node788 : node785;
										assign node785 = (inp[3]) ? 3'b010 : 3'b000;
										assign node788 = (inp[3]) ? 3'b000 : 3'b010;
									assign node791 = (inp[11]) ? node795 : node792;
										assign node792 = (inp[3]) ? 3'b010 : 3'b000;
										assign node795 = (inp[3]) ? 3'b001 : 3'b010;
								assign node798 = (inp[3]) ? node804 : node799;
									assign node799 = (inp[11]) ? 3'b011 : node800;
										assign node800 = (inp[2]) ? 3'b001 : 3'b000;
									assign node804 = (inp[11]) ? node808 : node805;
										assign node805 = (inp[2]) ? 3'b010 : 3'b011;
										assign node808 = (inp[2]) ? 3'b001 : 3'b000;
							assign node811 = (inp[2]) ? node823 : node812;
								assign node812 = (inp[3]) ? node818 : node813;
									assign node813 = (inp[11]) ? node815 : 3'b001;
										assign node815 = (inp[7]) ? 3'b011 : 3'b010;
									assign node818 = (inp[11]) ? 3'b000 : node819;
										assign node819 = (inp[7]) ? 3'b010 : 3'b011;
								assign node823 = (inp[3]) ? node831 : node824;
									assign node824 = (inp[11]) ? node828 : node825;
										assign node825 = (inp[7]) ? 3'b000 : 3'b001;
										assign node828 = (inp[7]) ? 3'b011 : 3'b010;
									assign node831 = (inp[11]) ? 3'b001 : 3'b011;
						assign node834 = (inp[2]) ? node866 : node835;
							assign node835 = (inp[10]) ? node859 : node836;
								assign node836 = (inp[7]) ? node848 : node837;
									assign node837 = (inp[1]) ? node843 : node838;
										assign node838 = (inp[11]) ? 3'b001 : node839;
											assign node839 = (inp[3]) ? 3'b011 : 3'b001;
										assign node843 = (inp[0]) ? 3'b011 : node844;
											assign node844 = (inp[11]) ? 3'b011 : 3'b001;
									assign node848 = (inp[1]) ? node854 : node849;
										assign node849 = (inp[3]) ? node851 : 3'b001;
											assign node851 = (inp[0]) ? 3'b001 : 3'b010;
										assign node854 = (inp[3]) ? node856 : 3'b010;
											assign node856 = (inp[11]) ? 3'b001 : 3'b010;
								assign node859 = (inp[3]) ? node861 : 3'b000;
									assign node861 = (inp[11]) ? 3'b001 : node862;
										assign node862 = (inp[7]) ? 3'b011 : 3'b010;
							assign node866 = (inp[3]) ? node882 : node867;
								assign node867 = (inp[11]) ? node879 : node868;
									assign node868 = (inp[0]) ? node874 : node869;
										assign node869 = (inp[7]) ? 3'b001 : node870;
											assign node870 = (inp[10]) ? 3'b000 : 3'b001;
										assign node874 = (inp[10]) ? node876 : 3'b000;
											assign node876 = (inp[7]) ? 3'b001 : 3'b000;
									assign node879 = (inp[7]) ? 3'b010 : 3'b011;
								assign node882 = (inp[11]) ? 3'b000 : node883;
									assign node883 = (inp[10]) ? 3'b010 : 3'b011;
				assign node887 = (inp[11]) ? node959 : node888;
					assign node888 = (inp[6]) ? node952 : node889;
						assign node889 = (inp[7]) ? node919 : node890;
							assign node890 = (inp[10]) ? node898 : node891;
								assign node891 = (inp[1]) ? node895 : node892;
									assign node892 = (inp[2]) ? 3'b001 : 3'b000;
									assign node895 = (inp[2]) ? 3'b000 : 3'b001;
								assign node898 = (inp[9]) ? node908 : node899;
									assign node899 = (inp[3]) ? node901 : 3'b000;
										assign node901 = (inp[1]) ? node905 : node902;
											assign node902 = (inp[2]) ? 3'b000 : 3'b001;
											assign node905 = (inp[2]) ? 3'b001 : 3'b000;
									assign node908 = (inp[0]) ? node914 : node909;
										assign node909 = (inp[2]) ? node911 : 3'b001;
											assign node911 = (inp[3]) ? 3'b001 : 3'b000;
										assign node914 = (inp[3]) ? 3'b000 : node915;
											assign node915 = (inp[1]) ? 3'b000 : 3'b001;
							assign node919 = (inp[10]) ? node937 : node920;
								assign node920 = (inp[0]) ? node928 : node921;
									assign node921 = (inp[2]) ? 3'b011 : node922;
										assign node922 = (inp[3]) ? node924 : 3'b010;
											assign node924 = (inp[1]) ? 3'b010 : 3'b011;
									assign node928 = (inp[2]) ? node930 : 3'b011;
										assign node930 = (inp[9]) ? node934 : node931;
											assign node931 = (inp[1]) ? 3'b010 : 3'b011;
											assign node934 = (inp[1]) ? 3'b011 : 3'b010;
								assign node937 = (inp[9]) ? node945 : node938;
									assign node938 = (inp[1]) ? node942 : node939;
										assign node939 = (inp[2]) ? 3'b011 : 3'b010;
										assign node942 = (inp[2]) ? 3'b010 : 3'b011;
									assign node945 = (inp[2]) ? node949 : node946;
										assign node946 = (inp[1]) ? 3'b011 : 3'b010;
										assign node949 = (inp[1]) ? 3'b010 : 3'b011;
						assign node952 = (inp[10]) ? node956 : node953;
							assign node953 = (inp[2]) ? 3'b011 : 3'b010;
							assign node956 = (inp[2]) ? 3'b010 : 3'b011;
					assign node959 = (inp[6]) ? node1017 : node960;
						assign node960 = (inp[7]) ? node1002 : node961;
							assign node961 = (inp[9]) ? node983 : node962;
								assign node962 = (inp[0]) ? node976 : node963;
									assign node963 = (inp[10]) ? node971 : node964;
										assign node964 = (inp[1]) ? node968 : node965;
											assign node965 = (inp[2]) ? 3'b011 : 3'b010;
											assign node968 = (inp[2]) ? 3'b010 : 3'b011;
										assign node971 = (inp[2]) ? 3'b010 : node972;
											assign node972 = (inp[3]) ? 3'b010 : 3'b010;
									assign node976 = (inp[2]) ? node978 : 3'b010;
										assign node978 = (inp[3]) ? 3'b010 : node979;
											assign node979 = (inp[10]) ? 3'b011 : 3'b010;
								assign node983 = (inp[1]) ? node995 : node984;
									assign node984 = (inp[2]) ? node990 : node985;
										assign node985 = (inp[10]) ? node987 : 3'b010;
											assign node987 = (inp[3]) ? 3'b010 : 3'b011;
										assign node990 = (inp[3]) ? 3'b011 : node991;
											assign node991 = (inp[10]) ? 3'b010 : 3'b011;
									assign node995 = (inp[2]) ? 3'b010 : node996;
										assign node996 = (inp[3]) ? 3'b011 : node997;
											assign node997 = (inp[10]) ? 3'b010 : 3'b011;
							assign node1002 = (inp[2]) ? node1012 : node1003;
								assign node1003 = (inp[10]) ? node1009 : node1004;
									assign node1004 = (inp[3]) ? 3'b000 : node1005;
										assign node1005 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1009 = (inp[1]) ? 3'b001 : 3'b000;
								assign node1012 = (inp[1]) ? node1014 : 3'b001;
									assign node1014 = (inp[3]) ? 3'b000 : 3'b001;
						assign node1017 = (inp[2]) ? node1023 : node1018;
							assign node1018 = (inp[7]) ? 3'b001 : node1019;
								assign node1019 = (inp[3]) ? 3'b001 : 3'b000;
							assign node1023 = (inp[7]) ? 3'b000 : node1024;
								assign node1024 = (inp[3]) ? 3'b000 : 3'b001;
		assign node1028 = (inp[4]) ? node1536 : node1029;
			assign node1029 = (inp[6]) ? node1319 : node1030;
				assign node1030 = (inp[3]) ? node1184 : node1031;
					assign node1031 = (inp[7]) ? node1115 : node1032;
						assign node1032 = (inp[8]) ? node1078 : node1033;
							assign node1033 = (inp[11]) ? node1057 : node1034;
								assign node1034 = (inp[10]) ? node1044 : node1035;
									assign node1035 = (inp[1]) ? node1041 : node1036;
										assign node1036 = (inp[2]) ? 3'b101 : node1037;
											assign node1037 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1041 = (inp[2]) ? 3'b100 : 3'b101;
									assign node1044 = (inp[9]) ? node1050 : node1045;
										assign node1045 = (inp[1]) ? 3'b111 : node1046;
											assign node1046 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1050 = (inp[0]) ? node1054 : node1051;
											assign node1051 = (inp[2]) ? 3'b110 : 3'b111;
											assign node1054 = (inp[2]) ? 3'b111 : 3'b110;
								assign node1057 = (inp[10]) ? node1069 : node1058;
									assign node1058 = (inp[9]) ? node1064 : node1059;
										assign node1059 = (inp[0]) ? node1061 : 3'b110;
											assign node1061 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1064 = (inp[1]) ? 3'b111 : node1065;
											assign node1065 = (inp[2]) ? 3'b110 : 3'b110;
									assign node1069 = (inp[1]) ? node1073 : node1070;
										assign node1070 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1073 = (inp[2]) ? 3'b100 : node1074;
											assign node1074 = (inp[9]) ? 3'b100 : 3'b101;
							assign node1078 = (inp[11]) ? node1100 : node1079;
								assign node1079 = (inp[10]) ? node1093 : node1080;
									assign node1080 = (inp[2]) ? node1088 : node1081;
										assign node1081 = (inp[0]) ? node1085 : node1082;
											assign node1082 = (inp[1]) ? 3'b101 : 3'b100;
											assign node1085 = (inp[9]) ? 3'b100 : 3'b100;
										assign node1088 = (inp[0]) ? 3'b101 : node1089;
											assign node1089 = (inp[1]) ? 3'b100 : 3'b100;
									assign node1093 = (inp[2]) ? 3'b101 : node1094;
										assign node1094 = (inp[1]) ? 3'b101 : node1095;
											assign node1095 = (inp[0]) ? 3'b100 : 3'b101;
								assign node1100 = (inp[2]) ? node1108 : node1101;
									assign node1101 = (inp[1]) ? node1105 : node1102;
										assign node1102 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1105 = (inp[9]) ? 3'b100 : 3'b101;
									assign node1108 = (inp[0]) ? node1110 : 3'b100;
										assign node1110 = (inp[10]) ? 3'b100 : node1111;
											assign node1111 = (inp[1]) ? 3'b101 : 3'b100;
						assign node1115 = (inp[10]) ? node1153 : node1116;
							assign node1116 = (inp[8]) ? node1138 : node1117;
								assign node1117 = (inp[2]) ? node1131 : node1118;
									assign node1118 = (inp[0]) ? node1124 : node1119;
										assign node1119 = (inp[11]) ? node1121 : 3'b101;
											assign node1121 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1124 = (inp[1]) ? node1128 : node1125;
											assign node1125 = (inp[9]) ? 3'b100 : 3'b100;
											assign node1128 = (inp[9]) ? 3'b100 : 3'b100;
									assign node1131 = (inp[11]) ? 3'b101 : node1132;
										assign node1132 = (inp[9]) ? node1134 : 3'b101;
											assign node1134 = (inp[1]) ? 3'b101 : 3'b100;
								assign node1138 = (inp[11]) ? 3'b111 : node1139;
									assign node1139 = (inp[2]) ? node1145 : node1140;
										assign node1140 = (inp[9]) ? 3'b110 : node1141;
											assign node1141 = (inp[1]) ? 3'b111 : 3'b110;
										assign node1145 = (inp[1]) ? node1149 : node1146;
											assign node1146 = (inp[9]) ? 3'b110 : 3'b111;
											assign node1149 = (inp[9]) ? 3'b111 : 3'b110;
							assign node1153 = (inp[11]) ? node1167 : node1154;
								assign node1154 = (inp[9]) ? node1162 : node1155;
									assign node1155 = (inp[1]) ? 3'b111 : node1156;
										assign node1156 = (inp[8]) ? 3'b110 : node1157;
											assign node1157 = (inp[2]) ? 3'b111 : 3'b110;
									assign node1162 = (inp[1]) ? node1164 : 3'b111;
										assign node1164 = (inp[0]) ? 3'b110 : 3'b111;
								assign node1167 = (inp[8]) ? node1177 : node1168;
									assign node1168 = (inp[2]) ? 3'b110 : node1169;
										assign node1169 = (inp[0]) ? node1173 : node1170;
											assign node1170 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1173 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1177 = (inp[9]) ? node1181 : node1178;
										assign node1178 = (inp[1]) ? 3'b111 : 3'b110;
										assign node1181 = (inp[1]) ? 3'b110 : 3'b111;
					assign node1184 = (inp[7]) ? node1262 : node1185;
						assign node1185 = (inp[8]) ? node1237 : node1186;
							assign node1186 = (inp[1]) ? node1216 : node1187;
								assign node1187 = (inp[2]) ? node1201 : node1188;
									assign node1188 = (inp[9]) ? node1194 : node1189;
										assign node1189 = (inp[0]) ? 3'b111 : node1190;
											assign node1190 = (inp[10]) ? 3'b101 : 3'b100;
										assign node1194 = (inp[10]) ? node1198 : node1195;
											assign node1195 = (inp[0]) ? 3'b101 : 3'b111;
											assign node1198 = (inp[11]) ? 3'b110 : 3'b100;
									assign node1201 = (inp[0]) ? node1209 : node1202;
										assign node1202 = (inp[9]) ? node1206 : node1203;
											assign node1203 = (inp[11]) ? 3'b100 : 3'b100;
											assign node1206 = (inp[11]) ? 3'b101 : 3'b111;
										assign node1209 = (inp[9]) ? node1213 : node1210;
											assign node1210 = (inp[10]) ? 3'b100 : 3'b101;
											assign node1213 = (inp[10]) ? 3'b100 : 3'b100;
								assign node1216 = (inp[11]) ? node1226 : node1217;
									assign node1217 = (inp[10]) ? node1223 : node1218;
										assign node1218 = (inp[9]) ? 3'b110 : node1219;
											assign node1219 = (inp[0]) ? 3'b110 : 3'b110;
										assign node1223 = (inp[2]) ? 3'b101 : 3'b100;
									assign node1226 = (inp[10]) ? node1232 : node1227;
										assign node1227 = (inp[9]) ? 3'b100 : node1228;
											assign node1228 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1232 = (inp[0]) ? 3'b110 : node1233;
											assign node1233 = (inp[9]) ? 3'b111 : 3'b110;
							assign node1237 = (inp[10]) ? node1249 : node1238;
								assign node1238 = (inp[1]) ? 3'b110 : node1239;
									assign node1239 = (inp[9]) ? node1245 : node1240;
										assign node1240 = (inp[11]) ? node1242 : 3'b110;
											assign node1242 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1245 = (inp[11]) ? 3'b110 : 3'b111;
								assign node1249 = (inp[1]) ? node1257 : node1250;
									assign node1250 = (inp[9]) ? node1254 : node1251;
										assign node1251 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1254 = (inp[2]) ? 3'b111 : 3'b110;
									assign node1257 = (inp[9]) ? node1259 : 3'b111;
										assign node1259 = (inp[2]) ? 3'b110 : 3'b111;
						assign node1262 = (inp[8]) ? node1284 : node1263;
							assign node1263 = (inp[10]) ? node1277 : node1264;
								assign node1264 = (inp[2]) ? node1270 : node1265;
									assign node1265 = (inp[0]) ? 3'b110 : node1266;
										assign node1266 = (inp[11]) ? 3'b111 : 3'b110;
									assign node1270 = (inp[9]) ? 3'b111 : node1271;
										assign node1271 = (inp[1]) ? 3'b111 : node1272;
											assign node1272 = (inp[0]) ? 3'b111 : 3'b110;
								assign node1277 = (inp[0]) ? node1281 : node1278;
									assign node1278 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1281 = (inp[9]) ? 3'b100 : 3'b101;
							assign node1284 = (inp[11]) ? node1304 : node1285;
								assign node1285 = (inp[10]) ? node1299 : node1286;
									assign node1286 = (inp[9]) ? node1294 : node1287;
										assign node1287 = (inp[0]) ? node1291 : node1288;
											assign node1288 = (inp[1]) ? 3'b100 : 3'b101;
											assign node1291 = (inp[1]) ? 3'b101 : 3'b100;
										assign node1294 = (inp[2]) ? 3'b100 : node1295;
											assign node1295 = (inp[1]) ? 3'b100 : 3'b101;
									assign node1299 = (inp[1]) ? 3'b100 : node1300;
										assign node1300 = (inp[9]) ? 3'b101 : 3'b100;
								assign node1304 = (inp[0]) ? node1310 : node1305;
									assign node1305 = (inp[2]) ? 3'b101 : node1306;
										assign node1306 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1310 = (inp[1]) ? node1316 : node1311;
										assign node1311 = (inp[10]) ? 3'b100 : node1312;
											assign node1312 = (inp[9]) ? 3'b100 : 3'b100;
										assign node1316 = (inp[9]) ? 3'b100 : 3'b101;
				assign node1319 = (inp[3]) ? node1433 : node1320;
					assign node1320 = (inp[8]) ? node1398 : node1321;
						assign node1321 = (inp[10]) ? node1353 : node1322;
							assign node1322 = (inp[11]) ? node1338 : node1323;
								assign node1323 = (inp[7]) ? node1333 : node1324;
									assign node1324 = (inp[0]) ? node1330 : node1325;
										assign node1325 = (inp[9]) ? node1327 : 3'b011;
											assign node1327 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1330 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1333 = (inp[9]) ? node1335 : 3'b000;
										assign node1335 = (inp[0]) ? 3'b000 : 3'b001;
								assign node1338 = (inp[0]) ? 3'b001 : node1339;
									assign node1339 = (inp[2]) ? node1347 : node1340;
										assign node1340 = (inp[1]) ? node1344 : node1341;
											assign node1341 = (inp[7]) ? 3'b000 : 3'b000;
											assign node1344 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1347 = (inp[1]) ? node1349 : 3'b001;
											assign node1349 = (inp[9]) ? 3'b000 : 3'b001;
							assign node1353 = (inp[11]) ? node1379 : node1354;
								assign node1354 = (inp[7]) ? node1368 : node1355;
									assign node1355 = (inp[9]) ? node1361 : node1356;
										assign node1356 = (inp[0]) ? 3'b001 : node1357;
											assign node1357 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1361 = (inp[0]) ? node1365 : node1362;
											assign node1362 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1365 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1368 = (inp[2]) ? node1374 : node1369;
										assign node1369 = (inp[1]) ? node1371 : 3'b010;
											assign node1371 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1374 = (inp[0]) ? node1376 : 3'b011;
											assign node1376 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1379 = (inp[2]) ? node1385 : node1380;
									assign node1380 = (inp[0]) ? node1382 : 3'b010;
										assign node1382 = (inp[7]) ? 3'b011 : 3'b010;
									assign node1385 = (inp[9]) ? node1393 : node1386;
										assign node1386 = (inp[7]) ? node1390 : node1387;
											assign node1387 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1390 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1393 = (inp[1]) ? 3'b011 : node1394;
											assign node1394 = (inp[7]) ? 3'b011 : 3'b010;
						assign node1398 = (inp[9]) ? node1420 : node1399;
							assign node1399 = (inp[7]) ? node1415 : node1400;
								assign node1400 = (inp[11]) ? 3'b010 : node1401;
									assign node1401 = (inp[1]) ? node1409 : node1402;
										assign node1402 = (inp[2]) ? node1406 : node1403;
											assign node1403 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1406 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1409 = (inp[2]) ? node1411 : 3'b011;
											assign node1411 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1415 = (inp[10]) ? 3'b011 : node1416;
									assign node1416 = (inp[11]) ? 3'b011 : 3'b010;
							assign node1420 = (inp[7]) ? node1428 : node1421;
								assign node1421 = (inp[11]) ? 3'b011 : node1422;
									assign node1422 = (inp[10]) ? node1424 : 3'b010;
										assign node1424 = (inp[2]) ? 3'b011 : 3'b010;
								assign node1428 = (inp[10]) ? 3'b010 : node1429;
									assign node1429 = (inp[2]) ? 3'b010 : 3'b011;
					assign node1433 = (inp[8]) ? node1511 : node1434;
						assign node1434 = (inp[10]) ? node1474 : node1435;
							assign node1435 = (inp[7]) ? node1453 : node1436;
								assign node1436 = (inp[11]) ? node1444 : node1437;
									assign node1437 = (inp[0]) ? 3'b001 : node1438;
										assign node1438 = (inp[1]) ? 3'b000 : node1439;
											assign node1439 = (inp[9]) ? 3'b000 : 3'b000;
									assign node1444 = (inp[9]) ? node1448 : node1445;
										assign node1445 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1448 = (inp[2]) ? 3'b011 : node1449;
											assign node1449 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1453 = (inp[1]) ? node1461 : node1454;
									assign node1454 = (inp[11]) ? node1456 : 3'b011;
										assign node1456 = (inp[9]) ? node1458 : 3'b011;
											assign node1458 = (inp[2]) ? 3'b011 : 3'b010;
									assign node1461 = (inp[9]) ? node1469 : node1462;
										assign node1462 = (inp[0]) ? node1466 : node1463;
											assign node1463 = (inp[11]) ? 3'b010 : 3'b011;
											assign node1466 = (inp[11]) ? 3'b011 : 3'b010;
										assign node1469 = (inp[2]) ? 3'b010 : node1470;
											assign node1470 = (inp[11]) ? 3'b010 : 3'b011;
							assign node1474 = (inp[11]) ? node1494 : node1475;
								assign node1475 = (inp[7]) ? node1489 : node1476;
									assign node1476 = (inp[0]) ? node1484 : node1477;
										assign node1477 = (inp[9]) ? node1481 : node1478;
											assign node1478 = (inp[1]) ? 3'b010 : 3'b011;
											assign node1481 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1484 = (inp[9]) ? 3'b011 : node1485;
											assign node1485 = (inp[1]) ? 3'b011 : 3'b010;
									assign node1489 = (inp[0]) ? 3'b001 : node1490;
										assign node1490 = (inp[1]) ? 3'b001 : 3'b000;
								assign node1494 = (inp[1]) ? node1502 : node1495;
									assign node1495 = (inp[2]) ? 3'b001 : node1496;
										assign node1496 = (inp[7]) ? node1498 : 3'b000;
											assign node1498 = (inp[0]) ? 3'b000 : 3'b001;
									assign node1502 = (inp[2]) ? node1506 : node1503;
										assign node1503 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1506 = (inp[0]) ? 3'b000 : node1507;
											assign node1507 = (inp[9]) ? 3'b001 : 3'b000;
						assign node1511 = (inp[9]) ? node1525 : node1512;
							assign node1512 = (inp[11]) ? 3'b001 : node1513;
								assign node1513 = (inp[10]) ? node1519 : node1514;
									assign node1514 = (inp[7]) ? 3'b000 : node1515;
										assign node1515 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1519 = (inp[7]) ? 3'b001 : node1520;
										assign node1520 = (inp[2]) ? 3'b001 : 3'b000;
							assign node1525 = (inp[11]) ? 3'b000 : node1526;
								assign node1526 = (inp[10]) ? node1528 : 3'b001;
									assign node1528 = (inp[0]) ? node1530 : 3'b001;
										assign node1530 = (inp[1]) ? 3'b000 : node1531;
											assign node1531 = (inp[7]) ? 3'b000 : 3'b001;
			assign node1536 = (inp[10]) ? node1710 : node1537;
				assign node1537 = (inp[8]) ? node1663 : node1538;
					assign node1538 = (inp[7]) ? node1612 : node1539;
						assign node1539 = (inp[6]) ? node1581 : node1540;
							assign node1540 = (inp[2]) ? node1564 : node1541;
								assign node1541 = (inp[1]) ? node1553 : node1542;
									assign node1542 = (inp[9]) ? node1548 : node1543;
										assign node1543 = (inp[0]) ? 3'b000 : node1544;
											assign node1544 = (inp[11]) ? 3'b001 : 3'b000;
										assign node1548 = (inp[3]) ? node1550 : 3'b001;
											assign node1550 = (inp[0]) ? 3'b000 : 3'b001;
									assign node1553 = (inp[9]) ? node1559 : node1554;
										assign node1554 = (inp[0]) ? 3'b001 : node1555;
											assign node1555 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1559 = (inp[3]) ? 3'b000 : node1560;
											assign node1560 = (inp[0]) ? 3'b000 : 3'b000;
								assign node1564 = (inp[9]) ? node1576 : node1565;
									assign node1565 = (inp[3]) ? node1571 : node1566;
										assign node1566 = (inp[0]) ? 3'b001 : node1567;
											assign node1567 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1571 = (inp[0]) ? 3'b000 : node1572;
											assign node1572 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1576 = (inp[11]) ? node1578 : 3'b001;
										assign node1578 = (inp[1]) ? 3'b001 : 3'b000;
							assign node1581 = (inp[9]) ? node1599 : node1582;
								assign node1582 = (inp[1]) ? node1588 : node1583;
									assign node1583 = (inp[0]) ? node1585 : 3'b011;
										assign node1585 = (inp[3]) ? 3'b010 : 3'b011;
									assign node1588 = (inp[11]) ? node1594 : node1589;
										assign node1589 = (inp[2]) ? 3'b010 : node1590;
											assign node1590 = (inp[0]) ? 3'b010 : 3'b011;
										assign node1594 = (inp[2]) ? node1596 : 3'b010;
											assign node1596 = (inp[3]) ? 3'b011 : 3'b010;
								assign node1599 = (inp[3]) ? node1605 : node1600;
									assign node1600 = (inp[0]) ? node1602 : 3'b010;
										assign node1602 = (inp[11]) ? 3'b011 : 3'b010;
									assign node1605 = (inp[0]) ? 3'b010 : node1606;
										assign node1606 = (inp[1]) ? node1608 : 3'b011;
											assign node1608 = (inp[11]) ? 3'b011 : 3'b010;
						assign node1612 = (inp[3]) ? node1656 : node1613;
							assign node1613 = (inp[6]) ? node1637 : node1614;
								assign node1614 = (inp[1]) ? node1624 : node1615;
									assign node1615 = (inp[2]) ? node1621 : node1616;
										assign node1616 = (inp[0]) ? 3'b011 : node1617;
											assign node1617 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1621 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1624 = (inp[9]) ? node1630 : node1625;
										assign node1625 = (inp[0]) ? 3'b010 : node1626;
											assign node1626 = (inp[11]) ? 3'b011 : 3'b010;
										assign node1630 = (inp[0]) ? node1634 : node1631;
											assign node1631 = (inp[11]) ? 3'b011 : 3'b010;
											assign node1634 = (inp[11]) ? 3'b010 : 3'b011;
								assign node1637 = (inp[2]) ? node1651 : node1638;
									assign node1638 = (inp[9]) ? node1646 : node1639;
										assign node1639 = (inp[1]) ? node1643 : node1640;
											assign node1640 = (inp[0]) ? 3'b010 : 3'b010;
											assign node1643 = (inp[11]) ? 3'b011 : 3'b010;
										assign node1646 = (inp[0]) ? node1648 : 3'b011;
											assign node1648 = (inp[11]) ? 3'b010 : 3'b011;
									assign node1651 = (inp[11]) ? node1653 : 3'b011;
										assign node1653 = (inp[0]) ? 3'b010 : 3'b011;
							assign node1656 = (inp[11]) ? node1660 : node1657;
								assign node1657 = (inp[0]) ? 3'b011 : 3'b010;
								assign node1660 = (inp[0]) ? 3'b010 : 3'b011;
					assign node1663 = (inp[6]) ? node1699 : node1664;
						assign node1664 = (inp[7]) ? node1672 : node1665;
							assign node1665 = (inp[1]) ? node1669 : node1666;
								assign node1666 = (inp[3]) ? 3'b011 : 3'b010;
								assign node1669 = (inp[3]) ? 3'b010 : 3'b011;
							assign node1672 = (inp[3]) ? node1690 : node1673;
								assign node1673 = (inp[9]) ? node1681 : node1674;
									assign node1674 = (inp[11]) ? node1678 : node1675;
										assign node1675 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1678 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1681 = (inp[0]) ? node1683 : 3'b001;
										assign node1683 = (inp[1]) ? node1687 : node1684;
											assign node1684 = (inp[11]) ? 3'b001 : 3'b000;
											assign node1687 = (inp[11]) ? 3'b000 : 3'b001;
								assign node1690 = (inp[2]) ? 3'b000 : node1691;
									assign node1691 = (inp[1]) ? node1695 : node1692;
										assign node1692 = (inp[11]) ? 3'b001 : 3'b000;
										assign node1695 = (inp[11]) ? 3'b000 : 3'b001;
						assign node1699 = (inp[11]) ? node1705 : node1700;
							assign node1700 = (inp[7]) ? 3'b001 : node1701;
								assign node1701 = (inp[3]) ? 3'b001 : 3'b000;
							assign node1705 = (inp[3]) ? 3'b000 : node1706;
								assign node1706 = (inp[7]) ? 3'b000 : 3'b001;
				assign node1710 = (inp[7]) ? node1780 : node1711;
					assign node1711 = (inp[6]) ? node1753 : node1712;
						assign node1712 = (inp[8]) ? node1746 : node1713;
							assign node1713 = (inp[11]) ? node1721 : node1714;
								assign node1714 = (inp[3]) ? node1718 : node1715;
									assign node1715 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1718 = (inp[0]) ? 3'b010 : 3'b011;
								assign node1721 = (inp[0]) ? node1731 : node1722;
									assign node1722 = (inp[2]) ? node1728 : node1723;
										assign node1723 = (inp[9]) ? 3'b011 : node1724;
											assign node1724 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1728 = (inp[9]) ? 3'b010 : 3'b011;
									assign node1731 = (inp[2]) ? node1739 : node1732;
										assign node1732 = (inp[3]) ? node1736 : node1733;
											assign node1733 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1736 = (inp[1]) ? 3'b010 : 3'b011;
										assign node1739 = (inp[3]) ? node1743 : node1740;
											assign node1740 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1743 = (inp[1]) ? 3'b010 : 3'b011;
							assign node1746 = (inp[3]) ? node1750 : node1747;
								assign node1747 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1750 = (inp[1]) ? 3'b010 : 3'b011;
						assign node1753 = (inp[3]) ? node1767 : node1754;
							assign node1754 = (inp[8]) ? 3'b001 : node1755;
								assign node1755 = (inp[0]) ? node1761 : node1756;
									assign node1756 = (inp[11]) ? 3'b000 : node1757;
										assign node1757 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1761 = (inp[11]) ? 3'b001 : node1762;
										assign node1762 = (inp[1]) ? 3'b001 : 3'b000;
							assign node1767 = (inp[8]) ? 3'b000 : node1768;
								assign node1768 = (inp[0]) ? node1774 : node1769;
									assign node1769 = (inp[1]) ? 3'b001 : node1770;
										assign node1770 = (inp[11]) ? 3'b001 : 3'b000;
									assign node1774 = (inp[11]) ? 3'b000 : node1775;
										assign node1775 = (inp[1]) ? 3'b000 : 3'b001;
					assign node1780 = (inp[1]) ? node1792 : node1781;
						assign node1781 = (inp[6]) ? node1787 : node1782;
							assign node1782 = (inp[0]) ? 3'b001 : node1783;
								assign node1783 = (inp[8]) ? 3'b001 : 3'b000;
							assign node1787 = (inp[0]) ? 3'b000 : node1788;
								assign node1788 = (inp[8]) ? 3'b000 : 3'b001;
						assign node1792 = (inp[8]) ? 3'b000 : node1793;
							assign node1793 = (inp[0]) ? 3'b000 : 3'b001;

endmodule