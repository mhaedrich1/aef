module dtc_split125_bm82 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;

	assign outp = (inp[0]) ? node160 : node1;
		assign node1 = (inp[3]) ? node97 : node2;
			assign node2 = (inp[6]) ? node40 : node3;
				assign node3 = (inp[1]) ? node15 : node4;
					assign node4 = (inp[7]) ? node8 : node5;
						assign node5 = (inp[4]) ? 3'b111 : 3'b001;
						assign node8 = (inp[4]) ? node10 : 3'b111;
							assign node10 = (inp[10]) ? node12 : 3'b011;
								assign node12 = (inp[5]) ? 3'b111 : 3'b011;
					assign node15 = (inp[4]) ? node25 : node16;
						assign node16 = (inp[7]) ? node18 : 3'b001;
							assign node18 = (inp[9]) ? node22 : node19;
								assign node19 = (inp[2]) ? 3'b010 : 3'b001;
								assign node22 = (inp[11]) ? 3'b101 : 3'b011;
						assign node25 = (inp[8]) ? node33 : node26;
							assign node26 = (inp[5]) ? node30 : node27;
								assign node27 = (inp[7]) ? 3'b011 : 3'b111;
								assign node30 = (inp[10]) ? 3'b001 : 3'b001;
							assign node33 = (inp[10]) ? node37 : node34;
								assign node34 = (inp[7]) ? 3'b110 : 3'b101;
								assign node37 = (inp[5]) ? 3'b111 : 3'b001;
				assign node40 = (inp[9]) ? node70 : node41;
					assign node41 = (inp[1]) ? node57 : node42;
						assign node42 = (inp[4]) ? node50 : node43;
							assign node43 = (inp[11]) ? node47 : node44;
								assign node44 = (inp[10]) ? 3'b101 : 3'b100;
								assign node47 = (inp[7]) ? 3'b100 : 3'b110;
							assign node50 = (inp[10]) ? node54 : node51;
								assign node51 = (inp[7]) ? 3'b110 : 3'b001;
								assign node54 = (inp[8]) ? 3'b001 : 3'b011;
						assign node57 = (inp[4]) ? node65 : node58;
							assign node58 = (inp[10]) ? node62 : node59;
								assign node59 = (inp[2]) ? 3'b100 : 3'b000;
								assign node62 = (inp[7]) ? 3'b000 : 3'b100;
							assign node65 = (inp[7]) ? 3'b100 : node66;
								assign node66 = (inp[2]) ? 3'b100 : 3'b110;
					assign node70 = (inp[4]) ? node82 : node71;
						assign node71 = (inp[2]) ? node77 : node72;
							assign node72 = (inp[7]) ? 3'b010 : node73;
								assign node73 = (inp[1]) ? 3'b101 : 3'b011;
							assign node77 = (inp[5]) ? node79 : 3'b110;
								assign node79 = (inp[7]) ? 3'b100 : 3'b110;
						assign node82 = (inp[1]) ? node90 : node83;
							assign node83 = (inp[11]) ? node87 : node84;
								assign node84 = (inp[2]) ? 3'b011 : 3'b001;
								assign node87 = (inp[7]) ? 3'b001 : 3'b111;
							assign node90 = (inp[8]) ? node94 : node91;
								assign node91 = (inp[7]) ? 3'b001 : 3'b001;
								assign node94 = (inp[7]) ? 3'b010 : 3'b000;
			assign node97 = (inp[6]) ? node113 : node98;
				assign node98 = (inp[8]) ? node100 : 3'b111;
					assign node100 = (inp[2]) ? node102 : 3'b111;
						assign node102 = (inp[10]) ? node108 : node103;
							assign node103 = (inp[1]) ? 3'b001 : node104;
								assign node104 = (inp[11]) ? 3'b111 : 3'b011;
							assign node108 = (inp[11]) ? node110 : 3'b111;
								assign node110 = (inp[4]) ? 3'b111 : 3'b011;
				assign node113 = (inp[9]) ? node143 : node114;
					assign node114 = (inp[4]) ? node128 : node115;
						assign node115 = (inp[5]) ? node123 : node116;
							assign node116 = (inp[1]) ? node120 : node117;
								assign node117 = (inp[11]) ? 3'b001 : 3'b010;
								assign node120 = (inp[7]) ? 3'b110 : 3'b000;
							assign node123 = (inp[11]) ? 3'b001 : node124;
								assign node124 = (inp[8]) ? 3'b001 : 3'b101;
						assign node128 = (inp[1]) ? node136 : node129;
							assign node129 = (inp[2]) ? node133 : node130;
								assign node130 = (inp[10]) ? 3'b111 : 3'b011;
								assign node133 = (inp[11]) ? 3'b111 : 3'b101;
							assign node136 = (inp[10]) ? node140 : node137;
								assign node137 = (inp[2]) ? 3'b100 : 3'b101;
								assign node140 = (inp[7]) ? 3'b001 : 3'b011;
					assign node143 = (inp[1]) ? node149 : node144;
						assign node144 = (inp[7]) ? node146 : 3'b111;
							assign node146 = (inp[2]) ? 3'b101 : 3'b111;
						assign node149 = (inp[2]) ? node155 : node150;
							assign node150 = (inp[4]) ? node152 : 3'b011;
								assign node152 = (inp[11]) ? 3'b111 : 3'b111;
							assign node155 = (inp[10]) ? node157 : 3'b001;
								assign node157 = (inp[5]) ? 3'b011 : 3'b011;
		assign node160 = (inp[6]) ? node262 : node161;
			assign node161 = (inp[4]) ? node213 : node162;
				assign node162 = (inp[3]) ? node186 : node163;
					assign node163 = (inp[1]) ? node177 : node164;
						assign node164 = (inp[7]) ? node170 : node165;
							assign node165 = (inp[11]) ? 3'b001 : node166;
								assign node166 = (inp[5]) ? 3'b000 : 3'b001;
							assign node170 = (inp[10]) ? node174 : node171;
								assign node171 = (inp[5]) ? 3'b110 : 3'b100;
								assign node174 = (inp[2]) ? 3'b000 : 3'b010;
						assign node177 = (inp[7]) ? 3'b000 : node178;
							assign node178 = (inp[11]) ? node182 : node179;
								assign node179 = (inp[2]) ? 3'b000 : 3'b010;
								assign node182 = (inp[5]) ? 3'b110 : 3'b010;
					assign node186 = (inp[7]) ? node200 : node187;
						assign node187 = (inp[10]) ? node193 : node188;
							assign node188 = (inp[2]) ? 3'b101 : node189;
								assign node189 = (inp[9]) ? 3'b111 : 3'b101;
							assign node193 = (inp[2]) ? node197 : node194;
								assign node194 = (inp[9]) ? 3'b111 : 3'b011;
								assign node197 = (inp[5]) ? 3'b011 : 3'b110;
						assign node200 = (inp[5]) ? node206 : node201;
							assign node201 = (inp[10]) ? node203 : 3'b010;
								assign node203 = (inp[9]) ? 3'b001 : 3'b000;
							assign node206 = (inp[9]) ? node210 : node207;
								assign node207 = (inp[10]) ? 3'b110 : 3'b100;
								assign node210 = (inp[1]) ? 3'b001 : 3'b001;
				assign node213 = (inp[3]) ? node241 : node214;
					assign node214 = (inp[10]) ? node228 : node215;
						assign node215 = (inp[2]) ? node223 : node216;
							assign node216 = (inp[1]) ? node220 : node217;
								assign node217 = (inp[8]) ? 3'b010 : 3'b101;
								assign node220 = (inp[9]) ? 3'b010 : 3'b000;
							assign node223 = (inp[9]) ? node225 : 3'b100;
								assign node225 = (inp[5]) ? 3'b100 : 3'b110;
						assign node228 = (inp[9]) ? node236 : node229;
							assign node229 = (inp[7]) ? node233 : node230;
								assign node230 = (inp[1]) ? 3'b000 : 3'b101;
								assign node233 = (inp[11]) ? 3'b110 : 3'b010;
							assign node236 = (inp[2]) ? 3'b101 : node237;
								assign node237 = (inp[5]) ? 3'b111 : 3'b011;
					assign node241 = (inp[9]) ? node255 : node242;
						assign node242 = (inp[10]) ? node248 : node243;
							assign node243 = (inp[5]) ? node245 : 3'b001;
								assign node245 = (inp[1]) ? 3'b110 : 3'b011;
							assign node248 = (inp[7]) ? node252 : node249;
								assign node249 = (inp[1]) ? 3'b101 : 3'b111;
								assign node252 = (inp[1]) ? 3'b001 : 3'b101;
						assign node255 = (inp[1]) ? node257 : 3'b111;
							assign node257 = (inp[2]) ? 3'b011 : node258;
								assign node258 = (inp[7]) ? 3'b101 : 3'b011;
			assign node262 = (inp[3]) ? node294 : node263;
				assign node263 = (inp[4]) ? node273 : node264;
					assign node264 = (inp[1]) ? 3'b000 : node265;
						assign node265 = (inp[2]) ? node267 : 3'b000;
							assign node267 = (inp[7]) ? 3'b000 : node268;
								assign node268 = (inp[9]) ? 3'b010 : 3'b000;
					assign node273 = (inp[9]) ? node281 : node274;
						assign node274 = (inp[1]) ? 3'b000 : node275;
							assign node275 = (inp[11]) ? node277 : 3'b000;
								assign node277 = (inp[7]) ? 3'b000 : 3'b100;
						assign node281 = (inp[1]) ? node289 : node282;
							assign node282 = (inp[10]) ? node286 : node283;
								assign node283 = (inp[5]) ? 3'b000 : 3'b100;
								assign node286 = (inp[5]) ? 3'b010 : 3'b000;
							assign node289 = (inp[7]) ? 3'b000 : node290;
								assign node290 = (inp[10]) ? 3'b100 : 3'b000;
				assign node294 = (inp[9]) ? node320 : node295;
					assign node295 = (inp[1]) ? node311 : node296;
						assign node296 = (inp[2]) ? node304 : node297;
							assign node297 = (inp[5]) ? node301 : node298;
								assign node298 = (inp[8]) ? 3'b000 : 3'b010;
								assign node301 = (inp[8]) ? 3'b100 : 3'b001;
							assign node304 = (inp[5]) ? node308 : node305;
								assign node305 = (inp[10]) ? 3'b100 : 3'b000;
								assign node308 = (inp[4]) ? 3'b010 : 3'b100;
						assign node311 = (inp[7]) ? 3'b000 : node312;
							assign node312 = (inp[8]) ? node316 : node313;
								assign node313 = (inp[5]) ? 3'b010 : 3'b100;
								assign node316 = (inp[10]) ? 3'b100 : 3'b000;
					assign node320 = (inp[7]) ? node332 : node321;
						assign node321 = (inp[8]) ? node327 : node322;
							assign node322 = (inp[1]) ? 3'b110 : node323;
								assign node323 = (inp[11]) ? 3'b101 : 3'b001;
							assign node327 = (inp[11]) ? 3'b010 : node328;
								assign node328 = (inp[1]) ? 3'b100 : 3'b010;
						assign node332 = (inp[5]) ? node340 : node333;
							assign node333 = (inp[10]) ? node337 : node334;
								assign node334 = (inp[4]) ? 3'b010 : 3'b010;
								assign node337 = (inp[8]) ? 3'b100 : 3'b000;
							assign node340 = (inp[1]) ? node344 : node341;
								assign node341 = (inp[4]) ? 3'b100 : 3'b110;
								assign node344 = (inp[10]) ? 3'b110 : 3'b010;

endmodule