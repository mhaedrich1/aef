module dtc_split875_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node5;
	wire [40-1:0] node6;
	wire [40-1:0] node8;
	wire [40-1:0] node10;
	wire [40-1:0] node11;
	wire [40-1:0] node12;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node50;
	wire [40-1:0] node52;
	wire [40-1:0] node53;
	wire [40-1:0] node55;
	wire [40-1:0] node56;
	wire [40-1:0] node58;
	wire [40-1:0] node61;
	wire [40-1:0] node62;
	wire [40-1:0] node65;
	wire [40-1:0] node69;
	wire [40-1:0] node70;
	wire [40-1:0] node72;
	wire [40-1:0] node74;
	wire [40-1:0] node75;
	wire [40-1:0] node76;
	wire [40-1:0] node79;
	wire [40-1:0] node82;
	wire [40-1:0] node83;
	wire [40-1:0] node86;
	wire [40-1:0] node89;
	wire [40-1:0] node90;
	wire [40-1:0] node92;
	wire [40-1:0] node94;
	wire [40-1:0] node95;
	wire [40-1:0] node98;
	wire [40-1:0] node101;
	wire [40-1:0] node104;
	wire [40-1:0] node105;
	wire [40-1:0] node108;
	wire [40-1:0] node109;
	wire [40-1:0] node111;
	wire [40-1:0] node112;
	wire [40-1:0] node114;
	wire [40-1:0] node116;
	wire [40-1:0] node118;
	wire [40-1:0] node122;
	wire [40-1:0] node123;
	wire [40-1:0] node125;
	wire [40-1:0] node127;
	wire [40-1:0] node128;
	wire [40-1:0] node130;
	wire [40-1:0] node133;
	wire [40-1:0] node134;
	wire [40-1:0] node137;
	wire [40-1:0] node140;
	wire [40-1:0] node141;
	wire [40-1:0] node143;
	wire [40-1:0] node145;
	wire [40-1:0] node146;
	wire [40-1:0] node149;
	wire [40-1:0] node152;
	wire [40-1:0] node155;
	wire [40-1:0] node156;
	wire [40-1:0] node158;
	wire [40-1:0] node159;
	wire [40-1:0] node161;
	wire [40-1:0] node162;
	wire [40-1:0] node164;
	wire [40-1:0] node166;
	wire [40-1:0] node167;
	wire [40-1:0] node169;
	wire [40-1:0] node172;
	wire [40-1:0] node173;
	wire [40-1:0] node176;
	wire [40-1:0] node179;
	wire [40-1:0] node180;
	wire [40-1:0] node182;
	wire [40-1:0] node184;
	wire [40-1:0] node185;
	wire [40-1:0] node188;
	wire [40-1:0] node191;
	wire [40-1:0] node195;
	wire [40-1:0] node196;
	wire [40-1:0] node198;
	wire [40-1:0] node200;
	wire [40-1:0] node201;
	wire [40-1:0] node203;
	wire [40-1:0] node206;
	wire [40-1:0] node207;
	wire [40-1:0] node210;
	wire [40-1:0] node213;
	wire [40-1:0] node214;
	wire [40-1:0] node217;
	wire [40-1:0] node218;
	wire [40-1:0] node220;
	wire [40-1:0] node222;
	wire [40-1:0] node224;
	wire [40-1:0] node226;
	wire [40-1:0] node228;
	wire [40-1:0] node231;
	wire [40-1:0] node232;
	wire [40-1:0] node234;
	wire [40-1:0] node236;
	wire [40-1:0] node237;
	wire [40-1:0] node239;
	wire [40-1:0] node242;
	wire [40-1:0] node243;
	wire [40-1:0] node246;
	wire [40-1:0] node249;
	wire [40-1:0] node250;
	wire [40-1:0] node252;
	wire [40-1:0] node254;
	wire [40-1:0] node255;
	wire [40-1:0] node258;
	wire [40-1:0] node261;
	wire [40-1:0] node264;
	wire [40-1:0] node265;
	wire [40-1:0] node266;
	wire [40-1:0] node269;
	wire [40-1:0] node270;
	wire [40-1:0] node271;
	wire [40-1:0] node272;
	wire [40-1:0] node273;
	wire [40-1:0] node276;
	wire [40-1:0] node279;
	wire [40-1:0] node280;
	wire [40-1:0] node283;
	wire [40-1:0] node286;
	wire [40-1:0] node287;
	wire [40-1:0] node288;
	wire [40-1:0] node291;
	wire [40-1:0] node294;
	wire [40-1:0] node295;
	wire [40-1:0] node298;
	wire [40-1:0] node301;
	wire [40-1:0] node302;
	wire [40-1:0] node303;
	wire [40-1:0] node304;
	wire [40-1:0] node307;
	wire [40-1:0] node310;
	wire [40-1:0] node311;
	wire [40-1:0] node314;
	wire [40-1:0] node317;
	wire [40-1:0] node318;
	wire [40-1:0] node319;
	wire [40-1:0] node322;
	wire [40-1:0] node325;
	wire [40-1:0] node326;
	wire [40-1:0] node329;
	wire [40-1:0] node332;
	wire [40-1:0] node333;
	wire [40-1:0] node336;
	wire [40-1:0] node338;
	wire [40-1:0] node339;
	wire [40-1:0] node340;
	wire [40-1:0] node341;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node344;
	wire [40-1:0] node345;
	wire [40-1:0] node346;
	wire [40-1:0] node347;
	wire [40-1:0] node350;
	wire [40-1:0] node353;
	wire [40-1:0] node354;
	wire [40-1:0] node357;
	wire [40-1:0] node360;
	wire [40-1:0] node361;
	wire [40-1:0] node362;
	wire [40-1:0] node365;
	wire [40-1:0] node368;
	wire [40-1:0] node369;
	wire [40-1:0] node372;
	wire [40-1:0] node375;
	wire [40-1:0] node376;
	wire [40-1:0] node377;
	wire [40-1:0] node378;
	wire [40-1:0] node381;
	wire [40-1:0] node384;
	wire [40-1:0] node385;
	wire [40-1:0] node388;
	wire [40-1:0] node391;
	wire [40-1:0] node392;
	wire [40-1:0] node393;
	wire [40-1:0] node396;
	wire [40-1:0] node399;
	wire [40-1:0] node400;
	wire [40-1:0] node403;
	wire [40-1:0] node406;
	wire [40-1:0] node407;
	wire [40-1:0] node408;
	wire [40-1:0] node409;
	wire [40-1:0] node410;
	wire [40-1:0] node413;
	wire [40-1:0] node416;
	wire [40-1:0] node417;
	wire [40-1:0] node420;
	wire [40-1:0] node423;
	wire [40-1:0] node424;
	wire [40-1:0] node425;
	wire [40-1:0] node428;
	wire [40-1:0] node431;
	wire [40-1:0] node432;
	wire [40-1:0] node435;
	wire [40-1:0] node438;
	wire [40-1:0] node439;
	wire [40-1:0] node440;
	wire [40-1:0] node441;
	wire [40-1:0] node444;
	wire [40-1:0] node447;
	wire [40-1:0] node448;
	wire [40-1:0] node451;
	wire [40-1:0] node454;
	wire [40-1:0] node455;
	wire [40-1:0] node456;
	wire [40-1:0] node459;
	wire [40-1:0] node462;
	wire [40-1:0] node463;
	wire [40-1:0] node466;
	wire [40-1:0] node469;
	wire [40-1:0] node470;
	wire [40-1:0] node471;
	wire [40-1:0] node472;
	wire [40-1:0] node473;
	wire [40-1:0] node474;
	wire [40-1:0] node477;
	wire [40-1:0] node480;
	wire [40-1:0] node481;
	wire [40-1:0] node484;
	wire [40-1:0] node487;
	wire [40-1:0] node488;
	wire [40-1:0] node489;
	wire [40-1:0] node492;
	wire [40-1:0] node495;
	wire [40-1:0] node496;
	wire [40-1:0] node499;
	wire [40-1:0] node502;
	wire [40-1:0] node503;
	wire [40-1:0] node504;
	wire [40-1:0] node505;
	wire [40-1:0] node508;
	wire [40-1:0] node511;
	wire [40-1:0] node512;
	wire [40-1:0] node515;
	wire [40-1:0] node518;
	wire [40-1:0] node519;
	wire [40-1:0] node520;
	wire [40-1:0] node523;
	wire [40-1:0] node526;
	wire [40-1:0] node527;
	wire [40-1:0] node530;
	wire [40-1:0] node533;
	wire [40-1:0] node534;
	wire [40-1:0] node535;
	wire [40-1:0] node536;
	wire [40-1:0] node537;
	wire [40-1:0] node540;
	wire [40-1:0] node543;
	wire [40-1:0] node544;
	wire [40-1:0] node547;
	wire [40-1:0] node550;
	wire [40-1:0] node551;
	wire [40-1:0] node552;
	wire [40-1:0] node555;
	wire [40-1:0] node558;
	wire [40-1:0] node559;
	wire [40-1:0] node562;
	wire [40-1:0] node565;
	wire [40-1:0] node566;
	wire [40-1:0] node567;
	wire [40-1:0] node568;
	wire [40-1:0] node571;
	wire [40-1:0] node574;
	wire [40-1:0] node575;
	wire [40-1:0] node578;
	wire [40-1:0] node581;
	wire [40-1:0] node582;
	wire [40-1:0] node583;
	wire [40-1:0] node586;
	wire [40-1:0] node589;
	wire [40-1:0] node590;
	wire [40-1:0] node593;
	wire [40-1:0] node596;
	wire [40-1:0] node597;
	wire [40-1:0] node599;
	wire [40-1:0] node600;
	wire [40-1:0] node601;
	wire [40-1:0] node602;
	wire [40-1:0] node603;
	wire [40-1:0] node606;
	wire [40-1:0] node612;
	wire [40-1:0] node613;
	wire [40-1:0] node614;
	wire [40-1:0] node615;
	wire [40-1:0] node616;
	wire [40-1:0] node617;
	wire [40-1:0] node620;
	wire [40-1:0] node623;
	wire [40-1:0] node624;
	wire [40-1:0] node627;
	wire [40-1:0] node630;
	wire [40-1:0] node631;
	wire [40-1:0] node632;
	wire [40-1:0] node635;
	wire [40-1:0] node638;
	wire [40-1:0] node639;
	wire [40-1:0] node642;
	wire [40-1:0] node645;
	wire [40-1:0] node646;
	wire [40-1:0] node647;
	wire [40-1:0] node648;
	wire [40-1:0] node651;
	wire [40-1:0] node654;
	wire [40-1:0] node655;
	wire [40-1:0] node658;
	wire [40-1:0] node661;
	wire [40-1:0] node662;
	wire [40-1:0] node663;
	wire [40-1:0] node666;
	wire [40-1:0] node669;
	wire [40-1:0] node670;
	wire [40-1:0] node673;
	wire [40-1:0] node676;
	wire [40-1:0] node677;
	wire [40-1:0] node678;
	wire [40-1:0] node679;
	wire [40-1:0] node680;
	wire [40-1:0] node683;
	wire [40-1:0] node686;
	wire [40-1:0] node687;
	wire [40-1:0] node690;
	wire [40-1:0] node693;
	wire [40-1:0] node694;
	wire [40-1:0] node695;
	wire [40-1:0] node698;
	wire [40-1:0] node701;
	wire [40-1:0] node702;
	wire [40-1:0] node705;
	wire [40-1:0] node708;
	wire [40-1:0] node709;
	wire [40-1:0] node710;
	wire [40-1:0] node711;
	wire [40-1:0] node714;
	wire [40-1:0] node717;
	wire [40-1:0] node718;
	wire [40-1:0] node721;
	wire [40-1:0] node724;
	wire [40-1:0] node725;
	wire [40-1:0] node726;
	wire [40-1:0] node729;
	wire [40-1:0] node732;
	wire [40-1:0] node733;
	wire [40-1:0] node736;
	wire [40-1:0] node739;
	wire [40-1:0] node740;
	wire [40-1:0] node741;
	wire [40-1:0] node742;
	wire [40-1:0] node743;
	wire [40-1:0] node745;
	wire [40-1:0] node746;
	wire [40-1:0] node747;
	wire [40-1:0] node751;
	wire [40-1:0] node752;
	wire [40-1:0] node755;
	wire [40-1:0] node758;
	wire [40-1:0] node759;
	wire [40-1:0] node760;
	wire [40-1:0] node761;
	wire [40-1:0] node764;
	wire [40-1:0] node767;
	wire [40-1:0] node768;
	wire [40-1:0] node773;
	wire [40-1:0] node774;
	wire [40-1:0] node775;
	wire [40-1:0] node777;
	wire [40-1:0] node779;
	wire [40-1:0] node782;
	wire [40-1:0] node783;
	wire [40-1:0] node784;
	wire [40-1:0] node791;
	wire [40-1:0] node792;
	wire [40-1:0] node794;
	wire [40-1:0] node796;
	wire [40-1:0] node797;
	wire [40-1:0] node799;
	wire [40-1:0] node800;
	wire [40-1:0] node803;
	wire [40-1:0] node807;
	wire [40-1:0] node808;
	wire [40-1:0] node809;
	wire [40-1:0] node810;
	wire [40-1:0] node811;
	wire [40-1:0] node812;
	wire [40-1:0] node815;
	wire [40-1:0] node818;
	wire [40-1:0] node819;
	wire [40-1:0] node822;
	wire [40-1:0] node825;
	wire [40-1:0] node826;
	wire [40-1:0] node827;
	wire [40-1:0] node830;
	wire [40-1:0] node833;
	wire [40-1:0] node834;
	wire [40-1:0] node837;
	wire [40-1:0] node840;
	wire [40-1:0] node841;
	wire [40-1:0] node842;
	wire [40-1:0] node843;
	wire [40-1:0] node846;
	wire [40-1:0] node849;
	wire [40-1:0] node850;
	wire [40-1:0] node853;
	wire [40-1:0] node856;
	wire [40-1:0] node857;
	wire [40-1:0] node858;
	wire [40-1:0] node861;
	wire [40-1:0] node864;
	wire [40-1:0] node865;
	wire [40-1:0] node868;
	wire [40-1:0] node871;
	wire [40-1:0] node872;
	wire [40-1:0] node873;
	wire [40-1:0] node874;
	wire [40-1:0] node875;
	wire [40-1:0] node878;
	wire [40-1:0] node881;
	wire [40-1:0] node882;
	wire [40-1:0] node885;
	wire [40-1:0] node888;
	wire [40-1:0] node889;
	wire [40-1:0] node890;
	wire [40-1:0] node893;
	wire [40-1:0] node896;
	wire [40-1:0] node897;
	wire [40-1:0] node900;
	wire [40-1:0] node903;
	wire [40-1:0] node904;
	wire [40-1:0] node905;
	wire [40-1:0] node906;
	wire [40-1:0] node909;
	wire [40-1:0] node912;
	wire [40-1:0] node913;
	wire [40-1:0] node916;
	wire [40-1:0] node919;
	wire [40-1:0] node920;
	wire [40-1:0] node921;
	wire [40-1:0] node924;
	wire [40-1:0] node927;
	wire [40-1:0] node928;
	wire [40-1:0] node931;
	wire [40-1:0] node934;
	wire [40-1:0] node935;
	wire [40-1:0] node936;
	wire [40-1:0] node938;
	wire [40-1:0] node939;
	wire [40-1:0] node941;
	wire [40-1:0] node943;
	wire [40-1:0] node945;
	wire [40-1:0] node946;
	wire [40-1:0] node949;
	wire [40-1:0] node952;
	wire [40-1:0] node953;
	wire [40-1:0] node955;
	wire [40-1:0] node957;
	wire [40-1:0] node958;
	wire [40-1:0] node961;
	wire [40-1:0] node964;
	wire [40-1:0] node965;
	wire [40-1:0] node967;
	wire [40-1:0] node968;
	wire [40-1:0] node971;
	wire [40-1:0] node974;
	wire [40-1:0] node975;
	wire [40-1:0] node976;
	wire [40-1:0] node979;
	wire [40-1:0] node983;
	wire [40-1:0] node984;
	wire [40-1:0] node985;
	wire [40-1:0] node986;
	wire [40-1:0] node988;
	wire [40-1:0] node991;
	wire [40-1:0] node992;
	wire [40-1:0] node996;
	wire [40-1:0] node997;
	wire [40-1:0] node999;
	wire [40-1:0] node1002;
	wire [40-1:0] node1003;
	wire [40-1:0] node1008;
	wire [40-1:0] node1009;
	wire [40-1:0] node1011;
	wire [40-1:0] node1012;
	wire [40-1:0] node1013;
	wire [40-1:0] node1014;
	wire [40-1:0] node1015;
	wire [40-1:0] node1016;
	wire [40-1:0] node1019;
	wire [40-1:0] node1022;
	wire [40-1:0] node1023;
	wire [40-1:0] node1026;
	wire [40-1:0] node1029;
	wire [40-1:0] node1030;
	wire [40-1:0] node1031;
	wire [40-1:0] node1034;
	wire [40-1:0] node1037;
	wire [40-1:0] node1038;
	wire [40-1:0] node1041;
	wire [40-1:0] node1044;
	wire [40-1:0] node1045;
	wire [40-1:0] node1046;
	wire [40-1:0] node1047;
	wire [40-1:0] node1050;
	wire [40-1:0] node1053;
	wire [40-1:0] node1054;
	wire [40-1:0] node1057;
	wire [40-1:0] node1060;
	wire [40-1:0] node1061;
	wire [40-1:0] node1062;
	wire [40-1:0] node1065;
	wire [40-1:0] node1068;
	wire [40-1:0] node1069;
	wire [40-1:0] node1072;
	wire [40-1:0] node1075;
	wire [40-1:0] node1076;
	wire [40-1:0] node1077;
	wire [40-1:0] node1078;
	wire [40-1:0] node1079;
	wire [40-1:0] node1082;
	wire [40-1:0] node1085;
	wire [40-1:0] node1086;
	wire [40-1:0] node1089;
	wire [40-1:0] node1092;
	wire [40-1:0] node1093;
	wire [40-1:0] node1094;
	wire [40-1:0] node1097;
	wire [40-1:0] node1100;
	wire [40-1:0] node1101;
	wire [40-1:0] node1104;
	wire [40-1:0] node1107;
	wire [40-1:0] node1108;
	wire [40-1:0] node1109;
	wire [40-1:0] node1110;
	wire [40-1:0] node1113;
	wire [40-1:0] node1116;
	wire [40-1:0] node1117;
	wire [40-1:0] node1120;
	wire [40-1:0] node1123;
	wire [40-1:0] node1124;
	wire [40-1:0] node1125;
	wire [40-1:0] node1128;
	wire [40-1:0] node1131;
	wire [40-1:0] node1132;
	wire [40-1:0] node1135;
	wire [40-1:0] node1138;
	wire [40-1:0] node1139;
	wire [40-1:0] node1140;
	wire [40-1:0] node1141;
	wire [40-1:0] node1142;
	wire [40-1:0] node1143;
	wire [40-1:0] node1144;
	wire [40-1:0] node1147;
	wire [40-1:0] node1150;
	wire [40-1:0] node1151;
	wire [40-1:0] node1154;
	wire [40-1:0] node1157;
	wire [40-1:0] node1158;
	wire [40-1:0] node1159;
	wire [40-1:0] node1162;
	wire [40-1:0] node1165;
	wire [40-1:0] node1166;
	wire [40-1:0] node1169;
	wire [40-1:0] node1172;
	wire [40-1:0] node1173;
	wire [40-1:0] node1174;
	wire [40-1:0] node1175;
	wire [40-1:0] node1178;
	wire [40-1:0] node1181;
	wire [40-1:0] node1182;
	wire [40-1:0] node1185;
	wire [40-1:0] node1188;
	wire [40-1:0] node1189;
	wire [40-1:0] node1190;
	wire [40-1:0] node1193;
	wire [40-1:0] node1196;
	wire [40-1:0] node1197;
	wire [40-1:0] node1200;
	wire [40-1:0] node1203;
	wire [40-1:0] node1204;
	wire [40-1:0] node1205;
	wire [40-1:0] node1206;
	wire [40-1:0] node1207;
	wire [40-1:0] node1210;
	wire [40-1:0] node1213;
	wire [40-1:0] node1214;
	wire [40-1:0] node1217;
	wire [40-1:0] node1220;
	wire [40-1:0] node1221;
	wire [40-1:0] node1222;
	wire [40-1:0] node1225;
	wire [40-1:0] node1228;
	wire [40-1:0] node1229;
	wire [40-1:0] node1232;
	wire [40-1:0] node1235;
	wire [40-1:0] node1236;
	wire [40-1:0] node1237;
	wire [40-1:0] node1238;
	wire [40-1:0] node1241;
	wire [40-1:0] node1244;
	wire [40-1:0] node1245;
	wire [40-1:0] node1248;
	wire [40-1:0] node1251;
	wire [40-1:0] node1252;
	wire [40-1:0] node1253;
	wire [40-1:0] node1256;
	wire [40-1:0] node1259;
	wire [40-1:0] node1260;
	wire [40-1:0] node1263;

	assign outp = (inp[9]) ? node264 : node1;
		assign node1 = (inp[4]) ? node5 : node2;
			assign node2 = (inp[1]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
			assign node5 = (inp[1]) ? node17 : node6;
				assign node6 = (inp[8]) ? node8 : 40'b0000000000000000000000000000000000000000;
					assign node8 = (inp[7]) ? node10 : 40'b0000000000000000000000000000000000000000;
						assign node10 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node11;
							assign node11 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node12;
								assign node12 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
				assign node17 = (inp[7]) ? node155 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[11]) ? node24 : node21;
								assign node21 = (inp[3]) ? 40'b0000000000100010000000000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[3]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000000010000001000000000000000000;
							assign node27 = (inp[11]) ? node31 : node28;
								assign node28 = (inp[3]) ? 40'b0000000000100000000000000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[3]) ? node33 : 40'b0000000000000000000001000000000010000000;
									assign node33 = (inp[10]) ? node39 : node34;
										assign node34 = (inp[0]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[13]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[13]) ? node43 : node40;
											assign node40 = (inp[0]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000010000000;
						assign node46 = (inp[14]) ? node104 : node47;
							assign node47 = (inp[0]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[3]) ? node69 : node50;
									assign node50 = (inp[15]) ? node52 : 40'b0000000000000000000000000000000000000000;
										assign node52 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node53;
											assign node53 = (inp[12]) ? node55 : 40'b0000000000000000000000000000000000000000;
												assign node55 = (inp[2]) ? node61 : node56;
													assign node56 = (inp[6]) ? node58 : 40'b0000000000000000000000000000000000000000;
														assign node58 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node61 = (inp[10]) ? node65 : node62;
														assign node62 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node65 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node69 = (inp[13]) ? node89 : node70;
										assign node70 = (inp[12]) ? node72 : 40'b0000000000000000000000000000000000000000;
											assign node72 = (inp[15]) ? node74 : 40'b0000000000000000000000000000000000000000;
												assign node74 = (inp[10]) ? node82 : node75;
													assign node75 = (inp[6]) ? node79 : node76;
														assign node76 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node79 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node82 = (inp[5]) ? node86 : node83;
														assign node83 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node86 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node89 = (inp[10]) ? node101 : node90;
											assign node90 = (inp[15]) ? node92 : 40'b0000000000000000000000000000000000000000;
												assign node92 = (inp[12]) ? node94 : 40'b0000000000000000000000000000000000000000;
													assign node94 = (inp[5]) ? node98 : node95;
														assign node95 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node98 = (inp[11]) ? 40'b0000000000000010010000100000010000000000 : 40'b0000000000000000000000000000000000000000;
											assign node101 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000001000000000;
							assign node104 = (inp[3]) ? node108 : node105;
								assign node105 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node108 = (inp[0]) ? node122 : node109;
									assign node109 = (inp[5]) ? node111 : 40'b0000000000000000000000000000000000000000;
										assign node111 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node112;
											assign node112 = (inp[15]) ? node114 : 40'b0000000000000000000000000000000000000000;
												assign node114 = (inp[12]) ? node116 : 40'b0000000000000000000000000000000000000000;
													assign node116 = (inp[6]) ? node118 : 40'b0000000000000000000000000000000000000000;
														assign node118 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node122 = (inp[10]) ? node140 : node123;
										assign node123 = (inp[15]) ? node125 : 40'b0000000000000000000000000000000000000000;
											assign node125 = (inp[12]) ? node127 : 40'b0000000000000000000000000000000000000000;
												assign node127 = (inp[5]) ? node133 : node128;
													assign node128 = (inp[6]) ? node130 : 40'b0000000000000000000000000000000000000000;
														assign node130 = (inp[2]) ? 40'b0000000000000000010000000000000001000010 : 40'b0000000000000000000000000000000000000000;
													assign node133 = (inp[13]) ? node137 : node134;
														assign node134 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node137 = (inp[2]) ? 40'b0000000000000010010000100000001001000000 : 40'b0000000010000010010000100000000001000000;
										assign node140 = (inp[13]) ? node152 : node141;
											assign node141 = (inp[15]) ? node143 : 40'b0000000000000000000000000000000000000000;
												assign node143 = (inp[12]) ? node145 : 40'b0000000000000000000000000000000000000000;
													assign node145 = (inp[6]) ? node149 : node146;
														assign node146 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node149 = (inp[11]) ? 40'b0000000000001000010000100000000011000000 : 40'b0000000000000000010100100000000011000000;
											assign node152 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node155 = (inp[14]) ? node195 : node156;
						assign node156 = (inp[8]) ? node158 : 40'b0000000000000000000000000000000000000000;
							assign node158 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node159;
								assign node159 = (inp[0]) ? node161 : 40'b0000000000000000000000000000000000000000;
									assign node161 = (inp[13]) ? node179 : node162;
										assign node162 = (inp[12]) ? node164 : 40'b0000000000000000000000000000000000000000;
											assign node164 = (inp[15]) ? node166 : 40'b0000000000000000000000000000000000000000;
												assign node166 = (inp[5]) ? node172 : node167;
													assign node167 = (inp[6]) ? node169 : 40'b0000000000000000000000000000000000000000;
														assign node169 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node172 = (inp[10]) ? node176 : node173;
														assign node173 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node176 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node179 = (inp[10]) ? node191 : node180;
											assign node180 = (inp[15]) ? node182 : 40'b0000000000000000000000000000000000000000;
												assign node182 = (inp[12]) ? node184 : 40'b0000000000000000000000000000000000000000;
													assign node184 = (inp[5]) ? node188 : node185;
														assign node185 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node188 = (inp[6]) ? 40'b0000000010000010000000100000000100000000 : 40'b0000000000000000000000000000000000000000;
											assign node191 = (inp[3]) ? 40'b0000000000000000000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
						assign node195 = (inp[8]) ? node213 : node196;
							assign node196 = (inp[11]) ? node198 : 40'b0000000000000000000000000000000000000000;
								assign node198 = (inp[3]) ? node200 : 40'b0000000000000000000000000000000000000000;
									assign node200 = (inp[10]) ? node206 : node201;
										assign node201 = (inp[0]) ? node203 : 40'b0000000000000000000000000000000000000000;
											assign node203 = (inp[13]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node206 = (inp[0]) ? node210 : node207;
											assign node207 = (inp[13]) ? 40'b0000000000000010000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node210 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000010000000110000000;
							assign node213 = (inp[3]) ? node217 : node214;
								assign node214 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node217 = (inp[0]) ? node231 : node218;
									assign node218 = (inp[6]) ? node220 : 40'b0000000000000000000000000000000000000000;
										assign node220 = (inp[12]) ? node222 : 40'b0000000000000000000000000000000000000000;
											assign node222 = (inp[5]) ? node224 : 40'b0000000000000000000000000000000000000000;
												assign node224 = (inp[15]) ? node226 : 40'b0000000000000000000000000000000000000000;
													assign node226 = (inp[2]) ? node228 : 40'b0000000000000000000000000000000000000000;
														assign node228 = (inp[10]) ? 40'b0100000000000000000000001000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node231 = (inp[13]) ? node249 : node232;
										assign node232 = (inp[15]) ? node234 : 40'b0000000000000000000000000000000000000000;
											assign node234 = (inp[12]) ? node236 : 40'b0000000000000000000000000000000000000000;
												assign node236 = (inp[2]) ? node242 : node237;
													assign node237 = (inp[5]) ? node239 : 40'b0000000000000000000000000000000000000000;
														assign node239 = (inp[6]) ? 40'b0100000010000000000000000000000100000000 : 40'b0000000000000000000000000000000000000000;
													assign node242 = (inp[10]) ? node246 : node243;
														assign node243 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node246 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node249 = (inp[10]) ? node261 : node250;
											assign node250 = (inp[15]) ? node252 : 40'b0000000000000000000000000000000000000000;
												assign node252 = (inp[12]) ? node254 : 40'b0000000000000000000000000000000000000000;
													assign node254 = (inp[6]) ? node258 : node255;
														assign node255 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node258 = (inp[11]) ? 40'b0100000000000010000000100000000100000001 : 40'b0000000000000000000000000000000000000000;
											assign node261 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node264 = (inp[1]) ? node332 : node265;
			assign node265 = (inp[8]) ? node269 : node266;
				assign node266 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node269 = (inp[7]) ? node301 : node270;
					assign node270 = (inp[11]) ? node286 : node271;
						assign node271 = (inp[3]) ? node279 : node272;
							assign node272 = (inp[14]) ? node276 : node273;
								assign node273 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node276 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
							assign node279 = (inp[14]) ? node283 : node280;
								assign node280 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node283 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
						assign node286 = (inp[14]) ? node294 : node287;
							assign node287 = (inp[3]) ? node291 : node288;
								assign node288 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node291 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
							assign node294 = (inp[3]) ? node298 : node295;
								assign node295 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
								assign node298 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node301 = (inp[14]) ? node317 : node302;
						assign node302 = (inp[3]) ? node310 : node303;
							assign node303 = (inp[11]) ? node307 : node304;
								assign node304 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node307 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
							assign node310 = (inp[11]) ? node314 : node311;
								assign node311 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node314 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
						assign node317 = (inp[3]) ? node325 : node318;
							assign node318 = (inp[11]) ? node322 : node319;
								assign node319 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node322 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
							assign node325 = (inp[11]) ? node329 : node326;
								assign node326 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
								assign node329 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node332 = (inp[4]) ? node336 : node333;
				assign node333 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node336 = (inp[8]) ? node338 : 40'b0000100000000000000000000000000000000000;
					assign node338 = (inp[7]) ? node934 : node339;
						assign node339 = (inp[3]) ? node739 : node340;
							assign node340 = (inp[14]) ? node596 : node341;
								assign node341 = (inp[11]) ? node469 : node342;
									assign node342 = (inp[13]) ? node406 : node343;
										assign node343 = (inp[10]) ? node375 : node344;
											assign node344 = (inp[15]) ? node360 : node345;
												assign node345 = (inp[0]) ? node353 : node346;
													assign node346 = (inp[5]) ? node350 : node347;
														assign node347 = (inp[6]) ? 40'b0001000000011101010010000010101000010000 : 40'b1001000000010101010010000000101000010000;
														assign node350 = (inp[6]) ? 40'b0001000000010101010010000001101000010000 : 40'b0001000000010101010110000010101000010000;
													assign node353 = (inp[2]) ? node357 : node354;
														assign node354 = (inp[12]) ? 40'b0000000000011101010010000010101000010000 : 40'b1000000000010101010010000000101000010000;
														assign node357 = (inp[12]) ? 40'b0000000000010101010010000001101000010000 : 40'b0000000000010101010110000010101000010000;
												assign node360 = (inp[0]) ? node368 : node361;
													assign node361 = (inp[5]) ? node365 : node362;
														assign node362 = (inp[6]) ? 40'b0001000000001101010010000010101000010000 : 40'b1001000000000101010010000000101000010000;
														assign node365 = (inp[6]) ? 40'b0001000000000101010010000001101000010000 : 40'b0001000000000101010110000010101000010000;
													assign node368 = (inp[6]) ? node372 : node369;
														assign node369 = (inp[5]) ? 40'b0000000000000101010110000010101000010000 : 40'b1000000000000101010010000000101000010000;
														assign node372 = (inp[5]) ? 40'b0000000000000101010010000001101000010000 : 40'b0000000000001101010010000010101000010000;
											assign node375 = (inp[0]) ? node391 : node376;
												assign node376 = (inp[15]) ? node384 : node377;
													assign node377 = (inp[12]) ? node381 : node378;
														assign node378 = (inp[2]) ? 40'b0001000000010001010110000010101000010000 : 40'b1001000000010001010010000000101000010000;
														assign node381 = (inp[6]) ? 40'b0001000000011001010010000011101000010000 : 40'b0001000000010001010010000001101000010000;
													assign node384 = (inp[12]) ? node388 : node385;
														assign node385 = (inp[2]) ? 40'b0001000000000001010110000010101000010000 : 40'b1001000000000001010010000010101000010000;
														assign node388 = (inp[2]) ? 40'b0001000000000001010010000001101000010000 : 40'b0001000000001001010010000010101000010000;
												assign node391 = (inp[15]) ? node399 : node392;
													assign node392 = (inp[5]) ? node396 : node393;
														assign node393 = (inp[6]) ? 40'b0000000000011001010010000010101000010000 : 40'b1000000000010001010010000000101000010000;
														assign node396 = (inp[6]) ? 40'b0000000000010001010010000001101000010000 : 40'b0000000000010001010110000010101000010000;
													assign node399 = (inp[5]) ? node403 : node400;
														assign node400 = (inp[6]) ? 40'b0000000000001001010010000010101000010000 : 40'b1000000000000001010010000000101000010000;
														assign node403 = (inp[6]) ? 40'b0000000000000001010010000001101000010000 : 40'b0000000000000001010110000010101000010000;
										assign node406 = (inp[0]) ? node438 : node407;
											assign node407 = (inp[10]) ? node423 : node408;
												assign node408 = (inp[15]) ? node416 : node409;
													assign node409 = (inp[6]) ? node413 : node410;
														assign node410 = (inp[5]) ? 40'b0001000000010101010110000010001000010000 : 40'b1001000000010101010010000010001000010000;
														assign node413 = (inp[5]) ? 40'b0001000000010101010010000001001000010000 : 40'b0001000000011101010010000010001000010000;
													assign node416 = (inp[12]) ? node420 : node417;
														assign node417 = (inp[2]) ? 40'b0001000000000101010110000010001000010000 : 40'b1001000000000101010010000000001000010000;
														assign node420 = (inp[2]) ? 40'b0001000000000101010010000001001000010000 : 40'b0001000000001101010010000010001000010000;
												assign node423 = (inp[15]) ? node431 : node424;
													assign node424 = (inp[6]) ? node428 : node425;
														assign node425 = (inp[5]) ? 40'b0001000000010001010110000010001000010000 : 40'b1001000000010001010010000000001000010000;
														assign node428 = (inp[5]) ? 40'b0001000000010001010010000001001000010000 : 40'b0001000000011001010010000010001000010000;
													assign node431 = (inp[5]) ? node435 : node432;
														assign node432 = (inp[6]) ? 40'b0001000000001001010010000010001000010000 : 40'b1001000000000001010010000010001000010000;
														assign node435 = (inp[6]) ? 40'b0001000000000001010010000001001000010000 : 40'b0001000000000001010110000010001000010000;
											assign node438 = (inp[15]) ? node454 : node439;
												assign node439 = (inp[10]) ? node447 : node440;
													assign node440 = (inp[5]) ? node444 : node441;
														assign node441 = (inp[6]) ? 40'b0000000000011101010010000010001000010000 : 40'b1000000000010101010010000000001000010000;
														assign node444 = (inp[6]) ? 40'b0000000000010101010010000001001000010000 : 40'b0000000000010101010110000010001000010000;
													assign node447 = (inp[5]) ? node451 : node448;
														assign node448 = (inp[6]) ? 40'b0000000000011001010010000010001000010000 : 40'b1000000000010001010010000000001000010000;
														assign node451 = (inp[6]) ? 40'b0000000000010001010010000001001000010000 : 40'b0000000000010001010110000010001000010000;
												assign node454 = (inp[10]) ? node462 : node455;
													assign node455 = (inp[5]) ? node459 : node456;
														assign node456 = (inp[6]) ? 40'b0000000000001101010010000010001000010000 : 40'b1000000000000101010010000000001000010000;
														assign node459 = (inp[6]) ? 40'b1000000000000101010010000001001000010000 : 40'b0000000000000101010110000010001000010000;
													assign node462 = (inp[12]) ? node466 : node463;
														assign node463 = (inp[2]) ? 40'b0000000000000001010110000010001000010000 : 40'b1000000000000001010010000000001000010000;
														assign node466 = (inp[2]) ? 40'b0000000000000001010010000001001000010000 : 40'b0000000000001001010010000010001000010000;
									assign node469 = (inp[13]) ? node533 : node470;
										assign node470 = (inp[15]) ? node502 : node471;
											assign node471 = (inp[0]) ? node487 : node472;
												assign node472 = (inp[10]) ? node480 : node473;
													assign node473 = (inp[6]) ? node477 : node474;
														assign node474 = (inp[12]) ? 40'b0001000000010101010110000010101000000000 : 40'b1001000000010101010110000010101000000000;
														assign node477 = (inp[5]) ? 40'b0001000000010101010010000001101000000000 : 40'b0001000000011101010010000010101000000000;
													assign node480 = (inp[12]) ? node484 : node481;
														assign node481 = (inp[2]) ? 40'b0001000000010001010110000010101000000000 : 40'b1001000000010001010010000000101000000000;
														assign node484 = (inp[2]) ? 40'b0001000000010001010010000001101000000000 : 40'b0001000000011001010010000010101000000000;
												assign node487 = (inp[10]) ? node495 : node488;
													assign node488 = (inp[2]) ? node492 : node489;
														assign node489 = (inp[12]) ? 40'b0000000000011101010010000010101000000000 : 40'b1000000000010101010010000000101000000000;
														assign node492 = (inp[12]) ? 40'b0000000000010101010010000001101000000000 : 40'b0000000000010101010110000010101000000000;
													assign node495 = (inp[12]) ? node499 : node496;
														assign node496 = (inp[2]) ? 40'b0000000000010001010110000010101000000000 : 40'b1000000000010001010010000000101000000000;
														assign node499 = (inp[2]) ? 40'b0000000000010001010010000001101000000000 : 40'b0000000000011001010010000010101000000000;
											assign node502 = (inp[0]) ? node518 : node503;
												assign node503 = (inp[10]) ? node511 : node504;
													assign node504 = (inp[12]) ? node508 : node505;
														assign node505 = (inp[6]) ? 40'b0001000000001101010010000010101000000000 : 40'b1001000000000101010110000010101000000000;
														assign node508 = (inp[2]) ? 40'b0001000000000101010010000011101000000000 : 40'b0001000000001101010010000010101000000000;
													assign node511 = (inp[6]) ? node515 : node512;
														assign node512 = (inp[5]) ? 40'b0001000000000001010110000010101000000000 : 40'b1001000000000001010010000000101000000000;
														assign node515 = (inp[5]) ? 40'b0001000000000001010010000001101000000000 : 40'b0001000000001001010010000010101000000000;
												assign node518 = (inp[10]) ? node526 : node519;
													assign node519 = (inp[2]) ? node523 : node520;
														assign node520 = (inp[12]) ? 40'b0000000000001101010010000010101000000000 : 40'b1000000000000101010010000000101000000000;
														assign node523 = (inp[12]) ? 40'b0000000000000101010010000001101000000000 : 40'b0000000000000101010110000010101000000000;
													assign node526 = (inp[5]) ? node530 : node527;
														assign node527 = (inp[6]) ? 40'b0000000000001001010010000010101000000000 : 40'b1000000000000001010010000000101000000000;
														assign node530 = (inp[6]) ? 40'b0000000000000001010010000001101000000000 : 40'b0000000000000001010110000010101000000000;
										assign node533 = (inp[15]) ? node565 : node534;
											assign node534 = (inp[0]) ? node550 : node535;
												assign node535 = (inp[10]) ? node543 : node536;
													assign node536 = (inp[6]) ? node540 : node537;
														assign node537 = (inp[5]) ? 40'b0001000000010101010110000010001000000000 : 40'b1001000000010101010010000000001000000000;
														assign node540 = (inp[5]) ? 40'b0001000000010101010010000001001000000000 : 40'b0001000000011101010010000010001000000000;
													assign node543 = (inp[5]) ? node547 : node544;
														assign node544 = (inp[6]) ? 40'b0001000000011001010010000010001000000000 : 40'b1001000000010001010010000000001000000000;
														assign node547 = (inp[6]) ? 40'b0001000000010001010010000001001000000000 : 40'b0001000000010001010110000010001000000000;
												assign node550 = (inp[10]) ? node558 : node551;
													assign node551 = (inp[2]) ? node555 : node552;
														assign node552 = (inp[12]) ? 40'b0000000000011101010010000010001000000000 : 40'b1000000000010101010010000000001000000000;
														assign node555 = (inp[5]) ? 40'b0000000000010101010110000011001000000000 : 40'b0000000000011101010010000010001000000000;
													assign node558 = (inp[6]) ? node562 : node559;
														assign node559 = (inp[5]) ? 40'b0000000000010001010110000010001000000000 : 40'b1000000000010001010010000000001000000000;
														assign node562 = (inp[5]) ? 40'b0000000000010001010010000011001000000000 : 40'b0000000000011001010010000010001000000000;
											assign node565 = (inp[0]) ? node581 : node566;
												assign node566 = (inp[10]) ? node574 : node567;
													assign node567 = (inp[5]) ? node571 : node568;
														assign node568 = (inp[6]) ? 40'b0001000000001101010010000010001000000000 : 40'b1001000000000101010010000000001000000000;
														assign node571 = (inp[6]) ? 40'b0001000000000101010010000011001000000000 : 40'b0001000000000101010110000010001000000000;
													assign node574 = (inp[5]) ? node578 : node575;
														assign node575 = (inp[6]) ? 40'b0001000000001001010010000010001000000000 : 40'b1001000000000001010010000000001000000000;
														assign node578 = (inp[6]) ? 40'b0001000000000001010010000001001000000000 : 40'b0001000000000001010110000010001000000000;
												assign node581 = (inp[10]) ? node589 : node582;
													assign node582 = (inp[12]) ? node586 : node583;
														assign node583 = (inp[2]) ? 40'b0000000000000101010110000010001000000000 : 40'b1000000000000101010010000000001000000000;
														assign node586 = (inp[2]) ? 40'b0000000000000101010010000001001000000000 : 40'b0000000000001101010010000010001000000000;
													assign node589 = (inp[12]) ? node593 : node590;
														assign node590 = (inp[2]) ? 40'b0000000000000001010110000010001000000000 : 40'b1000000000000001010010000000001000000000;
														assign node593 = (inp[2]) ? 40'b0000000000000001010010000001001000000000 : 40'b0000000000001001010010000010001000000000;
								assign node596 = (inp[11]) ? node612 : node597;
									assign node597 = (inp[2]) ? node599 : 40'b0000000000000000000000000000000000000000;
										assign node599 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node600;
											assign node600 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node601;
												assign node601 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node602;
													assign node602 = (inp[15]) ? node606 : node603;
														assign node603 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node606 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node612 = (inp[0]) ? node676 : node613;
										assign node613 = (inp[13]) ? node645 : node614;
											assign node614 = (inp[10]) ? node630 : node615;
												assign node615 = (inp[15]) ? node623 : node616;
													assign node616 = (inp[2]) ? node620 : node617;
														assign node617 = (inp[12]) ? 40'b0001010000011100000000000010100000000000 : 40'b1001010000010100000000000000100000000000;
														assign node620 = (inp[12]) ? 40'b0001010000010100000000000001100000000000 : 40'b0001010000010100000100000010100000000000;
													assign node623 = (inp[2]) ? node627 : node624;
														assign node624 = (inp[12]) ? 40'b0001010000001100000000000010100000000000 : 40'b1001010000000100000000000010100000000000;
														assign node627 = (inp[12]) ? 40'b0001010000000100000000000001100000000000 : 40'b0001010000000100000100000010100000000000;
												assign node630 = (inp[15]) ? node638 : node631;
													assign node631 = (inp[12]) ? node635 : node632;
														assign node632 = (inp[2]) ? 40'b0001010000010000000100000010100000000000 : 40'b1001010000010000000000000000100000000000;
														assign node635 = (inp[2]) ? 40'b0001010000010000000000000001100000000000 : 40'b0001010000011000000000000010100000000000;
													assign node638 = (inp[5]) ? node642 : node639;
														assign node639 = (inp[6]) ? 40'b0001010000001000000000000010100000000000 : 40'b1001010000000000000000000000100000000000;
														assign node642 = (inp[6]) ? 40'b0001010000000000000000000001100000000000 : 40'b0001010000000000000100000010100000000000;
											assign node645 = (inp[15]) ? node661 : node646;
												assign node646 = (inp[10]) ? node654 : node647;
													assign node647 = (inp[5]) ? node651 : node648;
														assign node648 = (inp[6]) ? 40'b0001010000011100000000000010000000000000 : 40'b1001010000010100000000000000000000000000;
														assign node651 = (inp[6]) ? 40'b0001010000010100000000000001000000000000 : 40'b0001010000010100000100000010000000000000;
													assign node654 = (inp[2]) ? node658 : node655;
														assign node655 = (inp[12]) ? 40'b0001010000011000000000000010000000000000 : 40'b1001010000010000000000000000000000000000;
														assign node658 = (inp[12]) ? 40'b0001010000010000000000000001000000000000 : 40'b0001010000010000000100000010000000000000;
												assign node661 = (inp[10]) ? node669 : node662;
													assign node662 = (inp[2]) ? node666 : node663;
														assign node663 = (inp[12]) ? 40'b0001010000001100000000000010000000000000 : 40'b1001010000000100000000000010000000000000;
														assign node666 = (inp[12]) ? 40'b0001010000000100000000000011000000000000 : 40'b0001010000000100000100000010000000000000;
													assign node669 = (inp[6]) ? node673 : node670;
														assign node670 = (inp[5]) ? 40'b0001010000000000000100000010000000000000 : 40'b1001010000000000000000000000000000000000;
														assign node673 = (inp[5]) ? 40'b0001010000000000000000000001000000000000 : 40'b0001010000001000000000000010000000000000;
										assign node676 = (inp[13]) ? node708 : node677;
											assign node677 = (inp[10]) ? node693 : node678;
												assign node678 = (inp[15]) ? node686 : node679;
													assign node679 = (inp[12]) ? node683 : node680;
														assign node680 = (inp[2]) ? 40'b0000010000010100000100000010100000000000 : 40'b1000010000010100000000000010100000000000;
														assign node683 = (inp[2]) ? 40'b0000010000010100000000000001100000000000 : 40'b0000010000011100000000000010100000000000;
													assign node686 = (inp[5]) ? node690 : node687;
														assign node687 = (inp[6]) ? 40'b0000010000001100000000000010100000000000 : 40'b1000010000000100000000000000100000000000;
														assign node690 = (inp[2]) ? 40'b0000010000000100000100000011100000000000 : 40'b0000010000000100000100000010100000000000;
												assign node693 = (inp[15]) ? node701 : node694;
													assign node694 = (inp[5]) ? node698 : node695;
														assign node695 = (inp[6]) ? 40'b0000010000011000000000000010100000000000 : 40'b1000010000010000000000000000100000000000;
														assign node698 = (inp[6]) ? 40'b0000010000010000000000000001100000000000 : 40'b0000010000010000000100000010100000000000;
													assign node701 = (inp[6]) ? node705 : node702;
														assign node702 = (inp[5]) ? 40'b0000010000000000000100000010100000000000 : 40'b1000010000000000000000000000100000000000;
														assign node705 = (inp[5]) ? 40'b0000010000000000000000000001100000000000 : 40'b0000010000001000000000000010100000000000;
											assign node708 = (inp[10]) ? node724 : node709;
												assign node709 = (inp[15]) ? node717 : node710;
													assign node710 = (inp[6]) ? node714 : node711;
														assign node711 = (inp[5]) ? 40'b0000010000010100000100000010000000000000 : 40'b1000010000010100000000000000000000000000;
														assign node714 = (inp[5]) ? 40'b0000010000010100000000000001000000000000 : 40'b0000010000011100000000000010000000000000;
													assign node717 = (inp[6]) ? node721 : node718;
														assign node718 = (inp[5]) ? 40'b0000010000000100000100000010000000000000 : 40'b1000010000000100000000000000000000000000;
														assign node721 = (inp[5]) ? 40'b0000010000000100000000000001000000000000 : 40'b0000010000001100000000000010000000000000;
												assign node724 = (inp[15]) ? node732 : node725;
													assign node725 = (inp[5]) ? node729 : node726;
														assign node726 = (inp[6]) ? 40'b0000010000011000000000000010000000000000 : 40'b1000010000010000000000000010000000000000;
														assign node729 = (inp[6]) ? 40'b0000010000010000000000000001000000000000 : 40'b0000010000010000000100000010000000000000;
													assign node732 = (inp[12]) ? node736 : node733;
														assign node733 = (inp[2]) ? 40'b0000010000000000000100000010000000000000 : 40'b1000010000000000000000000000000000000000;
														assign node736 = (inp[2]) ? 40'b0000010000000000000000000001000000000000 : 40'b0000010000001000000000000010000000000000;
							assign node739 = (inp[11]) ? node791 : node740;
								assign node740 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node741;
									assign node741 = (inp[12]) ? node773 : node742;
										assign node742 = (inp[13]) ? node758 : node743;
											assign node743 = (inp[15]) ? node745 : 40'b0000000000000000000000000000000000000000;
												assign node745 = (inp[2]) ? node751 : node746;
													assign node746 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node747;
														assign node747 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node751 = (inp[5]) ? node755 : node752;
														assign node752 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node755 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000100000010100000100000;
											assign node758 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node759;
												assign node759 = (inp[2]) ? node767 : node760;
													assign node760 = (inp[0]) ? node764 : node761;
														assign node761 = (inp[10]) ? 40'b1001000000010000000000000000000000100000 : 40'b0000000000000000000000000000000000000000;
														assign node764 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100000000000010000000100000;
													assign node767 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node768;
														assign node768 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node773 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node774;
											assign node774 = (inp[13]) ? node782 : node775;
												assign node775 = (inp[15]) ? node777 : 40'b0000000000000000000000000000000000000000;
													assign node777 = (inp[5]) ? node779 : 40'b0000000000000000000000000000000000000000;
														assign node779 = (inp[2]) ? 40'b0000000000000000000100000011100000100000 : 40'b0000000000000000000000000000000000000000;
												assign node782 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node783;
													assign node783 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node784;
														assign node784 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000011000000000000010000000100000;
								assign node791 = (inp[14]) ? node807 : node792;
									assign node792 = (inp[12]) ? node794 : 40'b0000000000000000000000000000000000000000;
										assign node794 = (inp[5]) ? node796 : 40'b0000000000000000000000000000000000000000;
											assign node796 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node797;
												assign node797 = (inp[2]) ? node799 : 40'b0000000000000000000000000000000000000000;
													assign node799 = (inp[15]) ? node803 : node800;
														assign node800 = (inp[10]) ? 40'b1001000000010000001000000000000000010000 : 40'b0000000000000000000000000000000000000000;
														assign node803 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node807 = (inp[13]) ? node871 : node808;
										assign node808 = (inp[10]) ? node840 : node809;
											assign node809 = (inp[15]) ? node825 : node810;
												assign node810 = (inp[0]) ? node818 : node811;
													assign node811 = (inp[2]) ? node815 : node812;
														assign node812 = (inp[12]) ? 40'b0011000000011100000000000010100000000000 : 40'b1011000000010100000000000000100000000000;
														assign node815 = (inp[12]) ? 40'b0011000000010100000000000001100000000000 : 40'b0011000000010100000100000010100000000000;
													assign node818 = (inp[12]) ? node822 : node819;
														assign node819 = (inp[2]) ? 40'b0010000000010100000100000010100000000000 : 40'b1010000000010100000000000000100000000000;
														assign node822 = (inp[2]) ? 40'b0010000000010100000000000001100000000000 : 40'b0010000000011100000000000010100000000000;
												assign node825 = (inp[0]) ? node833 : node826;
													assign node826 = (inp[12]) ? node830 : node827;
														assign node827 = (inp[2]) ? 40'b0011000000000100000100000010100000000000 : 40'b1011000000000100000000000000100000000000;
														assign node830 = (inp[2]) ? 40'b0011000000000100000000000001100000000000 : 40'b0011000000001100000000000010100000000000;
													assign node833 = (inp[12]) ? node837 : node834;
														assign node834 = (inp[2]) ? 40'b0010000000000100000100000010100000000000 : 40'b1010000000000100000000000000100000000000;
														assign node837 = (inp[2]) ? 40'b0010000000000100000000000001100000000000 : 40'b0010000000001100000000000010100000000000;
											assign node840 = (inp[0]) ? node856 : node841;
												assign node841 = (inp[15]) ? node849 : node842;
													assign node842 = (inp[2]) ? node846 : node843;
														assign node843 = (inp[12]) ? 40'b0011000000011000000000000010100000000000 : 40'b1011000000010000000000000010100000000000;
														assign node846 = (inp[12]) ? 40'b0011000000010000000000000001100000000000 : 40'b0011000000010000000100000010100000000000;
													assign node849 = (inp[12]) ? node853 : node850;
														assign node850 = (inp[2]) ? 40'b0011000000000000000100000010100000000000 : 40'b1011000000000000000000000000100000000000;
														assign node853 = (inp[2]) ? 40'b0011000000000000000000000001100000000000 : 40'b0011000000001000000000000010100000000000;
												assign node856 = (inp[15]) ? node864 : node857;
													assign node857 = (inp[2]) ? node861 : node858;
														assign node858 = (inp[12]) ? 40'b0010000000011000000000000010100000000000 : 40'b1010000000010000000000000001100000000000;
														assign node861 = (inp[12]) ? 40'b0010000000010000000000000001100000000000 : 40'b0010000000010000000100000010100000000000;
													assign node864 = (inp[6]) ? node868 : node865;
														assign node865 = (inp[5]) ? 40'b0010000000000000000100000010100000000000 : 40'b1010000000000000000000000000100000000000;
														assign node868 = (inp[5]) ? 40'b0010000000000000000000000001100000000000 : 40'b0010000000001000000000000010100000000000;
										assign node871 = (inp[0]) ? node903 : node872;
											assign node872 = (inp[10]) ? node888 : node873;
												assign node873 = (inp[15]) ? node881 : node874;
													assign node874 = (inp[2]) ? node878 : node875;
														assign node875 = (inp[12]) ? 40'b0011000000011100000000000010000000000000 : 40'b1011000000010100000000000000000000000000;
														assign node878 = (inp[5]) ? 40'b0011000000010100000100000011000000000000 : 40'b0011000000010100000000000001000000000000;
													assign node881 = (inp[2]) ? node885 : node882;
														assign node882 = (inp[12]) ? 40'b0011000000001100000000000010000000000000 : 40'b1011000000000100000000000010000000000000;
														assign node885 = (inp[12]) ? 40'b0011000000000100000000000001000000000000 : 40'b0011000000000100000100000010000000000000;
												assign node888 = (inp[15]) ? node896 : node889;
													assign node889 = (inp[5]) ? node893 : node890;
														assign node890 = (inp[6]) ? 40'b0011000000011000000000000010000000000000 : 40'b1011000000010000000000000000000000000000;
														assign node893 = (inp[6]) ? 40'b0011000000010000000000000001000000000000 : 40'b0011000000010000000100000010000000000000;
													assign node896 = (inp[12]) ? node900 : node897;
														assign node897 = (inp[2]) ? 40'b0011000000000000000100000010000000000000 : 40'b1011000000000000000000000000000000000000;
														assign node900 = (inp[2]) ? 40'b0011000000000000000000000011000000000000 : 40'b0011000000001000000000000010000000000000;
											assign node903 = (inp[10]) ? node919 : node904;
												assign node904 = (inp[15]) ? node912 : node905;
													assign node905 = (inp[5]) ? node909 : node906;
														assign node906 = (inp[6]) ? 40'b0010000000011100000000000010000000000000 : 40'b1010000000010100000000000000000000000000;
														assign node909 = (inp[2]) ? 40'b0010000000010100000100000011000000000000 : 40'b0010000000011100000000000010000000000000;
													assign node912 = (inp[2]) ? node916 : node913;
														assign node913 = (inp[12]) ? 40'b0010000000001100000000000010000000000000 : 40'b1010000000000100000000000010000000000000;
														assign node916 = (inp[5]) ? 40'b0010000000000100000100000011000000000000 : 40'b0010000000000100000100000010000000000000;
												assign node919 = (inp[15]) ? node927 : node920;
													assign node920 = (inp[2]) ? node924 : node921;
														assign node921 = (inp[12]) ? 40'b0010000000011000000000000010000000000000 : 40'b1010000000010000000000000000000000000000;
														assign node924 = (inp[12]) ? 40'b0010000000010000000000000011000000000000 : 40'b0010000000010000000100000010000000000000;
													assign node927 = (inp[5]) ? node931 : node928;
														assign node928 = (inp[6]) ? 40'b0010000000001000000000000010000000000000 : 40'b1010000000000000000000000010000000000000;
														assign node931 = (inp[6]) ? 40'b0010000000000000000000000001000000000000 : 40'b0010000000000000000100000010000000000000;
						assign node934 = (inp[3]) ? node1008 : node935;
							assign node935 = (inp[11]) ? node983 : node936;
								assign node936 = (inp[14]) ? node938 : 40'b0000000000000000000000000000000000000000;
									assign node938 = (inp[15]) ? node952 : node939;
										assign node939 = (inp[13]) ? node941 : 40'b0000000000000000000000000000000000000000;
											assign node941 = (inp[0]) ? node943 : 40'b0000000000000000000000000000000000000000;
												assign node943 = (inp[10]) ? node945 : 40'b0000000000000000000000000000000000000000;
													assign node945 = (inp[6]) ? node949 : node946;
														assign node946 = (inp[12]) ? 40'b0000001100011000000000000010000000000000 : 40'b1000001100010000000100000010000000000000;
														assign node949 = (inp[12]) ? 40'b0000001100011000000000000011000000000000 : 40'b0000001100011000000100000010000000000000;
										assign node952 = (inp[13]) ? node964 : node953;
											assign node953 = (inp[0]) ? node955 : 40'b0000000000000000000000000000000000000000;
												assign node955 = (inp[10]) ? node957 : 40'b0000000000000000000000000000000000000000;
													assign node957 = (inp[12]) ? node961 : node958;
														assign node958 = (inp[2]) ? 40'b0000001100000000000100000010100000000000 : 40'b1000001100000000000000000000100000000000;
														assign node961 = (inp[2]) ? 40'b0000001100000000000000000001100000000000 : 40'b0000001100001000000000000010100000000000;
											assign node964 = (inp[0]) ? node974 : node965;
												assign node965 = (inp[10]) ? node967 : 40'b0000000000000000000000000000000000000000;
													assign node967 = (inp[2]) ? node971 : node968;
														assign node968 = (inp[12]) ? 40'b0001001100001000000000000010000000000000 : 40'b1001001100000000000000000000000000000000;
														assign node971 = (inp[12]) ? 40'b0001001100000000000000000001000000000000 : 40'b0001001100000000000100000010000000000000;
												assign node974 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node975;
													assign node975 = (inp[12]) ? node979 : node976;
														assign node976 = (inp[2]) ? 40'b0000001100000100000100000010000000000000 : 40'b1000001100000100000000000000000000000000;
														assign node979 = (inp[2]) ? 40'b0000001100000100000000000001000000000000 : 40'b0000001100001100000000000010000000000000;
								assign node983 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node984;
									assign node984 = (inp[15]) ? node996 : node985;
										assign node985 = (inp[0]) ? node991 : node986;
											assign node986 = (inp[10]) ? node988 : 40'b0000000000000000000000000000000000000000;
												assign node988 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
											assign node991 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node992;
												assign node992 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
										assign node996 = (inp[0]) ? node1002 : node997;
											assign node997 = (inp[10]) ? node999 : 40'b0000000000000000000000000000000000000000;
												assign node999 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
											assign node1002 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node1003;
												assign node1003 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
							assign node1008 = (inp[11]) ? node1138 : node1009;
								assign node1009 = (inp[14]) ? node1011 : 40'b0000000000000000000000000000000000000000;
									assign node1011 = (inp[15]) ? node1075 : node1012;
										assign node1012 = (inp[13]) ? node1044 : node1013;
											assign node1013 = (inp[10]) ? node1029 : node1014;
												assign node1014 = (inp[0]) ? node1022 : node1015;
													assign node1015 = (inp[12]) ? node1019 : node1016;
														assign node1016 = (inp[2]) ? 40'b0001001000010100000100000010100000000000 : 40'b1001001000010100000000000010100000000000;
														assign node1019 = (inp[2]) ? 40'b0001001000010100000000000001100000000000 : 40'b0001001000011100000000000010100000000000;
													assign node1022 = (inp[6]) ? node1026 : node1023;
														assign node1023 = (inp[5]) ? 40'b0000001000010100000100000010100000000000 : 40'b1000001000010100000000000000100000000000;
														assign node1026 = (inp[5]) ? 40'b0000001000010100000000000011100000000000 : 40'b0000001000011100000000000010100000000000;
												assign node1029 = (inp[0]) ? node1037 : node1030;
													assign node1030 = (inp[2]) ? node1034 : node1031;
														assign node1031 = (inp[12]) ? 40'b0001001000011000000000000010100000000000 : 40'b1001001000010000000000000000100000000000;
														assign node1034 = (inp[12]) ? 40'b0001001000010000000000000001100000000000 : 40'b0001001000010000000100000010100000000000;
													assign node1037 = (inp[12]) ? node1041 : node1038;
														assign node1038 = (inp[2]) ? 40'b0000001000010000000100000010100000000000 : 40'b1000001000010000000000000000100000000000;
														assign node1041 = (inp[2]) ? 40'b0000001000010000000000000001100000000000 : 40'b0000001000011000000000000010100000000000;
											assign node1044 = (inp[10]) ? node1060 : node1045;
												assign node1045 = (inp[0]) ? node1053 : node1046;
													assign node1046 = (inp[12]) ? node1050 : node1047;
														assign node1047 = (inp[2]) ? 40'b0001001000010100000100000010000000000000 : 40'b1001001000010100000000000000000000000000;
														assign node1050 = (inp[2]) ? 40'b0001001000010100000000000001000000000000 : 40'b0001001000011100000000000010000000000000;
													assign node1053 = (inp[6]) ? node1057 : node1054;
														assign node1054 = (inp[5]) ? 40'b0000001000010100000100000010000000000000 : 40'b1000001000010100000000000000000000000000;
														assign node1057 = (inp[5]) ? 40'b0000001000010100000000000001000000000000 : 40'b0000001000011100000000000010000000000000;
												assign node1060 = (inp[0]) ? node1068 : node1061;
													assign node1061 = (inp[5]) ? node1065 : node1062;
														assign node1062 = (inp[6]) ? 40'b0001001000011000000000000010000000000000 : 40'b1001001000010000000000000000000000000000;
														assign node1065 = (inp[6]) ? 40'b0001001000010000000000000001000000000000 : 40'b0001001000010000000100000010000000000000;
													assign node1068 = (inp[2]) ? node1072 : node1069;
														assign node1069 = (inp[12]) ? 40'b0000001000011000000000000010000000000000 : 40'b1000001000010000000000000000000000000000;
														assign node1072 = (inp[12]) ? 40'b0000001000010000000000000001000000000000 : 40'b0000001000010000000100000010000000000000;
										assign node1075 = (inp[13]) ? node1107 : node1076;
											assign node1076 = (inp[0]) ? node1092 : node1077;
												assign node1077 = (inp[10]) ? node1085 : node1078;
													assign node1078 = (inp[12]) ? node1082 : node1079;
														assign node1079 = (inp[2]) ? 40'b0001001000000100000100000010100000000000 : 40'b1001001000000100000000000000100000000000;
														assign node1082 = (inp[2]) ? 40'b0001001000000100000000000001100000000000 : 40'b0001001000001100000000000010100000000000;
													assign node1085 = (inp[5]) ? node1089 : node1086;
														assign node1086 = (inp[6]) ? 40'b0001001000001000000000000010100000000000 : 40'b1001001000000000000000000000100000000000;
														assign node1089 = (inp[6]) ? 40'b0001001000000000000000000001100000000000 : 40'b0001001000000000000100000010100000000000;
												assign node1092 = (inp[10]) ? node1100 : node1093;
													assign node1093 = (inp[2]) ? node1097 : node1094;
														assign node1094 = (inp[12]) ? 40'b0000001000001100000000000010100000000000 : 40'b1000001000000100000000000000100000000000;
														assign node1097 = (inp[12]) ? 40'b0000001000000100000000000001100000000000 : 40'b0000001000000100000100000010100000000000;
													assign node1100 = (inp[5]) ? node1104 : node1101;
														assign node1101 = (inp[6]) ? 40'b0000001000001000000000000010100000000000 : 40'b1000001000000000000000000000100000000000;
														assign node1104 = (inp[6]) ? 40'b0000001000000000000000000011100000000000 : 40'b0000001000000000000100000010100000000000;
											assign node1107 = (inp[10]) ? node1123 : node1108;
												assign node1108 = (inp[0]) ? node1116 : node1109;
													assign node1109 = (inp[2]) ? node1113 : node1110;
														assign node1110 = (inp[12]) ? 40'b0001001000001100000000000010000000000000 : 40'b1001001000000100000000000000000000000000;
														assign node1113 = (inp[12]) ? 40'b0001001000000100000000000001000000000000 : 40'b0001001000000100000100000010000000000000;
													assign node1116 = (inp[2]) ? node1120 : node1117;
														assign node1117 = (inp[5]) ? 40'b0000001000000100000100000010000000000000 : 40'b1000001000001100000000000010000000000000;
														assign node1120 = (inp[12]) ? 40'b0000001000000100000000000001000000000000 : 40'b0000001000000100000100000010000000000000;
												assign node1123 = (inp[0]) ? node1131 : node1124;
													assign node1124 = (inp[12]) ? node1128 : node1125;
														assign node1125 = (inp[2]) ? 40'b0001001000000000000100000010000000000000 : 40'b1001001000000000000000000000000000000000;
														assign node1128 = (inp[2]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000001000000000000010000000000000;
													assign node1131 = (inp[6]) ? node1135 : node1132;
														assign node1132 = (inp[5]) ? 40'b0000001000000000000100000010000000000000 : 40'b1000001000000000000000000000000000000000;
														assign node1135 = (inp[5]) ? 40'b0000001000000000000000000001000000000000 : 40'b0000001000001000000000000010000000000000;
								assign node1138 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node1139;
									assign node1139 = (inp[13]) ? node1203 : node1140;
										assign node1140 = (inp[15]) ? node1172 : node1141;
											assign node1141 = (inp[0]) ? node1157 : node1142;
												assign node1142 = (inp[10]) ? node1150 : node1143;
													assign node1143 = (inp[12]) ? node1147 : node1144;
														assign node1144 = (inp[2]) ? 40'b0001001000010100000100000010100000001000 : 40'b1001001000010100000000000000100000001000;
														assign node1147 = (inp[2]) ? 40'b0001001000010100000000000001100000001000 : 40'b0001001000011100000000000010100000001000;
													assign node1150 = (inp[5]) ? node1154 : node1151;
														assign node1151 = (inp[6]) ? 40'b0001001000011000000000000010100000001000 : 40'b1001001000010000000000000000100000001000;
														assign node1154 = (inp[6]) ? 40'b0001001000010000000000000001100000001000 : 40'b0001001000010000000100000010100000001000;
												assign node1157 = (inp[10]) ? node1165 : node1158;
													assign node1158 = (inp[12]) ? node1162 : node1159;
														assign node1159 = (inp[2]) ? 40'b0000001000010100000100000010100000001000 : 40'b1000001000010100000000000000100000001000;
														assign node1162 = (inp[2]) ? 40'b0000001000010100000000000001100000001000 : 40'b0000001000011100000000000010100000001000;
													assign node1165 = (inp[12]) ? node1169 : node1166;
														assign node1166 = (inp[2]) ? 40'b0000001000010000000100000010100000001000 : 40'b1000001000010000000000000000100000001000;
														assign node1169 = (inp[2]) ? 40'b0000001000010000000000000011100000001000 : 40'b0000001000011000000000000010100000001000;
											assign node1172 = (inp[10]) ? node1188 : node1173;
												assign node1173 = (inp[0]) ? node1181 : node1174;
													assign node1174 = (inp[6]) ? node1178 : node1175;
														assign node1175 = (inp[5]) ? 40'b0001001000000100000100000010100000001000 : 40'b1001001000000100000000000000100000001000;
														assign node1178 = (inp[5]) ? 40'b0001001000000100000000000011100000001000 : 40'b0001001000001100000000000010100000001000;
													assign node1181 = (inp[6]) ? node1185 : node1182;
														assign node1182 = (inp[5]) ? 40'b0000001000000100000100000010100000001000 : 40'b1000001000000100000000000010100000001000;
														assign node1185 = (inp[5]) ? 40'b0000001000000100000000000011100000001000 : 40'b0000001000001100000000000010100000001000;
												assign node1188 = (inp[0]) ? node1196 : node1189;
													assign node1189 = (inp[6]) ? node1193 : node1190;
														assign node1190 = (inp[5]) ? 40'b0001001000000000000100000010100000001000 : 40'b1001001000000000000000000010100000001000;
														assign node1193 = (inp[5]) ? 40'b0001001000000000000000000001100000001000 : 40'b0001001000001000000000000010100000001000;
													assign node1196 = (inp[12]) ? node1200 : node1197;
														assign node1197 = (inp[2]) ? 40'b0000001000000000000100000010100000001000 : 40'b1000001000000000000000000010100000001000;
														assign node1200 = (inp[2]) ? 40'b0000001000000000000000000001100000001000 : 40'b0000001000001000000000000010100000001000;
										assign node1203 = (inp[15]) ? node1235 : node1204;
											assign node1204 = (inp[0]) ? node1220 : node1205;
												assign node1205 = (inp[10]) ? node1213 : node1206;
													assign node1206 = (inp[12]) ? node1210 : node1207;
														assign node1207 = (inp[2]) ? 40'b0001001000010100000100000010000000001000 : 40'b1001001000010100000000000000000000001000;
														assign node1210 = (inp[2]) ? 40'b0001001000010100000000000001000000001000 : 40'b0001001000011100000000000010000000001000;
													assign node1213 = (inp[6]) ? node1217 : node1214;
														assign node1214 = (inp[5]) ? 40'b0001001000010000000100000010000000001000 : 40'b1001001000010000000000000000000000001000;
														assign node1217 = (inp[5]) ? 40'b0001001000010000000000000001000000001000 : 40'b0001001000011000000000000010000000001000;
												assign node1220 = (inp[10]) ? node1228 : node1221;
													assign node1221 = (inp[12]) ? node1225 : node1222;
														assign node1222 = (inp[2]) ? 40'b0000001000010100000100000010000000001000 : 40'b1000001000010100000000000000000000001000;
														assign node1225 = (inp[2]) ? 40'b0000001000010100000000000001000000001000 : 40'b0000001000011100000000000010000000001000;
													assign node1228 = (inp[12]) ? node1232 : node1229;
														assign node1229 = (inp[2]) ? 40'b0000001000010000000100000010000000001000 : 40'b1000001000010000000000000000000000001000;
														assign node1232 = (inp[2]) ? 40'b0000001000010000000000000011000000001000 : 40'b0000001000011000000000000010000000001000;
											assign node1235 = (inp[10]) ? node1251 : node1236;
												assign node1236 = (inp[0]) ? node1244 : node1237;
													assign node1237 = (inp[6]) ? node1241 : node1238;
														assign node1238 = (inp[5]) ? 40'b0001001000000100000100000010000000001000 : 40'b1001001000000100000000000000000000001000;
														assign node1241 = (inp[5]) ? 40'b0001001000000100000000000001000000001000 : 40'b0001001000001100000000000010000000001000;
													assign node1244 = (inp[2]) ? node1248 : node1245;
														assign node1245 = (inp[12]) ? 40'b0000001000001100000000000010000000001000 : 40'b1000001000000100000000000000000000001000;
														assign node1248 = (inp[12]) ? 40'b0000001000000100000000000001000000001000 : 40'b0000001000000100000100000010000000001000;
												assign node1251 = (inp[0]) ? node1259 : node1252;
													assign node1252 = (inp[5]) ? node1256 : node1253;
														assign node1253 = (inp[6]) ? 40'b0001001000001000000000000010000000001000 : 40'b1001001000000000000000000000000000001000;
														assign node1256 = (inp[6]) ? 40'b0001001000000000000000000001000000001000 : 40'b0001001000000000000100000010000000001000;
													assign node1259 = (inp[5]) ? node1263 : node1260;
														assign node1260 = (inp[6]) ? 40'b0000001000001000000000000010000000001000 : 40'b1000001000000000000000000000000000001000;
														assign node1263 = (inp[6]) ? 40'b0000001000000000000000000001000000001000 : 40'b0000001000000000000100000010000000001000;

endmodule