module dtc_split75_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node705;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node711;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node836;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node996;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1072;
	wire [3-1:0] node1074;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1083;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1093;
	wire [3-1:0] node1095;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1143;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1173;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1188;
	wire [3-1:0] node1192;
	wire [3-1:0] node1194;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1216;
	wire [3-1:0] node1219;
	wire [3-1:0] node1221;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1295;
	wire [3-1:0] node1298;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1319;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1350;
	wire [3-1:0] node1352;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1404;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1415;
	wire [3-1:0] node1417;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1424;
	wire [3-1:0] node1427;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1443;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1471;
	wire [3-1:0] node1473;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1487;
	wire [3-1:0] node1488;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1501;
	wire [3-1:0] node1504;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1523;
	wire [3-1:0] node1524;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1541;
	wire [3-1:0] node1543;
	wire [3-1:0] node1546;
	wire [3-1:0] node1548;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1563;
	wire [3-1:0] node1564;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1574;
	wire [3-1:0] node1577;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1581;
	wire [3-1:0] node1584;
	wire [3-1:0] node1585;
	wire [3-1:0] node1589;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1596;
	wire [3-1:0] node1597;
	wire [3-1:0] node1598;
	wire [3-1:0] node1599;
	wire [3-1:0] node1603;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1609;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1615;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1620;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1629;
	wire [3-1:0] node1630;
	wire [3-1:0] node1632;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1638;
	wire [3-1:0] node1641;
	wire [3-1:0] node1644;
	wire [3-1:0] node1646;
	wire [3-1:0] node1648;
	wire [3-1:0] node1650;
	wire [3-1:0] node1653;
	wire [3-1:0] node1654;
	wire [3-1:0] node1655;
	wire [3-1:0] node1657;
	wire [3-1:0] node1660;
	wire [3-1:0] node1661;
	wire [3-1:0] node1663;
	wire [3-1:0] node1667;
	wire [3-1:0] node1668;
	wire [3-1:0] node1669;
	wire [3-1:0] node1671;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1679;
	wire [3-1:0] node1680;
	wire [3-1:0] node1683;
	wire [3-1:0] node1686;
	wire [3-1:0] node1687;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1690;
	wire [3-1:0] node1692;
	wire [3-1:0] node1693;
	wire [3-1:0] node1696;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1703;
	wire [3-1:0] node1704;
	wire [3-1:0] node1707;
	wire [3-1:0] node1710;
	wire [3-1:0] node1712;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1719;
	wire [3-1:0] node1721;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1726;
	wire [3-1:0] node1730;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1740;
	wire [3-1:0] node1743;
	wire [3-1:0] node1744;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1750;
	wire [3-1:0] node1751;
	wire [3-1:0] node1753;
	wire [3-1:0] node1755;
	wire [3-1:0] node1759;
	wire [3-1:0] node1760;
	wire [3-1:0] node1761;
	wire [3-1:0] node1763;
	wire [3-1:0] node1766;
	wire [3-1:0] node1767;
	wire [3-1:0] node1771;
	wire [3-1:0] node1772;
	wire [3-1:0] node1775;
	wire [3-1:0] node1777;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1783;
	wire [3-1:0] node1784;
	wire [3-1:0] node1788;
	wire [3-1:0] node1791;
	wire [3-1:0] node1792;
	wire [3-1:0] node1794;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1802;
	wire [3-1:0] node1803;
	wire [3-1:0] node1805;
	wire [3-1:0] node1808;
	wire [3-1:0] node1810;
	wire [3-1:0] node1812;
	wire [3-1:0] node1815;
	wire [3-1:0] node1816;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1827;
	wire [3-1:0] node1830;
	wire [3-1:0] node1831;
	wire [3-1:0] node1833;
	wire [3-1:0] node1836;
	wire [3-1:0] node1837;
	wire [3-1:0] node1838;
	wire [3-1:0] node1841;
	wire [3-1:0] node1844;
	wire [3-1:0] node1845;
	wire [3-1:0] node1848;
	wire [3-1:0] node1851;
	wire [3-1:0] node1852;
	wire [3-1:0] node1854;
	wire [3-1:0] node1857;
	wire [3-1:0] node1858;
	wire [3-1:0] node1859;
	wire [3-1:0] node1860;
	wire [3-1:0] node1863;
	wire [3-1:0] node1866;
	wire [3-1:0] node1867;
	wire [3-1:0] node1871;
	wire [3-1:0] node1872;
	wire [3-1:0] node1873;
	wire [3-1:0] node1877;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1882;
	wire [3-1:0] node1883;
	wire [3-1:0] node1884;
	wire [3-1:0] node1885;
	wire [3-1:0] node1889;
	wire [3-1:0] node1892;
	wire [3-1:0] node1895;
	wire [3-1:0] node1896;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1903;
	wire [3-1:0] node1906;
	wire [3-1:0] node1907;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1912;
	wire [3-1:0] node1915;
	wire [3-1:0] node1917;
	wire [3-1:0] node1918;
	wire [3-1:0] node1922;
	wire [3-1:0] node1923;
	wire [3-1:0] node1924;
	wire [3-1:0] node1927;
	wire [3-1:0] node1930;
	wire [3-1:0] node1931;
	wire [3-1:0] node1935;
	wire [3-1:0] node1936;
	wire [3-1:0] node1937;
	wire [3-1:0] node1938;
	wire [3-1:0] node1939;
	wire [3-1:0] node1940;
	wire [3-1:0] node1942;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1949;
	wire [3-1:0] node1952;
	wire [3-1:0] node1953;
	wire [3-1:0] node1957;
	wire [3-1:0] node1958;
	wire [3-1:0] node1959;
	wire [3-1:0] node1962;
	wire [3-1:0] node1965;
	wire [3-1:0] node1966;
	wire [3-1:0] node1968;
	wire [3-1:0] node1971;
	wire [3-1:0] node1973;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1978;
	wire [3-1:0] node1980;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1985;
	wire [3-1:0] node1988;
	wire [3-1:0] node1991;
	wire [3-1:0] node1992;
	wire [3-1:0] node1996;
	wire [3-1:0] node1997;
	wire [3-1:0] node1998;
	wire [3-1:0] node1999;
	wire [3-1:0] node2004;
	wire [3-1:0] node2005;
	wire [3-1:0] node2009;
	wire [3-1:0] node2010;
	wire [3-1:0] node2011;
	wire [3-1:0] node2012;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2018;
	wire [3-1:0] node2020;
	wire [3-1:0] node2023;
	wire [3-1:0] node2024;
	wire [3-1:0] node2027;
	wire [3-1:0] node2030;
	wire [3-1:0] node2031;
	wire [3-1:0] node2032;
	wire [3-1:0] node2036;
	wire [3-1:0] node2037;
	wire [3-1:0] node2040;
	wire [3-1:0] node2042;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2047;
	wire [3-1:0] node2049;
	wire [3-1:0] node2051;
	wire [3-1:0] node2054;
	wire [3-1:0] node2055;
	wire [3-1:0] node2058;
	wire [3-1:0] node2060;
	wire [3-1:0] node2063;
	wire [3-1:0] node2064;
	wire [3-1:0] node2065;
	wire [3-1:0] node2068;
	wire [3-1:0] node2069;
	wire [3-1:0] node2073;
	wire [3-1:0] node2076;
	wire [3-1:0] node2077;
	wire [3-1:0] node2078;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2081;
	wire [3-1:0] node2082;
	wire [3-1:0] node2083;
	wire [3-1:0] node2084;
	wire [3-1:0] node2088;
	wire [3-1:0] node2089;
	wire [3-1:0] node2092;
	wire [3-1:0] node2093;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2101;
	wire [3-1:0] node2104;
	wire [3-1:0] node2107;
	wire [3-1:0] node2108;
	wire [3-1:0] node2109;
	wire [3-1:0] node2112;
	wire [3-1:0] node2115;
	wire [3-1:0] node2117;
	wire [3-1:0] node2120;
	wire [3-1:0] node2121;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2125;
	wire [3-1:0] node2130;
	wire [3-1:0] node2131;
	wire [3-1:0] node2132;
	wire [3-1:0] node2135;
	wire [3-1:0] node2136;
	wire [3-1:0] node2140;
	wire [3-1:0] node2142;
	wire [3-1:0] node2145;
	wire [3-1:0] node2146;
	wire [3-1:0] node2147;
	wire [3-1:0] node2149;
	wire [3-1:0] node2150;
	wire [3-1:0] node2154;
	wire [3-1:0] node2155;
	wire [3-1:0] node2158;
	wire [3-1:0] node2160;
	wire [3-1:0] node2163;
	wire [3-1:0] node2164;
	wire [3-1:0] node2165;
	wire [3-1:0] node2167;
	wire [3-1:0] node2169;
	wire [3-1:0] node2172;
	wire [3-1:0] node2174;
	wire [3-1:0] node2175;
	wire [3-1:0] node2178;
	wire [3-1:0] node2181;
	wire [3-1:0] node2182;
	wire [3-1:0] node2183;
	wire [3-1:0] node2187;
	wire [3-1:0] node2188;
	wire [3-1:0] node2191;
	wire [3-1:0] node2194;
	wire [3-1:0] node2195;
	wire [3-1:0] node2196;
	wire [3-1:0] node2197;
	wire [3-1:0] node2200;
	wire [3-1:0] node2201;
	wire [3-1:0] node2202;
	wire [3-1:0] node2204;
	wire [3-1:0] node2208;
	wire [3-1:0] node2209;
	wire [3-1:0] node2211;
	wire [3-1:0] node2215;
	wire [3-1:0] node2216;
	wire [3-1:0] node2217;
	wire [3-1:0] node2218;
	wire [3-1:0] node2221;
	wire [3-1:0] node2224;
	wire [3-1:0] node2225;
	wire [3-1:0] node2228;
	wire [3-1:0] node2231;
	wire [3-1:0] node2232;
	wire [3-1:0] node2233;
	wire [3-1:0] node2235;
	wire [3-1:0] node2238;
	wire [3-1:0] node2240;
	wire [3-1:0] node2243;
	wire [3-1:0] node2245;
	wire [3-1:0] node2248;
	wire [3-1:0] node2249;
	wire [3-1:0] node2250;
	wire [3-1:0] node2251;
	wire [3-1:0] node2252;
	wire [3-1:0] node2253;
	wire [3-1:0] node2258;
	wire [3-1:0] node2259;
	wire [3-1:0] node2261;
	wire [3-1:0] node2265;
	wire [3-1:0] node2266;
	wire [3-1:0] node2267;
	wire [3-1:0] node2269;
	wire [3-1:0] node2272;
	wire [3-1:0] node2275;
	wire [3-1:0] node2277;
	wire [3-1:0] node2280;
	wire [3-1:0] node2281;
	wire [3-1:0] node2282;
	wire [3-1:0] node2283;
	wire [3-1:0] node2287;
	wire [3-1:0] node2288;
	wire [3-1:0] node2290;
	wire [3-1:0] node2293;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2298;
	wire [3-1:0] node2303;
	wire [3-1:0] node2304;
	wire [3-1:0] node2305;
	wire [3-1:0] node2306;
	wire [3-1:0] node2307;
	wire [3-1:0] node2309;
	wire [3-1:0] node2311;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2318;
	wire [3-1:0] node2321;
	wire [3-1:0] node2322;
	wire [3-1:0] node2323;
	wire [3-1:0] node2324;
	wire [3-1:0] node2328;
	wire [3-1:0] node2329;
	wire [3-1:0] node2333;
	wire [3-1:0] node2334;
	wire [3-1:0] node2335;
	wire [3-1:0] node2339;
	wire [3-1:0] node2340;
	wire [3-1:0] node2344;
	wire [3-1:0] node2345;
	wire [3-1:0] node2346;
	wire [3-1:0] node2347;
	wire [3-1:0] node2348;
	wire [3-1:0] node2350;
	wire [3-1:0] node2354;
	wire [3-1:0] node2355;
	wire [3-1:0] node2358;
	wire [3-1:0] node2359;
	wire [3-1:0] node2362;
	wire [3-1:0] node2365;
	wire [3-1:0] node2366;
	wire [3-1:0] node2367;
	wire [3-1:0] node2370;
	wire [3-1:0] node2373;
	wire [3-1:0] node2375;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2380;
	wire [3-1:0] node2383;
	wire [3-1:0] node2385;
	wire [3-1:0] node2386;
	wire [3-1:0] node2390;
	wire [3-1:0] node2391;
	wire [3-1:0] node2393;
	wire [3-1:0] node2394;
	wire [3-1:0] node2398;
	wire [3-1:0] node2399;
	wire [3-1:0] node2402;
	wire [3-1:0] node2403;
	wire [3-1:0] node2407;
	wire [3-1:0] node2408;
	wire [3-1:0] node2409;
	wire [3-1:0] node2410;
	wire [3-1:0] node2411;
	wire [3-1:0] node2412;
	wire [3-1:0] node2415;
	wire [3-1:0] node2418;
	wire [3-1:0] node2421;
	wire [3-1:0] node2422;
	wire [3-1:0] node2423;
	wire [3-1:0] node2424;
	wire [3-1:0] node2429;
	wire [3-1:0] node2432;
	wire [3-1:0] node2433;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2441;
	wire [3-1:0] node2442;
	wire [3-1:0] node2446;
	wire [3-1:0] node2447;
	wire [3-1:0] node2448;
	wire [3-1:0] node2449;
	wire [3-1:0] node2453;
	wire [3-1:0] node2455;
	wire [3-1:0] node2458;
	wire [3-1:0] node2459;
	wire [3-1:0] node2460;
	wire [3-1:0] node2464;
	wire [3-1:0] node2465;
	wire [3-1:0] node2469;
	wire [3-1:0] node2470;
	wire [3-1:0] node2471;
	wire [3-1:0] node2472;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2478;
	wire [3-1:0] node2479;
	wire [3-1:0] node2482;
	wire [3-1:0] node2486;
	wire [3-1:0] node2487;
	wire [3-1:0] node2488;
	wire [3-1:0] node2489;
	wire [3-1:0] node2492;
	wire [3-1:0] node2495;
	wire [3-1:0] node2498;
	wire [3-1:0] node2500;
	wire [3-1:0] node2502;
	wire [3-1:0] node2505;
	wire [3-1:0] node2506;
	wire [3-1:0] node2507;
	wire [3-1:0] node2509;
	wire [3-1:0] node2512;
	wire [3-1:0] node2513;
	wire [3-1:0] node2515;
	wire [3-1:0] node2519;
	wire [3-1:0] node2520;
	wire [3-1:0] node2521;
	wire [3-1:0] node2525;
	wire [3-1:0] node2527;
	wire [3-1:0] node2530;
	wire [3-1:0] node2531;
	wire [3-1:0] node2532;
	wire [3-1:0] node2533;
	wire [3-1:0] node2534;
	wire [3-1:0] node2535;
	wire [3-1:0] node2536;
	wire [3-1:0] node2537;
	wire [3-1:0] node2539;
	wire [3-1:0] node2542;
	wire [3-1:0] node2544;
	wire [3-1:0] node2547;
	wire [3-1:0] node2548;
	wire [3-1:0] node2551;
	wire [3-1:0] node2554;
	wire [3-1:0] node2555;
	wire [3-1:0] node2556;
	wire [3-1:0] node2557;
	wire [3-1:0] node2560;
	wire [3-1:0] node2563;
	wire [3-1:0] node2564;
	wire [3-1:0] node2568;
	wire [3-1:0] node2569;
	wire [3-1:0] node2572;
	wire [3-1:0] node2575;
	wire [3-1:0] node2576;
	wire [3-1:0] node2578;
	wire [3-1:0] node2579;
	wire [3-1:0] node2582;
	wire [3-1:0] node2585;
	wire [3-1:0] node2586;
	wire [3-1:0] node2587;
	wire [3-1:0] node2589;
	wire [3-1:0] node2592;
	wire [3-1:0] node2595;
	wire [3-1:0] node2596;
	wire [3-1:0] node2599;
	wire [3-1:0] node2602;
	wire [3-1:0] node2603;
	wire [3-1:0] node2604;
	wire [3-1:0] node2605;
	wire [3-1:0] node2606;
	wire [3-1:0] node2610;
	wire [3-1:0] node2611;
	wire [3-1:0] node2614;
	wire [3-1:0] node2617;
	wire [3-1:0] node2619;
	wire [3-1:0] node2621;
	wire [3-1:0] node2624;
	wire [3-1:0] node2625;
	wire [3-1:0] node2626;
	wire [3-1:0] node2628;
	wire [3-1:0] node2629;
	wire [3-1:0] node2633;
	wire [3-1:0] node2635;
	wire [3-1:0] node2638;
	wire [3-1:0] node2639;
	wire [3-1:0] node2641;
	wire [3-1:0] node2644;
	wire [3-1:0] node2646;
	wire [3-1:0] node2649;
	wire [3-1:0] node2650;
	wire [3-1:0] node2651;
	wire [3-1:0] node2652;
	wire [3-1:0] node2653;
	wire [3-1:0] node2654;
	wire [3-1:0] node2656;
	wire [3-1:0] node2659;
	wire [3-1:0] node2662;
	wire [3-1:0] node2663;
	wire [3-1:0] node2666;
	wire [3-1:0] node2668;
	wire [3-1:0] node2671;
	wire [3-1:0] node2672;
	wire [3-1:0] node2673;
	wire [3-1:0] node2674;
	wire [3-1:0] node2678;
	wire [3-1:0] node2681;
	wire [3-1:0] node2682;
	wire [3-1:0] node2685;
	wire [3-1:0] node2688;
	wire [3-1:0] node2689;
	wire [3-1:0] node2690;
	wire [3-1:0] node2691;
	wire [3-1:0] node2695;
	wire [3-1:0] node2696;
	wire [3-1:0] node2699;
	wire [3-1:0] node2702;
	wire [3-1:0] node2704;
	wire [3-1:0] node2705;
	wire [3-1:0] node2706;
	wire [3-1:0] node2709;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2717;
	wire [3-1:0] node2718;
	wire [3-1:0] node2719;
	wire [3-1:0] node2720;
	wire [3-1:0] node2721;
	wire [3-1:0] node2725;
	wire [3-1:0] node2726;
	wire [3-1:0] node2728;
	wire [3-1:0] node2731;
	wire [3-1:0] node2734;
	wire [3-1:0] node2735;
	wire [3-1:0] node2736;
	wire [3-1:0] node2738;
	wire [3-1:0] node2742;
	wire [3-1:0] node2743;
	wire [3-1:0] node2745;
	wire [3-1:0] node2748;
	wire [3-1:0] node2749;
	wire [3-1:0] node2753;
	wire [3-1:0] node2754;
	wire [3-1:0] node2755;
	wire [3-1:0] node2756;
	wire [3-1:0] node2759;
	wire [3-1:0] node2761;
	wire [3-1:0] node2764;
	wire [3-1:0] node2765;
	wire [3-1:0] node2768;
	wire [3-1:0] node2771;
	wire [3-1:0] node2772;
	wire [3-1:0] node2774;
	wire [3-1:0] node2776;
	wire [3-1:0] node2779;
	wire [3-1:0] node2780;
	wire [3-1:0] node2781;
	wire [3-1:0] node2785;
	wire [3-1:0] node2788;
	wire [3-1:0] node2789;
	wire [3-1:0] node2790;
	wire [3-1:0] node2791;
	wire [3-1:0] node2792;
	wire [3-1:0] node2793;
	wire [3-1:0] node2794;
	wire [3-1:0] node2797;
	wire [3-1:0] node2800;
	wire [3-1:0] node2801;
	wire [3-1:0] node2802;
	wire [3-1:0] node2806;
	wire [3-1:0] node2807;
	wire [3-1:0] node2811;
	wire [3-1:0] node2812;
	wire [3-1:0] node2814;
	wire [3-1:0] node2817;
	wire [3-1:0] node2819;
	wire [3-1:0] node2822;
	wire [3-1:0] node2823;
	wire [3-1:0] node2824;
	wire [3-1:0] node2826;
	wire [3-1:0] node2829;
	wire [3-1:0] node2830;
	wire [3-1:0] node2835;
	wire [3-1:0] node2836;
	wire [3-1:0] node2837;
	wire [3-1:0] node2838;
	wire [3-1:0] node2839;
	wire [3-1:0] node2840;
	wire [3-1:0] node2845;
	wire [3-1:0] node2846;
	wire [3-1:0] node2848;
	wire [3-1:0] node2851;
	wire [3-1:0] node2854;
	wire [3-1:0] node2855;
	wire [3-1:0] node2856;
	wire [3-1:0] node2858;
	wire [3-1:0] node2861;
	wire [3-1:0] node2862;
	wire [3-1:0] node2866;
	wire [3-1:0] node2867;
	wire [3-1:0] node2870;
	wire [3-1:0] node2871;
	wire [3-1:0] node2875;
	wire [3-1:0] node2876;
	wire [3-1:0] node2877;
	wire [3-1:0] node2879;
	wire [3-1:0] node2881;
	wire [3-1:0] node2884;
	wire [3-1:0] node2887;
	wire [3-1:0] node2888;
	wire [3-1:0] node2891;
	wire [3-1:0] node2892;
	wire [3-1:0] node2896;
	wire [3-1:0] node2898;
	wire [3-1:0] node2899;
	wire [3-1:0] node2900;
	wire [3-1:0] node2901;
	wire [3-1:0] node2903;
	wire [3-1:0] node2906;
	wire [3-1:0] node2907;
	wire [3-1:0] node2910;
	wire [3-1:0] node2913;
	wire [3-1:0] node2914;
	wire [3-1:0] node2915;
	wire [3-1:0] node2919;
	wire [3-1:0] node2921;
	wire [3-1:0] node2924;
	wire [3-1:0] node2925;
	wire [3-1:0] node2926;
	wire [3-1:0] node2927;
	wire [3-1:0] node2931;
	wire [3-1:0] node2932;

	assign outp = (inp[6]) ? node1200 : node1;
		assign node1 = (inp[3]) ? node919 : node2;
			assign node2 = (inp[9]) ? node540 : node3;
				assign node3 = (inp[0]) ? node267 : node4;
					assign node4 = (inp[4]) ? node122 : node5;
						assign node5 = (inp[1]) ? node63 : node6;
							assign node6 = (inp[7]) ? node44 : node7;
								assign node7 = (inp[10]) ? node27 : node8;
									assign node8 = (inp[11]) ? node20 : node9;
										assign node9 = (inp[2]) ? node17 : node10;
											assign node10 = (inp[5]) ? node14 : node11;
												assign node11 = (inp[8]) ? 3'b111 : 3'b011;
												assign node14 = (inp[8]) ? 3'b011 : 3'b111;
											assign node17 = (inp[5]) ? 3'b001 : 3'b011;
										assign node20 = (inp[5]) ? 3'b101 : node21;
											assign node21 = (inp[8]) ? 3'b011 : node22;
												assign node22 = (inp[2]) ? 3'b101 : 3'b001;
									assign node27 = (inp[2]) ? node37 : node28;
										assign node28 = (inp[8]) ? node32 : node29;
											assign node29 = (inp[5]) ? 3'b001 : 3'b101;
											assign node32 = (inp[11]) ? 3'b001 : node33;
												assign node33 = (inp[5]) ? 3'b101 : 3'b001;
										assign node37 = (inp[11]) ? node41 : node38;
											assign node38 = (inp[5]) ? 3'b001 : 3'b101;
											assign node41 = (inp[5]) ? 3'b110 : 3'b001;
								assign node44 = (inp[2]) ? node56 : node45;
									assign node45 = (inp[5]) ? node51 : node46;
										assign node46 = (inp[10]) ? 3'b001 : node47;
											assign node47 = (inp[8]) ? 3'b000 : 3'b001;
										assign node51 = (inp[10]) ? node53 : 3'b001;
											assign node53 = (inp[8]) ? 3'b001 : 3'b000;
									assign node56 = (inp[8]) ? 3'b001 : node57;
										assign node57 = (inp[5]) ? node59 : 3'b001;
											assign node59 = (inp[10]) ? 3'b000 : 3'b001;
							assign node63 = (inp[7]) ? node87 : node64;
								assign node64 = (inp[10]) ? node80 : node65;
									assign node65 = (inp[11]) ? node73 : node66;
										assign node66 = (inp[8]) ? node68 : 3'b001;
											assign node68 = (inp[5]) ? node70 : 3'b011;
												assign node70 = (inp[2]) ? 3'b001 : 3'b101;
										assign node73 = (inp[8]) ? node77 : node74;
											assign node74 = (inp[5]) ? 3'b110 : 3'b101;
											assign node77 = (inp[5]) ? 3'b001 : 3'b101;
									assign node80 = (inp[8]) ? node82 : 3'b110;
										assign node82 = (inp[2]) ? 3'b110 : node83;
											assign node83 = (inp[5]) ? 3'b001 : 3'b101;
								assign node87 = (inp[10]) ? node107 : node88;
									assign node88 = (inp[8]) ? node96 : node89;
										assign node89 = (inp[5]) ? 3'b101 : node90;
											assign node90 = (inp[11]) ? 3'b101 : node91;
												assign node91 = (inp[2]) ? 3'b011 : 3'b111;
										assign node96 = (inp[5]) ? node102 : node97;
											assign node97 = (inp[2]) ? node99 : 3'b111;
												assign node99 = (inp[11]) ? 3'b011 : 3'b111;
											assign node102 = (inp[2]) ? node104 : 3'b011;
												assign node104 = (inp[11]) ? 3'b101 : 3'b011;
									assign node107 = (inp[11]) ? node113 : node108;
										assign node108 = (inp[8]) ? node110 : 3'b101;
											assign node110 = (inp[5]) ? 3'b101 : 3'b011;
										assign node113 = (inp[8]) ? node115 : 3'b001;
											assign node115 = (inp[5]) ? node119 : node116;
												assign node116 = (inp[2]) ? 3'b101 : 3'b001;
												assign node119 = (inp[2]) ? 3'b001 : 3'b101;
						assign node122 = (inp[7]) ? node206 : node123;
							assign node123 = (inp[11]) ? node165 : node124;
								assign node124 = (inp[1]) ? node146 : node125;
									assign node125 = (inp[8]) ? node139 : node126;
										assign node126 = (inp[2]) ? node134 : node127;
											assign node127 = (inp[10]) ? node131 : node128;
												assign node128 = (inp[5]) ? 3'b110 : 3'b100;
												assign node131 = (inp[5]) ? 3'b100 : 3'b110;
											assign node134 = (inp[10]) ? node136 : 3'b000;
												assign node136 = (inp[5]) ? 3'b000 : 3'b110;
										assign node139 = (inp[10]) ? node143 : node140;
											assign node140 = (inp[5]) ? 3'b000 : 3'b100;
											assign node143 = (inp[5]) ? 3'b110 : 3'b000;
									assign node146 = (inp[8]) ? node156 : node147;
										assign node147 = (inp[5]) ? node153 : node148;
											assign node148 = (inp[2]) ? node150 : 3'b010;
												assign node150 = (inp[10]) ? 3'b010 : 3'b110;
											assign node153 = (inp[2]) ? 3'b100 : 3'b000;
										assign node156 = (inp[2]) ? node158 : 3'b110;
											assign node158 = (inp[10]) ? node162 : node159;
												assign node159 = (inp[5]) ? 3'b110 : 3'b001;
												assign node162 = (inp[5]) ? 3'b010 : 3'b110;
								assign node165 = (inp[2]) ? node187 : node166;
									assign node166 = (inp[10]) ? node178 : node167;
										assign node167 = (inp[8]) ? node171 : node168;
											assign node168 = (inp[1]) ? 3'b110 : 3'b010;
											assign node171 = (inp[1]) ? node175 : node172;
												assign node172 = (inp[5]) ? 3'b000 : 3'b100;
												assign node175 = (inp[5]) ? 3'b110 : 3'b000;
										assign node178 = (inp[1]) ? node180 : 3'b110;
											assign node180 = (inp[8]) ? node184 : node181;
												assign node181 = (inp[5]) ? 3'b100 : 3'b010;
												assign node184 = (inp[5]) ? 3'b010 : 3'b110;
									assign node187 = (inp[1]) ? node199 : node188;
										assign node188 = (inp[10]) ? node194 : node189;
											assign node189 = (inp[8]) ? 3'b010 : node190;
												assign node190 = (inp[5]) ? 3'b110 : 3'b010;
											assign node194 = (inp[5]) ? node196 : 3'b110;
												assign node196 = (inp[8]) ? 3'b110 : 3'b010;
										assign node199 = (inp[8]) ? 3'b010 : node200;
											assign node200 = (inp[5]) ? 3'b100 : node201;
												assign node201 = (inp[10]) ? 3'b010 : 3'b110;
							assign node206 = (inp[1]) ? node244 : node207;
								assign node207 = (inp[10]) ? node223 : node208;
									assign node208 = (inp[11]) ? node216 : node209;
										assign node209 = (inp[2]) ? 3'b101 : node210;
											assign node210 = (inp[8]) ? node212 : 3'b111;
												assign node212 = (inp[5]) ? 3'b011 : 3'b111;
										assign node216 = (inp[8]) ? node220 : node217;
											assign node217 = (inp[2]) ? 3'b101 : 3'b001;
											assign node220 = (inp[5]) ? 3'b101 : 3'b011;
									assign node223 = (inp[2]) ? node231 : node224;
										assign node224 = (inp[11]) ? 3'b001 : node225;
											assign node225 = (inp[5]) ? node227 : 3'b001;
												assign node227 = (inp[8]) ? 3'b101 : 3'b001;
										assign node231 = (inp[11]) ? node237 : node232;
											assign node232 = (inp[8]) ? node234 : 3'b001;
												assign node234 = (inp[5]) ? 3'b001 : 3'b101;
											assign node237 = (inp[5]) ? node241 : node238;
												assign node238 = (inp[8]) ? 3'b101 : 3'b001;
												assign node241 = (inp[8]) ? 3'b000 : 3'b110;
								assign node244 = (inp[10]) ? node258 : node245;
									assign node245 = (inp[11]) ? node251 : node246;
										assign node246 = (inp[8]) ? node248 : 3'b001;
											assign node248 = (inp[5]) ? 3'b001 : 3'b101;
										assign node251 = (inp[5]) ? node255 : node252;
											assign node252 = (inp[2]) ? 3'b001 : 3'b101;
											assign node255 = (inp[8]) ? 3'b001 : 3'b110;
									assign node258 = (inp[5]) ? node262 : node259;
										assign node259 = (inp[8]) ? 3'b001 : 3'b110;
										assign node262 = (inp[8]) ? 3'b110 : node263;
											assign node263 = (inp[2]) ? 3'b010 : 3'b110;
					assign node267 = (inp[4]) ? node403 : node268;
						assign node268 = (inp[7]) ? node342 : node269;
							assign node269 = (inp[10]) ? node305 : node270;
								assign node270 = (inp[1]) ? node294 : node271;
									assign node271 = (inp[8]) ? node281 : node272;
										assign node272 = (inp[2]) ? node276 : node273;
											assign node273 = (inp[5]) ? 3'b110 : 3'b001;
											assign node276 = (inp[11]) ? node278 : 3'b110;
												assign node278 = (inp[5]) ? 3'b010 : 3'b110;
										assign node281 = (inp[11]) ? node287 : node282;
											assign node282 = (inp[5]) ? 3'b001 : node283;
												assign node283 = (inp[2]) ? 3'b001 : 3'b101;
											assign node287 = (inp[5]) ? node291 : node288;
												assign node288 = (inp[2]) ? 3'b001 : 3'b000;
												assign node291 = (inp[2]) ? 3'b110 : 3'b010;
									assign node294 = (inp[5]) ? 3'b010 : node295;
										assign node295 = (inp[2]) ? node299 : node296;
											assign node296 = (inp[11]) ? 3'b110 : 3'b001;
											assign node299 = (inp[8]) ? 3'b110 : node300;
												assign node300 = (inp[11]) ? 3'b010 : 3'b110;
								assign node305 = (inp[5]) ? node327 : node306;
									assign node306 = (inp[8]) ? node316 : node307;
										assign node307 = (inp[1]) ? node313 : node308;
											assign node308 = (inp[11]) ? node310 : 3'b110;
												assign node310 = (inp[2]) ? 3'b010 : 3'b110;
											assign node313 = (inp[11]) ? 3'b110 : 3'b010;
										assign node316 = (inp[11]) ? node322 : node317;
											assign node317 = (inp[1]) ? node319 : 3'b010;
												assign node319 = (inp[2]) ? 3'b010 : 3'b110;
											assign node322 = (inp[2]) ? node324 : 3'b010;
												assign node324 = (inp[1]) ? 3'b010 : 3'b110;
									assign node327 = (inp[8]) ? node335 : node328;
										assign node328 = (inp[1]) ? 3'b100 : node329;
											assign node329 = (inp[11]) ? node331 : 3'b010;
												assign node331 = (inp[2]) ? 3'b100 : 3'b000;
										assign node335 = (inp[1]) ? node339 : node336;
											assign node336 = (inp[11]) ? 3'b010 : 3'b110;
											assign node339 = (inp[11]) ? 3'b100 : 3'b010;
							assign node342 = (inp[1]) ? node380 : node343;
								assign node343 = (inp[2]) ? node365 : node344;
									assign node344 = (inp[11]) ? node356 : node345;
										assign node345 = (inp[8]) ? node349 : node346;
											assign node346 = (inp[5]) ? 3'b010 : 3'b001;
											assign node349 = (inp[5]) ? node353 : node350;
												assign node350 = (inp[10]) ? 3'b101 : 3'b010;
												assign node353 = (inp[10]) ? 3'b001 : 3'b101;
										assign node356 = (inp[10]) ? node362 : node357;
											assign node357 = (inp[8]) ? 3'b010 : node358;
												assign node358 = (inp[5]) ? 3'b001 : 3'b101;
											assign node362 = (inp[5]) ? 3'b110 : 3'b101;
									assign node365 = (inp[5]) ? node375 : node366;
										assign node366 = (inp[10]) ? node372 : node367;
											assign node367 = (inp[11]) ? 3'b101 : node368;
												assign node368 = (inp[8]) ? 3'b011 : 3'b101;
											assign node372 = (inp[8]) ? 3'b101 : 3'b001;
										assign node375 = (inp[11]) ? node377 : 3'b001;
											assign node377 = (inp[8]) ? 3'b001 : 3'b110;
								assign node380 = (inp[10]) ? node392 : node381;
									assign node381 = (inp[5]) ? node389 : node382;
										assign node382 = (inp[8]) ? 3'b101 : node383;
											assign node383 = (inp[2]) ? 3'b001 : node384;
												assign node384 = (inp[11]) ? 3'b001 : 3'b101;
										assign node389 = (inp[8]) ? 3'b001 : 3'b110;
									assign node392 = (inp[8]) ? node396 : node393;
										assign node393 = (inp[5]) ? 3'b010 : 3'b110;
										assign node396 = (inp[5]) ? 3'b110 : node397;
											assign node397 = (inp[11]) ? node399 : 3'b001;
												assign node399 = (inp[2]) ? 3'b110 : 3'b010;
						assign node403 = (inp[7]) ? node465 : node404;
							assign node404 = (inp[10]) ? node430 : node405;
								assign node405 = (inp[1]) ? node413 : node406;
									assign node406 = (inp[5]) ? node410 : node407;
										assign node407 = (inp[11]) ? 3'b010 : 3'b110;
										assign node410 = (inp[8]) ? 3'b010 : 3'b100;
									assign node413 = (inp[5]) ? node421 : node414;
										assign node414 = (inp[2]) ? node416 : 3'b100;
											assign node416 = (inp[11]) ? 3'b100 : node417;
												assign node417 = (inp[8]) ? 3'b010 : 3'b100;
										assign node421 = (inp[11]) ? node427 : node422;
											assign node422 = (inp[8]) ? node424 : 3'b100;
												assign node424 = (inp[2]) ? 3'b100 : 3'b000;
											assign node427 = (inp[8]) ? 3'b100 : 3'b000;
								assign node430 = (inp[1]) ? node454 : node431;
									assign node431 = (inp[11]) ? node441 : node432;
										assign node432 = (inp[8]) ? node438 : node433;
											assign node433 = (inp[5]) ? node435 : 3'b100;
												assign node435 = (inp[2]) ? 3'b000 : 3'b100;
											assign node438 = (inp[5]) ? 3'b100 : 3'b010;
										assign node441 = (inp[2]) ? node449 : node442;
											assign node442 = (inp[8]) ? node446 : node443;
												assign node443 = (inp[5]) ? 3'b000 : 3'b100;
												assign node446 = (inp[5]) ? 3'b100 : 3'b000;
											assign node449 = (inp[8]) ? 3'b100 : node450;
												assign node450 = (inp[5]) ? 3'b000 : 3'b100;
									assign node454 = (inp[11]) ? 3'b000 : node455;
										assign node455 = (inp[8]) ? node457 : 3'b000;
											assign node457 = (inp[2]) ? node461 : node458;
												assign node458 = (inp[5]) ? 3'b100 : 3'b000;
												assign node461 = (inp[5]) ? 3'b000 : 3'b100;
							assign node465 = (inp[10]) ? node507 : node466;
								assign node466 = (inp[5]) ? node484 : node467;
									assign node467 = (inp[1]) ? node479 : node468;
										assign node468 = (inp[11]) ? node472 : node469;
											assign node469 = (inp[8]) ? 3'b101 : 3'b001;
											assign node472 = (inp[8]) ? node476 : node473;
												assign node473 = (inp[2]) ? 3'b110 : 3'b010;
												assign node476 = (inp[2]) ? 3'b001 : 3'b000;
										assign node479 = (inp[8]) ? 3'b110 : node480;
											assign node480 = (inp[11]) ? 3'b100 : 3'b111;
									assign node484 = (inp[2]) ? node492 : node485;
										assign node485 = (inp[11]) ? 3'b010 : node486;
											assign node486 = (inp[8]) ? 3'b110 : node487;
												assign node487 = (inp[1]) ? 3'b010 : 3'b110;
										assign node492 = (inp[8]) ? node500 : node493;
											assign node493 = (inp[11]) ? node497 : node494;
												assign node494 = (inp[1]) ? 3'b010 : 3'b110;
												assign node497 = (inp[1]) ? 3'b100 : 3'b010;
											assign node500 = (inp[1]) ? node504 : node501;
												assign node501 = (inp[11]) ? 3'b110 : 3'b001;
												assign node504 = (inp[11]) ? 3'b010 : 3'b110;
								assign node507 = (inp[5]) ? node527 : node508;
									assign node508 = (inp[1]) ? node518 : node509;
										assign node509 = (inp[11]) ? node511 : 3'b110;
											assign node511 = (inp[8]) ? node515 : node512;
												assign node512 = (inp[2]) ? 3'b010 : 3'b110;
												assign node515 = (inp[2]) ? 3'b110 : 3'b010;
										assign node518 = (inp[11]) ? node520 : 3'b010;
											assign node520 = (inp[8]) ? node524 : node521;
												assign node521 = (inp[2]) ? 3'b100 : 3'b010;
												assign node524 = (inp[2]) ? 3'b010 : 3'b110;
									assign node527 = (inp[11]) ? node535 : node528;
										assign node528 = (inp[1]) ? node532 : node529;
											assign node529 = (inp[8]) ? 3'b110 : 3'b010;
											assign node532 = (inp[8]) ? 3'b010 : 3'b100;
										assign node535 = (inp[2]) ? 3'b100 : node536;
											assign node536 = (inp[1]) ? 3'b100 : 3'b000;
				assign node540 = (inp[4]) ? node764 : node541;
					assign node541 = (inp[7]) ? node651 : node542;
						assign node542 = (inp[0]) ? node602 : node543;
							assign node543 = (inp[1]) ? node577 : node544;
								assign node544 = (inp[10]) ? node558 : node545;
									assign node545 = (inp[5]) ? node553 : node546;
										assign node546 = (inp[2]) ? node548 : 3'b000;
											assign node548 = (inp[8]) ? 3'b010 : node549;
												assign node549 = (inp[11]) ? 3'b100 : 3'b010;
										assign node553 = (inp[8]) ? node555 : 3'b100;
											assign node555 = (inp[2]) ? 3'b100 : 3'b010;
									assign node558 = (inp[11]) ? node566 : node559;
										assign node559 = (inp[8]) ? node563 : node560;
											assign node560 = (inp[5]) ? 3'b000 : 3'b100;
											assign node563 = (inp[5]) ? 3'b100 : 3'b000;
										assign node566 = (inp[2]) ? node572 : node567;
											assign node567 = (inp[8]) ? 3'b100 : node568;
												assign node568 = (inp[5]) ? 3'b000 : 3'b100;
											assign node572 = (inp[8]) ? node574 : 3'b000;
												assign node574 = (inp[5]) ? 3'b000 : 3'b100;
								assign node577 = (inp[10]) ? node591 : node578;
									assign node578 = (inp[5]) ? node586 : node579;
										assign node579 = (inp[11]) ? 3'b110 : node580;
											assign node580 = (inp[2]) ? 3'b110 : node581;
												assign node581 = (inp[8]) ? 3'b111 : 3'b011;
										assign node586 = (inp[11]) ? node588 : 3'b010;
											assign node588 = (inp[8]) ? 3'b010 : 3'b100;
									assign node591 = (inp[5]) ? node597 : node592;
										assign node592 = (inp[8]) ? 3'b010 : node593;
											assign node593 = (inp[11]) ? 3'b100 : 3'b010;
										assign node597 = (inp[11]) ? 3'b100 : node598;
											assign node598 = (inp[2]) ? 3'b100 : 3'b110;
							assign node602 = (inp[11]) ? node624 : node603;
								assign node603 = (inp[10]) ? node615 : node604;
									assign node604 = (inp[1]) ? node610 : node605;
										assign node605 = (inp[8]) ? 3'b010 : node606;
											assign node606 = (inp[5]) ? 3'b100 : 3'b010;
										assign node610 = (inp[5]) ? node612 : 3'b100;
											assign node612 = (inp[8]) ? 3'b100 : 3'b000;
									assign node615 = (inp[1]) ? 3'b000 : node616;
										assign node616 = (inp[8]) ? node620 : node617;
											assign node617 = (inp[5]) ? 3'b000 : 3'b100;
											assign node620 = (inp[5]) ? 3'b100 : 3'b000;
								assign node624 = (inp[1]) ? node644 : node625;
									assign node625 = (inp[8]) ? node635 : node626;
										assign node626 = (inp[2]) ? 3'b000 : node627;
											assign node627 = (inp[10]) ? node631 : node628;
												assign node628 = (inp[5]) ? 3'b100 : 3'b000;
												assign node631 = (inp[5]) ? 3'b000 : 3'b100;
										assign node635 = (inp[5]) ? node639 : node636;
											assign node636 = (inp[10]) ? 3'b100 : 3'b010;
											assign node639 = (inp[2]) ? node641 : 3'b000;
												assign node641 = (inp[10]) ? 3'b000 : 3'b100;
									assign node644 = (inp[8]) ? node646 : 3'b000;
										assign node646 = (inp[2]) ? node648 : 3'b000;
											assign node648 = (inp[5]) ? 3'b000 : 3'b100;
						assign node651 = (inp[0]) ? node715 : node652;
							assign node652 = (inp[1]) ? node678 : node653;
								assign node653 = (inp[8]) ? node667 : node654;
									assign node654 = (inp[10]) ? node660 : node655;
										assign node655 = (inp[11]) ? 3'b000 : node656;
											assign node656 = (inp[5]) ? 3'b000 : 3'b001;
										assign node660 = (inp[11]) ? 3'b100 : node661;
											assign node661 = (inp[5]) ? node663 : 3'b000;
												assign node663 = (inp[2]) ? 3'b100 : 3'b000;
									assign node667 = (inp[10]) ? node675 : node668;
										assign node668 = (inp[5]) ? 3'b101 : node669;
											assign node669 = (inp[2]) ? 3'b101 : node670;
												assign node670 = (inp[11]) ? 3'b100 : 3'b000;
										assign node675 = (inp[2]) ? 3'b000 : 3'b001;
								assign node678 = (inp[11]) ? node698 : node679;
									assign node679 = (inp[8]) ? node693 : node680;
										assign node680 = (inp[2]) ? node688 : node681;
											assign node681 = (inp[5]) ? node685 : node682;
												assign node682 = (inp[10]) ? 3'b110 : 3'b101;
												assign node685 = (inp[10]) ? 3'b101 : 3'b110;
											assign node688 = (inp[10]) ? node690 : 3'b110;
												assign node690 = (inp[5]) ? 3'b001 : 3'b110;
										assign node693 = (inp[10]) ? node695 : 3'b001;
											assign node695 = (inp[5]) ? 3'b110 : 3'b001;
									assign node698 = (inp[8]) ? node708 : node699;
										assign node699 = (inp[2]) ? node705 : node700;
											assign node700 = (inp[10]) ? 3'b110 : node701;
												assign node701 = (inp[5]) ? 3'b110 : 3'b010;
											assign node705 = (inp[10]) ? 3'b010 : 3'b110;
										assign node708 = (inp[2]) ? 3'b110 : node709;
											assign node709 = (inp[10]) ? node711 : 3'b001;
												assign node711 = (inp[5]) ? 3'b110 : 3'b001;
							assign node715 = (inp[10]) ? node737 : node716;
								assign node716 = (inp[2]) ? node730 : node717;
									assign node717 = (inp[1]) ? node721 : node718;
										assign node718 = (inp[8]) ? 3'b110 : 3'b010;
										assign node721 = (inp[5]) ? node727 : node722;
											assign node722 = (inp[8]) ? 3'b110 : node723;
												assign node723 = (inp[11]) ? 3'b010 : 3'b110;
											assign node727 = (inp[8]) ? 3'b010 : 3'b100;
									assign node730 = (inp[1]) ? 3'b010 : node731;
										assign node731 = (inp[8]) ? node733 : 3'b010;
											assign node733 = (inp[5]) ? 3'b110 : 3'b010;
								assign node737 = (inp[1]) ? node753 : node738;
									assign node738 = (inp[5]) ? node746 : node739;
										assign node739 = (inp[8]) ? node741 : 3'b010;
											assign node741 = (inp[2]) ? node743 : 3'b110;
												assign node743 = (inp[11]) ? 3'b010 : 3'b110;
										assign node746 = (inp[8]) ? 3'b010 : node747;
											assign node747 = (inp[2]) ? 3'b100 : node748;
												assign node748 = (inp[11]) ? 3'b100 : 3'b000;
									assign node753 = (inp[5]) ? node761 : node754;
										assign node754 = (inp[8]) ? node756 : 3'b100;
											assign node756 = (inp[2]) ? 3'b100 : node757;
												assign node757 = (inp[11]) ? 3'b000 : 3'b010;
										assign node761 = (inp[8]) ? 3'b100 : 3'b000;
					assign node764 = (inp[0]) ? node860 : node765;
						assign node765 = (inp[10]) ? node819 : node766;
							assign node766 = (inp[1]) ? node782 : node767;
								assign node767 = (inp[7]) ? node769 : 3'b010;
									assign node769 = (inp[5]) ? node775 : node770;
										assign node770 = (inp[2]) ? 3'b010 : node771;
											assign node771 = (inp[11]) ? 3'b000 : 3'b110;
										assign node775 = (inp[8]) ? node779 : node776;
											assign node776 = (inp[11]) ? 3'b000 : 3'b100;
											assign node779 = (inp[11]) ? 3'b100 : 3'b010;
								assign node782 = (inp[7]) ? node800 : node783;
									assign node783 = (inp[2]) ? node791 : node784;
										assign node784 = (inp[8]) ? node788 : node785;
											assign node785 = (inp[5]) ? 3'b000 : 3'b100;
											assign node788 = (inp[5]) ? 3'b100 : 3'b000;
										assign node791 = (inp[5]) ? node797 : node792;
											assign node792 = (inp[8]) ? node794 : 3'b100;
												assign node794 = (inp[11]) ? 3'b000 : 3'b010;
											assign node797 = (inp[8]) ? 3'b100 : 3'b000;
									assign node800 = (inp[11]) ? node812 : node801;
										assign node801 = (inp[5]) ? node807 : node802;
											assign node802 = (inp[2]) ? 3'b010 : node803;
												assign node803 = (inp[8]) ? 3'b001 : 3'b011;
											assign node807 = (inp[8]) ? node809 : 3'b010;
												assign node809 = (inp[2]) ? 3'b010 : 3'b110;
										assign node812 = (inp[5]) ? node816 : node813;
											assign node813 = (inp[8]) ? 3'b110 : 3'b010;
											assign node816 = (inp[8]) ? 3'b010 : 3'b100;
							assign node819 = (inp[7]) ? node829 : node820;
								assign node820 = (inp[1]) ? node824 : node821;
									assign node821 = (inp[5]) ? 3'b000 : 3'b010;
									assign node824 = (inp[8]) ? node826 : 3'b000;
										assign node826 = (inp[5]) ? 3'b000 : 3'b100;
								assign node829 = (inp[1]) ? node841 : node830;
									assign node830 = (inp[5]) ? node836 : node831;
										assign node831 = (inp[8]) ? 3'b100 : node832;
											assign node832 = (inp[11]) ? 3'b000 : 3'b100;
										assign node836 = (inp[8]) ? node838 : 3'b000;
											assign node838 = (inp[11]) ? 3'b000 : 3'b100;
									assign node841 = (inp[8]) ? node847 : node842;
										assign node842 = (inp[11]) ? node844 : 3'b100;
											assign node844 = (inp[5]) ? 3'b000 : 3'b100;
										assign node847 = (inp[5]) ? node855 : node848;
											assign node848 = (inp[2]) ? node852 : node849;
												assign node849 = (inp[11]) ? 3'b010 : 3'b110;
												assign node852 = (inp[11]) ? 3'b010 : 3'b000;
											assign node855 = (inp[11]) ? 3'b100 : node856;
												assign node856 = (inp[2]) ? 3'b100 : 3'b010;
						assign node860 = (inp[7]) ? node870 : node861;
							assign node861 = (inp[1]) ? 3'b000 : node862;
								assign node862 = (inp[2]) ? node864 : 3'b000;
									assign node864 = (inp[11]) ? 3'b000 : node865;
										assign node865 = (inp[10]) ? 3'b000 : 3'b100;
							assign node870 = (inp[11]) ? node902 : node871;
								assign node871 = (inp[10]) ? node887 : node872;
									assign node872 = (inp[1]) ? node882 : node873;
										assign node873 = (inp[5]) ? node877 : node874;
											assign node874 = (inp[8]) ? 3'b110 : 3'b010;
											assign node877 = (inp[2]) ? node879 : 3'b010;
												assign node879 = (inp[8]) ? 3'b110 : 3'b100;
										assign node882 = (inp[8]) ? 3'b100 : node883;
											assign node883 = (inp[5]) ? 3'b000 : 3'b100;
									assign node887 = (inp[1]) ? 3'b000 : node888;
										assign node888 = (inp[2]) ? node896 : node889;
											assign node889 = (inp[5]) ? node893 : node890;
												assign node890 = (inp[8]) ? 3'b000 : 3'b100;
												assign node893 = (inp[8]) ? 3'b100 : 3'b000;
											assign node896 = (inp[8]) ? 3'b100 : node897;
												assign node897 = (inp[5]) ? 3'b000 : 3'b100;
								assign node902 = (inp[5]) ? 3'b000 : node903;
									assign node903 = (inp[1]) ? node913 : node904;
										assign node904 = (inp[8]) ? node908 : node905;
											assign node905 = (inp[10]) ? 3'b000 : 3'b100;
											assign node908 = (inp[10]) ? 3'b100 : node909;
												assign node909 = (inp[2]) ? 3'b010 : 3'b000;
										assign node913 = (inp[2]) ? node915 : 3'b000;
											assign node915 = (inp[8]) ? 3'b100 : 3'b000;
			assign node919 = (inp[9]) ? node1173 : node920;
				assign node920 = (inp[7]) ? node1002 : node921;
					assign node921 = (inp[4]) ? node987 : node922;
						assign node922 = (inp[10]) ? node968 : node923;
							assign node923 = (inp[11]) ? node943 : node924;
								assign node924 = (inp[1]) ? node930 : node925;
									assign node925 = (inp[8]) ? 3'b100 : node926;
										assign node926 = (inp[5]) ? 3'b000 : 3'b100;
									assign node930 = (inp[0]) ? node936 : node931;
										assign node931 = (inp[5]) ? node933 : 3'b010;
											assign node933 = (inp[8]) ? 3'b010 : 3'b100;
										assign node936 = (inp[5]) ? 3'b000 : node937;
											assign node937 = (inp[2]) ? node939 : 3'b000;
												assign node939 = (inp[8]) ? 3'b100 : 3'b000;
								assign node943 = (inp[2]) ? node951 : node944;
									assign node944 = (inp[0]) ? 3'b000 : node945;
										assign node945 = (inp[5]) ? 3'b000 : node946;
											assign node946 = (inp[8]) ? 3'b000 : 3'b100;
									assign node951 = (inp[5]) ? node961 : node952;
										assign node952 = (inp[1]) ? node956 : node953;
											assign node953 = (inp[8]) ? 3'b100 : 3'b000;
											assign node956 = (inp[8]) ? node958 : 3'b100;
												assign node958 = (inp[0]) ? 3'b000 : 3'b010;
										assign node961 = (inp[1]) ? node963 : 3'b000;
											assign node963 = (inp[0]) ? 3'b000 : node964;
												assign node964 = (inp[8]) ? 3'b100 : 3'b000;
							assign node968 = (inp[0]) ? 3'b000 : node969;
								assign node969 = (inp[1]) ? node971 : 3'b000;
									assign node971 = (inp[8]) ? node977 : node972;
										assign node972 = (inp[11]) ? 3'b000 : node973;
											assign node973 = (inp[5]) ? 3'b000 : 3'b100;
										assign node977 = (inp[11]) ? node983 : node978;
											assign node978 = (inp[2]) ? 3'b100 : node979;
												assign node979 = (inp[5]) ? 3'b100 : 3'b000;
											assign node983 = (inp[5]) ? 3'b000 : 3'b100;
						assign node987 = (inp[11]) ? 3'b000 : node988;
							assign node988 = (inp[1]) ? node990 : 3'b000;
								assign node990 = (inp[2]) ? node992 : 3'b000;
									assign node992 = (inp[5]) ? 3'b000 : node993;
										assign node993 = (inp[0]) ? 3'b000 : node994;
											assign node994 = (inp[8]) ? node996 : 3'b000;
												assign node996 = (inp[10]) ? 3'b000 : 3'b100;
					assign node1002 = (inp[4]) ? node1118 : node1003;
						assign node1003 = (inp[0]) ? node1077 : node1004;
							assign node1004 = (inp[5]) ? node1048 : node1005;
								assign node1005 = (inp[1]) ? node1021 : node1006;
									assign node1006 = (inp[10]) ? node1014 : node1007;
										assign node1007 = (inp[2]) ? node1009 : 3'b100;
											assign node1009 = (inp[8]) ? node1011 : 3'b000;
												assign node1011 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1014 = (inp[2]) ? node1016 : 3'b000;
											assign node1016 = (inp[8]) ? node1018 : 3'b110;
												assign node1018 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1021 = (inp[10]) ? node1035 : node1022;
										assign node1022 = (inp[2]) ? node1028 : node1023;
											assign node1023 = (inp[8]) ? 3'b000 : node1024;
												assign node1024 = (inp[11]) ? 3'b000 : 3'b010;
											assign node1028 = (inp[11]) ? node1032 : node1029;
												assign node1029 = (inp[8]) ? 3'b001 : 3'b110;
												assign node1032 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1035 = (inp[2]) ? node1043 : node1036;
											assign node1036 = (inp[11]) ? node1040 : node1037;
												assign node1037 = (inp[8]) ? 3'b110 : 3'b010;
												assign node1040 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1043 = (inp[8]) ? node1045 : 3'b010;
												assign node1045 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1048 = (inp[10]) ? node1062 : node1049;
									assign node1049 = (inp[11]) ? node1055 : node1050;
										assign node1050 = (inp[1]) ? node1052 : 3'b110;
											assign node1052 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1055 = (inp[1]) ? node1059 : node1056;
											assign node1056 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1059 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1062 = (inp[8]) ? node1072 : node1063;
										assign node1063 = (inp[1]) ? node1067 : node1064;
											assign node1064 = (inp[11]) ? 3'b010 : 3'b100;
											assign node1067 = (inp[2]) ? 3'b100 : node1068;
												assign node1068 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1072 = (inp[1]) ? node1074 : 3'b110;
											assign node1074 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1077 = (inp[10]) ? node1099 : node1078;
								assign node1078 = (inp[1]) ? node1086 : node1079;
									assign node1079 = (inp[8]) ? node1083 : node1080;
										assign node1080 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1083 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1086 = (inp[11]) ? 3'b100 : node1087;
										assign node1087 = (inp[8]) ? node1093 : node1088;
											assign node1088 = (inp[5]) ? 3'b100 : node1089;
												assign node1089 = (inp[2]) ? 3'b100 : 3'b000;
											assign node1093 = (inp[2]) ? node1095 : 3'b010;
												assign node1095 = (inp[5]) ? 3'b100 : 3'b010;
								assign node1099 = (inp[1]) ? node1113 : node1100;
									assign node1100 = (inp[11]) ? node1102 : 3'b100;
										assign node1102 = (inp[2]) ? node1108 : node1103;
											assign node1103 = (inp[8]) ? 3'b000 : node1104;
												assign node1104 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1108 = (inp[5]) ? node1110 : 3'b100;
												assign node1110 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1113 = (inp[11]) ? 3'b000 : node1114;
										assign node1114 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1118 = (inp[0]) ? node1162 : node1119;
							assign node1119 = (inp[1]) ? node1133 : node1120;
								assign node1120 = (inp[10]) ? 3'b000 : node1121;
									assign node1121 = (inp[11]) ? node1127 : node1122;
										assign node1122 = (inp[8]) ? 3'b100 : node1123;
											assign node1123 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1127 = (inp[2]) ? node1129 : 3'b000;
											assign node1129 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1133 = (inp[10]) ? node1149 : node1134;
									assign node1134 = (inp[11]) ? node1140 : node1135;
										assign node1135 = (inp[5]) ? node1137 : 3'b010;
											assign node1137 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1140 = (inp[5]) ? node1146 : node1141;
											assign node1141 = (inp[8]) ? node1143 : 3'b100;
												assign node1143 = (inp[2]) ? 3'b010 : 3'b000;
											assign node1146 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1149 = (inp[8]) ? node1155 : node1150;
										assign node1150 = (inp[11]) ? 3'b000 : node1151;
											assign node1151 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1155 = (inp[2]) ? 3'b100 : node1156;
											assign node1156 = (inp[5]) ? 3'b100 : node1157;
												assign node1157 = (inp[11]) ? 3'b100 : 3'b000;
							assign node1162 = (inp[10]) ? 3'b000 : node1163;
								assign node1163 = (inp[1]) ? 3'b000 : node1164;
									assign node1164 = (inp[11]) ? 3'b000 : node1165;
										assign node1165 = (inp[8]) ? 3'b100 : node1166;
											assign node1166 = (inp[5]) ? 3'b000 : 3'b100;
				assign node1173 = (inp[7]) ? node1175 : 3'b000;
					assign node1175 = (inp[0]) ? 3'b000 : node1176;
						assign node1176 = (inp[4]) ? 3'b000 : node1177;
							assign node1177 = (inp[1]) ? node1183 : node1178;
								assign node1178 = (inp[5]) ? node1180 : 3'b010;
									assign node1180 = (inp[10]) ? 3'b000 : 3'b010;
								assign node1183 = (inp[10]) ? 3'b000 : node1184;
									assign node1184 = (inp[5]) ? node1192 : node1185;
										assign node1185 = (inp[11]) ? 3'b100 : node1186;
											assign node1186 = (inp[8]) ? node1188 : 3'b100;
												assign node1188 = (inp[2]) ? 3'b010 : 3'b000;
										assign node1192 = (inp[8]) ? node1194 : 3'b000;
											assign node1194 = (inp[11]) ? 3'b000 : 3'b100;
		assign node1200 = (inp[3]) ? node2076 : node1201;
			assign node1201 = (inp[9]) ? node1551 : node1202;
				assign node1202 = (inp[0]) ? node1326 : node1203;
					assign node1203 = (inp[1]) ? node1225 : node1204;
						assign node1204 = (inp[7]) ? 3'b111 : node1205;
							assign node1205 = (inp[4]) ? node1207 : 3'b111;
								assign node1207 = (inp[11]) ? node1213 : node1208;
									assign node1208 = (inp[5]) ? node1210 : 3'b111;
										assign node1210 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1213 = (inp[10]) ? node1219 : node1214;
										assign node1214 = (inp[5]) ? node1216 : 3'b111;
											assign node1216 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1219 = (inp[2]) ? node1221 : 3'b011;
											assign node1221 = (inp[5]) ? 3'b111 : 3'b011;
						assign node1225 = (inp[7]) ? node1303 : node1226;
							assign node1226 = (inp[4]) ? node1272 : node1227;
								assign node1227 = (inp[11]) ? node1247 : node1228;
									assign node1228 = (inp[10]) ? node1238 : node1229;
										assign node1229 = (inp[8]) ? node1231 : 3'b111;
											assign node1231 = (inp[5]) ? node1235 : node1232;
												assign node1232 = (inp[2]) ? 3'b011 : 3'b111;
												assign node1235 = (inp[2]) ? 3'b111 : 3'b011;
										assign node1238 = (inp[8]) ? node1240 : 3'b011;
											assign node1240 = (inp[2]) ? node1244 : node1241;
												assign node1241 = (inp[5]) ? 3'b111 : 3'b011;
												assign node1244 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1247 = (inp[2]) ? node1259 : node1248;
										assign node1248 = (inp[10]) ? node1252 : node1249;
											assign node1249 = (inp[5]) ? 3'b011 : 3'b010;
											assign node1252 = (inp[5]) ? node1256 : node1253;
												assign node1253 = (inp[8]) ? 3'b111 : 3'b011;
												assign node1256 = (inp[8]) ? 3'b011 : 3'b010;
										assign node1259 = (inp[5]) ? node1267 : node1260;
											assign node1260 = (inp[10]) ? node1264 : node1261;
												assign node1261 = (inp[8]) ? 3'b011 : 3'b111;
												assign node1264 = (inp[8]) ? 3'b111 : 3'b011;
											assign node1267 = (inp[10]) ? node1269 : 3'b011;
												assign node1269 = (inp[8]) ? 3'b011 : 3'b110;
								assign node1272 = (inp[10]) ? node1292 : node1273;
									assign node1273 = (inp[8]) ? node1281 : node1274;
										assign node1274 = (inp[11]) ? 3'b101 : node1275;
											assign node1275 = (inp[5]) ? 3'b101 : node1276;
												assign node1276 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1281 = (inp[2]) ? node1287 : node1282;
											assign node1282 = (inp[5]) ? 3'b011 : node1283;
												assign node1283 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1287 = (inp[5]) ? 3'b101 : node1288;
												assign node1288 = (inp[11]) ? 3'b011 : 3'b111;
									assign node1292 = (inp[11]) ? node1298 : node1293;
										assign node1293 = (inp[8]) ? node1295 : 3'b101;
											assign node1295 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1298 = (inp[8]) ? node1300 : 3'b001;
											assign node1300 = (inp[2]) ? 3'b001 : 3'b101;
							assign node1303 = (inp[4]) ? node1305 : 3'b111;
								assign node1305 = (inp[8]) ? node1317 : node1306;
									assign node1306 = (inp[11]) ? node1310 : node1307;
										assign node1307 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1310 = (inp[5]) ? node1314 : node1311;
											assign node1311 = (inp[10]) ? 3'b011 : 3'b101;
											assign node1314 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1317 = (inp[5]) ? node1319 : 3'b111;
										assign node1319 = (inp[10]) ? node1321 : 3'b111;
											assign node1321 = (inp[2]) ? 3'b011 : node1322;
												assign node1322 = (inp[11]) ? 3'b011 : 3'b111;
					assign node1326 = (inp[4]) ? node1436 : node1327;
						assign node1327 = (inp[7]) ? node1401 : node1328;
							assign node1328 = (inp[1]) ? node1360 : node1329;
								assign node1329 = (inp[11]) ? node1345 : node1330;
									assign node1330 = (inp[10]) ? node1334 : node1331;
										assign node1331 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1334 = (inp[2]) ? node1340 : node1335;
											assign node1335 = (inp[5]) ? node1337 : 3'b111;
												assign node1337 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1340 = (inp[5]) ? 3'b101 : node1341;
												assign node1341 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1345 = (inp[8]) ? node1355 : node1346;
										assign node1346 = (inp[10]) ? node1350 : node1347;
											assign node1347 = (inp[5]) ? 3'b101 : 3'b111;
											assign node1350 = (inp[5]) ? node1352 : 3'b101;
												assign node1352 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1355 = (inp[5]) ? 3'b011 : node1356;
											assign node1356 = (inp[10]) ? 3'b011 : 3'b111;
								assign node1360 = (inp[10]) ? node1382 : node1361;
									assign node1361 = (inp[11]) ? node1367 : node1362;
										assign node1362 = (inp[5]) ? 3'b011 : node1363;
											assign node1363 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1367 = (inp[8]) ? node1375 : node1368;
											assign node1368 = (inp[5]) ? node1372 : node1369;
												assign node1369 = (inp[2]) ? 3'b101 : 3'b001;
												assign node1372 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1375 = (inp[5]) ? node1379 : node1376;
												assign node1376 = (inp[2]) ? 3'b011 : 3'b010;
												assign node1379 = (inp[2]) ? 3'b101 : 3'b001;
									assign node1382 = (inp[5]) ? node1394 : node1383;
										assign node1383 = (inp[11]) ? node1389 : node1384;
											assign node1384 = (inp[2]) ? 3'b101 : node1385;
												assign node1385 = (inp[8]) ? 3'b001 : 3'b101;
											assign node1389 = (inp[8]) ? 3'b001 : node1390;
												assign node1390 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1394 = (inp[11]) ? node1398 : node1395;
											assign node1395 = (inp[8]) ? 3'b101 : 3'b001;
											assign node1398 = (inp[8]) ? 3'b001 : 3'b110;
							assign node1401 = (inp[1]) ? node1411 : node1402;
								assign node1402 = (inp[11]) ? node1404 : 3'b111;
									assign node1404 = (inp[10]) ? node1406 : 3'b111;
										assign node1406 = (inp[2]) ? 3'b011 : node1407;
											assign node1407 = (inp[8]) ? 3'b111 : 3'b011;
								assign node1411 = (inp[11]) ? node1427 : node1412;
									assign node1412 = (inp[5]) ? node1420 : node1413;
										assign node1413 = (inp[2]) ? node1415 : 3'b101;
											assign node1415 = (inp[10]) ? node1417 : 3'b111;
												assign node1417 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1420 = (inp[8]) ? node1424 : node1421;
											assign node1421 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1424 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1427 = (inp[2]) ? 3'b011 : node1428;
										assign node1428 = (inp[10]) ? node1432 : node1429;
											assign node1429 = (inp[5]) ? 3'b111 : 3'b011;
											assign node1432 = (inp[5]) ? 3'b001 : 3'b111;
						assign node1436 = (inp[7]) ? node1492 : node1437;
							assign node1437 = (inp[1]) ? node1467 : node1438;
								assign node1438 = (inp[10]) ? node1450 : node1439;
									assign node1439 = (inp[8]) ? node1447 : node1440;
										assign node1440 = (inp[5]) ? 3'b001 : node1441;
											assign node1441 = (inp[2]) ? node1443 : 3'b001;
												assign node1443 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1447 = (inp[5]) ? 3'b101 : 3'b011;
									assign node1450 = (inp[11]) ? node1458 : node1451;
										assign node1451 = (inp[5]) ? node1455 : node1452;
											assign node1452 = (inp[8]) ? 3'b101 : 3'b001;
											assign node1455 = (inp[8]) ? 3'b001 : 3'b010;
										assign node1458 = (inp[5]) ? 3'b110 : node1459;
											assign node1459 = (inp[8]) ? node1463 : node1460;
												assign node1460 = (inp[2]) ? 3'b110 : 3'b000;
												assign node1463 = (inp[2]) ? 3'b001 : 3'b101;
								assign node1467 = (inp[8]) ? node1483 : node1468;
									assign node1468 = (inp[2]) ? node1476 : node1469;
										assign node1469 = (inp[11]) ? node1471 : 3'b110;
											assign node1471 = (inp[10]) ? node1473 : 3'b110;
												assign node1473 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1476 = (inp[5]) ? node1480 : node1477;
											assign node1477 = (inp[10]) ? 3'b110 : 3'b001;
											assign node1480 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1483 = (inp[10]) ? node1487 : node1484;
										assign node1484 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1487 = (inp[5]) ? 3'b110 : node1488;
											assign node1488 = (inp[2]) ? 3'b001 : 3'b010;
							assign node1492 = (inp[1]) ? node1528 : node1493;
								assign node1493 = (inp[5]) ? node1509 : node1494;
									assign node1494 = (inp[2]) ? node1504 : node1495;
										assign node1495 = (inp[10]) ? node1501 : node1496;
											assign node1496 = (inp[11]) ? 3'b111 : node1497;
												assign node1497 = (inp[8]) ? 3'b111 : 3'b011;
											assign node1501 = (inp[8]) ? 3'b011 : 3'b111;
										assign node1504 = (inp[8]) ? node1506 : 3'b011;
											assign node1506 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1509 = (inp[10]) ? node1519 : node1510;
										assign node1510 = (inp[8]) ? node1514 : node1511;
											assign node1511 = (inp[11]) ? 3'b101 : 3'b011;
											assign node1514 = (inp[11]) ? 3'b011 : node1515;
												assign node1515 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1519 = (inp[2]) ? node1523 : node1520;
											assign node1520 = (inp[11]) ? 3'b101 : 3'b011;
											assign node1523 = (inp[8]) ? 3'b101 : node1524;
												assign node1524 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1528 = (inp[11]) ? node1536 : node1529;
									assign node1529 = (inp[10]) ? node1533 : node1530;
										assign node1530 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1533 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1536 = (inp[8]) ? node1546 : node1537;
										assign node1537 = (inp[5]) ? node1541 : node1538;
											assign node1538 = (inp[10]) ? 3'b001 : 3'b101;
											assign node1541 = (inp[10]) ? node1543 : 3'b001;
												assign node1543 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1546 = (inp[2]) ? node1548 : 3'b101;
											assign node1548 = (inp[5]) ? 3'b101 : 3'b011;
				assign node1551 = (inp[0]) ? node1815 : node1552;
					assign node1552 = (inp[4]) ? node1686 : node1553;
						assign node1553 = (inp[7]) ? node1627 : node1554;
							assign node1554 = (inp[1]) ? node1596 : node1555;
								assign node1555 = (inp[8]) ? node1577 : node1556;
									assign node1556 = (inp[2]) ? node1568 : node1557;
										assign node1557 = (inp[5]) ? node1563 : node1558;
											assign node1558 = (inp[11]) ? 3'b011 : node1559;
												assign node1559 = (inp[10]) ? 3'b011 : 3'b101;
											assign node1563 = (inp[10]) ? 3'b101 : node1564;
												assign node1564 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1568 = (inp[11]) ? node1572 : node1569;
											assign node1569 = (inp[10]) ? 3'b111 : 3'b101;
											assign node1572 = (inp[10]) ? node1574 : 3'b101;
												assign node1574 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1577 = (inp[10]) ? node1589 : node1578;
										assign node1578 = (inp[5]) ? node1584 : node1579;
											assign node1579 = (inp[2]) ? node1581 : 3'b111;
												assign node1581 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1584 = (inp[11]) ? 3'b011 : node1585;
												assign node1585 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1589 = (inp[11]) ? node1591 : 3'b011;
											assign node1591 = (inp[5]) ? 3'b101 : node1592;
												assign node1592 = (inp[2]) ? 3'b111 : 3'b011;
								assign node1596 = (inp[10]) ? node1612 : node1597;
									assign node1597 = (inp[5]) ? node1603 : node1598;
										assign node1598 = (inp[8]) ? 3'b011 : node1599;
											assign node1599 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1603 = (inp[11]) ? node1609 : node1604;
											assign node1604 = (inp[2]) ? 3'b101 : node1605;
												assign node1605 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1609 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1612 = (inp[8]) ? node1618 : node1613;
										assign node1613 = (inp[11]) ? node1615 : 3'b001;
											assign node1615 = (inp[2]) ? 3'b111 : 3'b001;
										assign node1618 = (inp[5]) ? node1624 : node1619;
											assign node1619 = (inp[2]) ? 3'b101 : node1620;
												assign node1620 = (inp[11]) ? 3'b101 : 3'b001;
											assign node1624 = (inp[11]) ? 3'b001 : 3'b101;
							assign node1627 = (inp[10]) ? node1653 : node1628;
								assign node1628 = (inp[8]) ? node1644 : node1629;
									assign node1629 = (inp[11]) ? node1635 : node1630;
										assign node1630 = (inp[1]) ? node1632 : 3'b111;
											assign node1632 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1635 = (inp[5]) ? node1641 : node1636;
											assign node1636 = (inp[1]) ? node1638 : 3'b011;
												assign node1638 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1641 = (inp[2]) ? 3'b111 : 3'b011;
									assign node1644 = (inp[11]) ? node1646 : 3'b111;
										assign node1646 = (inp[1]) ? node1648 : 3'b111;
											assign node1648 = (inp[2]) ? node1650 : 3'b111;
												assign node1650 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1653 = (inp[1]) ? node1667 : node1654;
									assign node1654 = (inp[8]) ? node1660 : node1655;
										assign node1655 = (inp[11]) ? node1657 : 3'b011;
											assign node1657 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1660 = (inp[11]) ? 3'b111 : node1661;
											assign node1661 = (inp[2]) ? node1663 : 3'b111;
												assign node1663 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1667 = (inp[8]) ? node1675 : node1668;
										assign node1668 = (inp[5]) ? 3'b101 : node1669;
											assign node1669 = (inp[11]) ? node1671 : 3'b001;
												assign node1671 = (inp[2]) ? 3'b111 : 3'b011;
										assign node1675 = (inp[5]) ? node1679 : node1676;
											assign node1676 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1679 = (inp[11]) ? node1683 : node1680;
												assign node1680 = (inp[2]) ? 3'b001 : 3'b011;
												assign node1683 = (inp[2]) ? 3'b111 : 3'b011;
						assign node1686 = (inp[7]) ? node1748 : node1687;
							assign node1687 = (inp[1]) ? node1715 : node1688;
								assign node1688 = (inp[10]) ? node1700 : node1689;
									assign node1689 = (inp[11]) ? 3'b101 : node1690;
										assign node1690 = (inp[8]) ? node1692 : 3'b001;
											assign node1692 = (inp[2]) ? node1696 : node1693;
												assign node1693 = (inp[5]) ? 3'b101 : 3'b011;
												assign node1696 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1700 = (inp[11]) ? node1710 : node1701;
										assign node1701 = (inp[8]) ? node1703 : 3'b110;
											assign node1703 = (inp[2]) ? node1707 : node1704;
												assign node1704 = (inp[5]) ? 3'b001 : 3'b101;
												assign node1707 = (inp[5]) ? 3'b110 : 3'b011;
										assign node1710 = (inp[8]) ? node1712 : 3'b000;
											assign node1712 = (inp[5]) ? 3'b000 : 3'b001;
								assign node1715 = (inp[8]) ? node1733 : node1716;
									assign node1716 = (inp[11]) ? node1724 : node1717;
										assign node1717 = (inp[5]) ? node1719 : 3'b110;
											assign node1719 = (inp[10]) ? node1721 : 3'b110;
												assign node1721 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1724 = (inp[10]) ? node1730 : node1725;
											assign node1725 = (inp[5]) ? 3'b110 : node1726;
												assign node1726 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1730 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1733 = (inp[5]) ? node1743 : node1734;
										assign node1734 = (inp[2]) ? node1736 : 3'b001;
											assign node1736 = (inp[11]) ? node1740 : node1737;
												assign node1737 = (inp[10]) ? 3'b001 : 3'b101;
												assign node1740 = (inp[10]) ? 3'b110 : 3'b001;
										assign node1743 = (inp[2]) ? 3'b110 : node1744;
											assign node1744 = (inp[10]) ? 3'b110 : 3'b001;
							assign node1748 = (inp[10]) ? node1780 : node1749;
								assign node1749 = (inp[11]) ? node1759 : node1750;
									assign node1750 = (inp[2]) ? 3'b011 : node1751;
										assign node1751 = (inp[1]) ? node1753 : 3'b111;
											assign node1753 = (inp[5]) ? node1755 : 3'b011;
												assign node1755 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1759 = (inp[5]) ? node1771 : node1760;
										assign node1760 = (inp[1]) ? node1766 : node1761;
											assign node1761 = (inp[8]) ? node1763 : 3'b011;
												assign node1763 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1766 = (inp[8]) ? 3'b011 : node1767;
												assign node1767 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1771 = (inp[2]) ? node1775 : node1772;
											assign node1772 = (inp[8]) ? 3'b011 : 3'b101;
											assign node1775 = (inp[1]) ? node1777 : 3'b101;
												assign node1777 = (inp[8]) ? 3'b101 : 3'b001;
								assign node1780 = (inp[1]) ? node1802 : node1781;
									assign node1781 = (inp[8]) ? node1791 : node1782;
										assign node1782 = (inp[5]) ? node1788 : node1783;
											assign node1783 = (inp[2]) ? 3'b101 : node1784;
												assign node1784 = (inp[11]) ? 3'b101 : 3'b011;
											assign node1788 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1791 = (inp[11]) ? node1797 : node1792;
											assign node1792 = (inp[5]) ? node1794 : 3'b011;
												assign node1794 = (inp[2]) ? 3'b111 : 3'b011;
											assign node1797 = (inp[5]) ? 3'b101 : node1798;
												assign node1798 = (inp[2]) ? 3'b111 : 3'b011;
									assign node1802 = (inp[5]) ? node1808 : node1803;
										assign node1803 = (inp[11]) ? node1805 : 3'b101;
											assign node1805 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1808 = (inp[2]) ? node1810 : 3'b001;
											assign node1810 = (inp[11]) ? node1812 : 3'b001;
												assign node1812 = (inp[8]) ? 3'b000 : 3'b110;
					assign node1815 = (inp[7]) ? node1935 : node1816;
						assign node1816 = (inp[4]) ? node1880 : node1817;
							assign node1817 = (inp[10]) ? node1851 : node1818;
								assign node1818 = (inp[1]) ? node1830 : node1819;
									assign node1819 = (inp[11]) ? node1823 : node1820;
										assign node1820 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1823 = (inp[2]) ? node1827 : node1824;
											assign node1824 = (inp[8]) ? 3'b001 : 3'b101;
											assign node1827 = (inp[8]) ? 3'b101 : 3'b110;
									assign node1830 = (inp[11]) ? node1836 : node1831;
										assign node1831 = (inp[5]) ? node1833 : 3'b001;
											assign node1833 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1836 = (inp[8]) ? node1844 : node1837;
											assign node1837 = (inp[2]) ? node1841 : node1838;
												assign node1838 = (inp[5]) ? 3'b110 : 3'b010;
												assign node1841 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1844 = (inp[5]) ? node1848 : node1845;
												assign node1845 = (inp[2]) ? 3'b001 : 3'b000;
												assign node1848 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1851 = (inp[8]) ? node1857 : node1852;
									assign node1852 = (inp[5]) ? node1854 : 3'b110;
										assign node1854 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1857 = (inp[1]) ? node1871 : node1858;
										assign node1858 = (inp[5]) ? node1866 : node1859;
											assign node1859 = (inp[2]) ? node1863 : node1860;
												assign node1860 = (inp[11]) ? 3'b001 : 3'b101;
												assign node1863 = (inp[11]) ? 3'b001 : 3'b011;
											assign node1866 = (inp[11]) ? 3'b110 : node1867;
												assign node1867 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1871 = (inp[11]) ? node1877 : node1872;
											assign node1872 = (inp[2]) ? 3'b110 : node1873;
												assign node1873 = (inp[5]) ? 3'b110 : 3'b010;
											assign node1877 = (inp[5]) ? 3'b010 : 3'b110;
							assign node1880 = (inp[10]) ? node1906 : node1881;
								assign node1881 = (inp[1]) ? node1895 : node1882;
									assign node1882 = (inp[5]) ? node1892 : node1883;
										assign node1883 = (inp[2]) ? node1889 : node1884;
											assign node1884 = (inp[8]) ? 3'b001 : node1885;
												assign node1885 = (inp[11]) ? 3'b101 : 3'b010;
											assign node1889 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1892 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1895 = (inp[5]) ? node1903 : node1896;
										assign node1896 = (inp[8]) ? 3'b110 : node1897;
											assign node1897 = (inp[2]) ? 3'b010 : node1898;
												assign node1898 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1903 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1906 = (inp[1]) ? node1922 : node1907;
									assign node1907 = (inp[2]) ? node1915 : node1908;
										assign node1908 = (inp[8]) ? node1912 : node1909;
											assign node1909 = (inp[5]) ? 3'b100 : 3'b010;
											assign node1912 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1915 = (inp[8]) ? node1917 : 3'b100;
											assign node1917 = (inp[11]) ? 3'b100 : node1918;
												assign node1918 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1922 = (inp[2]) ? node1930 : node1923;
										assign node1923 = (inp[8]) ? node1927 : node1924;
											assign node1924 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1927 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1930 = (inp[8]) ? 3'b100 : node1931;
											assign node1931 = (inp[5]) ? 3'b000 : 3'b100;
						assign node1935 = (inp[10]) ? node2009 : node1936;
							assign node1936 = (inp[4]) ? node1976 : node1937;
								assign node1937 = (inp[8]) ? node1957 : node1938;
									assign node1938 = (inp[1]) ? node1946 : node1939;
										assign node1939 = (inp[5]) ? 3'b101 : node1940;
											assign node1940 = (inp[11]) ? node1942 : 3'b111;
												assign node1942 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1946 = (inp[2]) ? node1952 : node1947;
											assign node1947 = (inp[11]) ? node1949 : 3'b001;
												assign node1949 = (inp[5]) ? 3'b001 : 3'b011;
											assign node1952 = (inp[5]) ? 3'b001 : node1953;
												assign node1953 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1957 = (inp[1]) ? node1965 : node1958;
										assign node1958 = (inp[5]) ? node1962 : node1959;
											assign node1959 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1962 = (inp[2]) ? 3'b101 : 3'b011;
										assign node1965 = (inp[5]) ? node1971 : node1966;
											assign node1966 = (inp[11]) ? node1968 : 3'b011;
												assign node1968 = (inp[2]) ? 3'b101 : 3'b111;
											assign node1971 = (inp[2]) ? node1973 : 3'b101;
												assign node1973 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1976 = (inp[11]) ? node1996 : node1977;
									assign node1977 = (inp[8]) ? node1983 : node1978;
										assign node1978 = (inp[5]) ? node1980 : 3'b001;
											assign node1980 = (inp[1]) ? 3'b110 : 3'b001;
										assign node1983 = (inp[1]) ? node1991 : node1984;
											assign node1984 = (inp[2]) ? node1988 : node1985;
												assign node1985 = (inp[5]) ? 3'b101 : 3'b011;
												assign node1988 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1991 = (inp[5]) ? 3'b001 : node1992;
												assign node1992 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1996 = (inp[8]) ? node2004 : node1997;
										assign node1997 = (inp[5]) ? 3'b110 : node1998;
											assign node1998 = (inp[1]) ? 3'b110 : node1999;
												assign node1999 = (inp[2]) ? 3'b001 : 3'b101;
										assign node2004 = (inp[1]) ? 3'b001 : node2005;
											assign node2005 = (inp[5]) ? 3'b001 : 3'b101;
							assign node2009 = (inp[4]) ? node2045 : node2010;
								assign node2010 = (inp[1]) ? node2030 : node2011;
									assign node2011 = (inp[11]) ? node2023 : node2012;
										assign node2012 = (inp[2]) ? node2018 : node2013;
											assign node2013 = (inp[5]) ? 3'b101 : node2014;
												assign node2014 = (inp[8]) ? 3'b011 : 3'b101;
											assign node2018 = (inp[5]) ? node2020 : 3'b011;
												assign node2020 = (inp[8]) ? 3'b101 : 3'b011;
										assign node2023 = (inp[8]) ? node2027 : node2024;
											assign node2024 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2027 = (inp[2]) ? 3'b101 : 3'b011;
									assign node2030 = (inp[5]) ? node2036 : node2031;
										assign node2031 = (inp[2]) ? 3'b001 : node2032;
											assign node2032 = (inp[8]) ? 3'b101 : 3'b100;
										assign node2036 = (inp[8]) ? node2040 : node2037;
											assign node2037 = (inp[11]) ? 3'b110 : 3'b010;
											assign node2040 = (inp[11]) ? node2042 : 3'b001;
												assign node2042 = (inp[2]) ? 3'b110 : 3'b001;
								assign node2045 = (inp[8]) ? node2063 : node2046;
									assign node2046 = (inp[5]) ? node2054 : node2047;
										assign node2047 = (inp[1]) ? node2049 : 3'b110;
											assign node2049 = (inp[2]) ? node2051 : 3'b110;
												assign node2051 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2054 = (inp[1]) ? node2058 : node2055;
											assign node2055 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2058 = (inp[11]) ? node2060 : 3'b010;
												assign node2060 = (inp[2]) ? 3'b100 : 3'b000;
									assign node2063 = (inp[1]) ? node2073 : node2064;
										assign node2064 = (inp[5]) ? node2068 : node2065;
											assign node2065 = (inp[11]) ? 3'b001 : 3'b011;
											assign node2068 = (inp[2]) ? 3'b110 : node2069;
												assign node2069 = (inp[11]) ? 3'b110 : 3'b001;
										assign node2073 = (inp[2]) ? 3'b110 : 3'b010;
			assign node2076 = (inp[9]) ? node2530 : node2077;
				assign node2077 = (inp[7]) ? node2303 : node2078;
					assign node2078 = (inp[4]) ? node2194 : node2079;
						assign node2079 = (inp[10]) ? node2145 : node2080;
							assign node2080 = (inp[5]) ? node2120 : node2081;
								assign node2081 = (inp[0]) ? node2097 : node2082;
									assign node2082 = (inp[1]) ? node2088 : node2083;
										assign node2083 = (inp[2]) ? 3'b101 : node2084;
											assign node2084 = (inp[8]) ? 3'b111 : 3'b101;
										assign node2088 = (inp[11]) ? node2092 : node2089;
											assign node2089 = (inp[8]) ? 3'b011 : 3'b001;
											assign node2092 = (inp[8]) ? 3'b101 : node2093;
												assign node2093 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2097 = (inp[1]) ? node2107 : node2098;
										assign node2098 = (inp[8]) ? node2104 : node2099;
											assign node2099 = (inp[2]) ? node2101 : 3'b001;
												assign node2101 = (inp[11]) ? 3'b101 : 3'b001;
											assign node2104 = (inp[11]) ? 3'b001 : 3'b011;
										assign node2107 = (inp[2]) ? node2115 : node2108;
											assign node2108 = (inp[11]) ? node2112 : node2109;
												assign node2109 = (inp[8]) ? 3'b001 : 3'b111;
												assign node2112 = (inp[8]) ? 3'b110 : 3'b100;
											assign node2115 = (inp[11]) ? node2117 : 3'b110;
												assign node2117 = (inp[8]) ? 3'b110 : 3'b010;
								assign node2120 = (inp[1]) ? node2130 : node2121;
									assign node2121 = (inp[2]) ? 3'b110 : node2122;
										assign node2122 = (inp[8]) ? 3'b100 : node2123;
											assign node2123 = (inp[11]) ? node2125 : 3'b110;
												assign node2125 = (inp[0]) ? 3'b010 : 3'b110;
									assign node2130 = (inp[0]) ? node2140 : node2131;
										assign node2131 = (inp[8]) ? node2135 : node2132;
											assign node2132 = (inp[11]) ? 3'b110 : 3'b001;
											assign node2135 = (inp[11]) ? 3'b001 : node2136;
												assign node2136 = (inp[2]) ? 3'b001 : 3'b101;
										assign node2140 = (inp[8]) ? node2142 : 3'b010;
											assign node2142 = (inp[11]) ? 3'b010 : 3'b110;
							assign node2145 = (inp[5]) ? node2163 : node2146;
								assign node2146 = (inp[8]) ? node2154 : node2147;
									assign node2147 = (inp[0]) ? node2149 : 3'b110;
										assign node2149 = (inp[11]) ? 3'b010 : node2150;
											assign node2150 = (inp[1]) ? 3'b010 : 3'b110;
									assign node2154 = (inp[2]) ? node2158 : node2155;
										assign node2155 = (inp[1]) ? 3'b110 : 3'b100;
										assign node2158 = (inp[1]) ? node2160 : 3'b110;
											assign node2160 = (inp[11]) ? 3'b010 : 3'b001;
								assign node2163 = (inp[8]) ? node2181 : node2164;
									assign node2164 = (inp[0]) ? node2172 : node2165;
										assign node2165 = (inp[1]) ? node2167 : 3'b100;
											assign node2167 = (inp[2]) ? node2169 : 3'b110;
												assign node2169 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2172 = (inp[11]) ? node2174 : 3'b100;
											assign node2174 = (inp[1]) ? node2178 : node2175;
												assign node2175 = (inp[2]) ? 3'b100 : 3'b000;
												assign node2178 = (inp[2]) ? 3'b000 : 3'b100;
									assign node2181 = (inp[0]) ? node2187 : node2182;
										assign node2182 = (inp[11]) ? 3'b110 : node2183;
											assign node2183 = (inp[2]) ? 3'b110 : 3'b001;
										assign node2187 = (inp[11]) ? node2191 : node2188;
											assign node2188 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2191 = (inp[1]) ? 3'b100 : 3'b010;
						assign node2194 = (inp[0]) ? node2248 : node2195;
							assign node2195 = (inp[8]) ? node2215 : node2196;
								assign node2196 = (inp[10]) ? node2200 : node2197;
									assign node2197 = (inp[1]) ? 3'b010 : 3'b110;
									assign node2200 = (inp[1]) ? node2208 : node2201;
										assign node2201 = (inp[11]) ? 3'b010 : node2202;
											assign node2202 = (inp[5]) ? node2204 : 3'b110;
												assign node2204 = (inp[2]) ? 3'b000 : 3'b100;
										assign node2208 = (inp[11]) ? 3'b100 : node2209;
											assign node2209 = (inp[5]) ? node2211 : 3'b010;
												assign node2211 = (inp[2]) ? 3'b100 : 3'b000;
								assign node2215 = (inp[5]) ? node2231 : node2216;
									assign node2216 = (inp[1]) ? node2224 : node2217;
										assign node2217 = (inp[11]) ? node2221 : node2218;
											assign node2218 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2221 = (inp[10]) ? 3'b100 : 3'b000;
										assign node2224 = (inp[10]) ? node2228 : node2225;
											assign node2225 = (inp[11]) ? 3'b100 : 3'b001;
											assign node2228 = (inp[11]) ? 3'b010 : 3'b110;
									assign node2231 = (inp[1]) ? node2243 : node2232;
										assign node2232 = (inp[10]) ? node2238 : node2233;
											assign node2233 = (inp[11]) ? node2235 : 3'b000;
												assign node2235 = (inp[2]) ? 3'b110 : 3'b000;
											assign node2238 = (inp[2]) ? node2240 : 3'b110;
												assign node2240 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2243 = (inp[10]) ? node2245 : 3'b110;
											assign node2245 = (inp[11]) ? 3'b100 : 3'b010;
							assign node2248 = (inp[10]) ? node2280 : node2249;
								assign node2249 = (inp[1]) ? node2265 : node2250;
									assign node2250 = (inp[8]) ? node2258 : node2251;
										assign node2251 = (inp[5]) ? 3'b100 : node2252;
											assign node2252 = (inp[11]) ? 3'b010 : node2253;
												assign node2253 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2258 = (inp[5]) ? 3'b010 : node2259;
											assign node2259 = (inp[2]) ? node2261 : 3'b110;
												assign node2261 = (inp[11]) ? 3'b010 : 3'b110;
									assign node2265 = (inp[2]) ? node2275 : node2266;
										assign node2266 = (inp[8]) ? node2272 : node2267;
											assign node2267 = (inp[5]) ? node2269 : 3'b100;
												assign node2269 = (inp[11]) ? 3'b000 : 3'b100;
											assign node2272 = (inp[11]) ? 3'b100 : 3'b010;
										assign node2275 = (inp[5]) ? node2277 : 3'b100;
											assign node2277 = (inp[8]) ? 3'b100 : 3'b000;
								assign node2280 = (inp[1]) ? node2296 : node2281;
									assign node2281 = (inp[11]) ? node2287 : node2282;
										assign node2282 = (inp[5]) ? 3'b100 : node2283;
											assign node2283 = (inp[8]) ? 3'b010 : 3'b100;
										assign node2287 = (inp[5]) ? node2293 : node2288;
											assign node2288 = (inp[8]) ? node2290 : 3'b100;
												assign node2290 = (inp[2]) ? 3'b100 : 3'b000;
											assign node2293 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2296 = (inp[5]) ? 3'b000 : node2297;
										assign node2297 = (inp[11]) ? 3'b000 : node2298;
											assign node2298 = (inp[8]) ? 3'b100 : 3'b000;
					assign node2303 = (inp[0]) ? node2407 : node2304;
						assign node2304 = (inp[4]) ? node2344 : node2305;
							assign node2305 = (inp[1]) ? node2321 : node2306;
								assign node2306 = (inp[10]) ? node2314 : node2307;
									assign node2307 = (inp[11]) ? node2309 : 3'b111;
										assign node2309 = (inp[2]) ? node2311 : 3'b111;
											assign node2311 = (inp[5]) ? 3'b011 : 3'b111;
									assign node2314 = (inp[11]) ? node2318 : node2315;
										assign node2315 = (inp[5]) ? 3'b011 : 3'b111;
										assign node2318 = (inp[5]) ? 3'b111 : 3'b011;
								assign node2321 = (inp[8]) ? node2333 : node2322;
									assign node2322 = (inp[10]) ? node2328 : node2323;
										assign node2323 = (inp[5]) ? 3'b101 : node2324;
											assign node2324 = (inp[11]) ? 3'b101 : 3'b111;
										assign node2328 = (inp[11]) ? 3'b001 : node2329;
											assign node2329 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2333 = (inp[10]) ? node2339 : node2334;
										assign node2334 = (inp[5]) ? 3'b011 : node2335;
											assign node2335 = (inp[11]) ? 3'b011 : 3'b111;
										assign node2339 = (inp[5]) ? 3'b101 : node2340;
											assign node2340 = (inp[11]) ? 3'b101 : 3'b011;
							assign node2344 = (inp[8]) ? node2378 : node2345;
								assign node2345 = (inp[10]) ? node2365 : node2346;
									assign node2346 = (inp[11]) ? node2354 : node2347;
										assign node2347 = (inp[1]) ? 3'b001 : node2348;
											assign node2348 = (inp[5]) ? node2350 : 3'b011;
												assign node2350 = (inp[2]) ? 3'b101 : 3'b111;
										assign node2354 = (inp[2]) ? node2358 : node2355;
											assign node2355 = (inp[1]) ? 3'b101 : 3'b100;
											assign node2358 = (inp[5]) ? node2362 : node2359;
												assign node2359 = (inp[1]) ? 3'b001 : 3'b100;
												assign node2362 = (inp[1]) ? 3'b110 : 3'b001;
									assign node2365 = (inp[1]) ? node2373 : node2366;
										assign node2366 = (inp[5]) ? node2370 : node2367;
											assign node2367 = (inp[11]) ? 3'b001 : 3'b101;
											assign node2370 = (inp[11]) ? 3'b110 : 3'b001;
										assign node2373 = (inp[11]) ? node2375 : 3'b110;
											assign node2375 = (inp[2]) ? 3'b010 : 3'b110;
								assign node2378 = (inp[10]) ? node2390 : node2379;
									assign node2379 = (inp[5]) ? node2383 : node2380;
										assign node2380 = (inp[1]) ? 3'b101 : 3'b011;
										assign node2383 = (inp[1]) ? node2385 : 3'b101;
											assign node2385 = (inp[2]) ? 3'b001 : node2386;
												assign node2386 = (inp[11]) ? 3'b001 : 3'b101;
									assign node2390 = (inp[1]) ? node2398 : node2391;
										assign node2391 = (inp[5]) ? node2393 : 3'b101;
											assign node2393 = (inp[11]) ? 3'b001 : node2394;
												assign node2394 = (inp[2]) ? 3'b001 : 3'b101;
										assign node2398 = (inp[5]) ? node2402 : node2399;
											assign node2399 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2402 = (inp[11]) ? 3'b110 : node2403;
												assign node2403 = (inp[2]) ? 3'b110 : 3'b001;
						assign node2407 = (inp[4]) ? node2469 : node2408;
							assign node2408 = (inp[10]) ? node2432 : node2409;
								assign node2409 = (inp[1]) ? node2421 : node2410;
									assign node2410 = (inp[5]) ? node2418 : node2411;
										assign node2411 = (inp[2]) ? node2415 : node2412;
											assign node2412 = (inp[8]) ? 3'b011 : 3'b111;
											assign node2415 = (inp[11]) ? 3'b001 : 3'b101;
										assign node2418 = (inp[8]) ? 3'b101 : 3'b001;
									assign node2421 = (inp[8]) ? node2429 : node2422;
										assign node2422 = (inp[5]) ? 3'b110 : node2423;
											assign node2423 = (inp[2]) ? 3'b001 : node2424;
												assign node2424 = (inp[11]) ? 3'b001 : 3'b101;
										assign node2429 = (inp[5]) ? 3'b001 : 3'b101;
								assign node2432 = (inp[8]) ? node2446 : node2433;
									assign node2433 = (inp[5]) ? node2435 : 3'b110;
										assign node2435 = (inp[1]) ? node2441 : node2436;
											assign node2436 = (inp[11]) ? 3'b110 : node2437;
												assign node2437 = (inp[2]) ? 3'b110 : 3'b010;
											assign node2441 = (inp[2]) ? 3'b010 : node2442;
												assign node2442 = (inp[11]) ? 3'b010 : 3'b110;
									assign node2446 = (inp[11]) ? node2458 : node2447;
										assign node2447 = (inp[2]) ? node2453 : node2448;
											assign node2448 = (inp[5]) ? 3'b001 : node2449;
												assign node2449 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2453 = (inp[1]) ? node2455 : 3'b001;
												assign node2455 = (inp[5]) ? 3'b110 : 3'b001;
										assign node2458 = (inp[1]) ? node2464 : node2459;
											assign node2459 = (inp[5]) ? 3'b110 : node2460;
												assign node2460 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2464 = (inp[2]) ? 3'b110 : node2465;
												assign node2465 = (inp[5]) ? 3'b110 : 3'b010;
							assign node2469 = (inp[10]) ? node2505 : node2470;
								assign node2470 = (inp[11]) ? node2486 : node2471;
									assign node2471 = (inp[2]) ? 3'b110 : node2472;
										assign node2472 = (inp[8]) ? node2478 : node2473;
											assign node2473 = (inp[5]) ? 3'b010 : node2474;
												assign node2474 = (inp[1]) ? 3'b111 : 3'b110;
											assign node2478 = (inp[5]) ? node2482 : node2479;
												assign node2479 = (inp[1]) ? 3'b001 : 3'b101;
												assign node2482 = (inp[1]) ? 3'b110 : 3'b001;
									assign node2486 = (inp[5]) ? node2498 : node2487;
										assign node2487 = (inp[8]) ? node2495 : node2488;
											assign node2488 = (inp[1]) ? node2492 : node2489;
												assign node2489 = (inp[2]) ? 3'b110 : 3'b010;
												assign node2492 = (inp[2]) ? 3'b010 : 3'b100;
											assign node2495 = (inp[1]) ? 3'b110 : 3'b001;
										assign node2498 = (inp[8]) ? node2500 : 3'b010;
											assign node2500 = (inp[1]) ? node2502 : 3'b110;
												assign node2502 = (inp[2]) ? 3'b010 : 3'b110;
								assign node2505 = (inp[5]) ? node2519 : node2506;
									assign node2506 = (inp[8]) ? node2512 : node2507;
										assign node2507 = (inp[11]) ? node2509 : 3'b010;
											assign node2509 = (inp[1]) ? 3'b010 : 3'b000;
										assign node2512 = (inp[11]) ? 3'b110 : node2513;
											assign node2513 = (inp[2]) ? node2515 : 3'b001;
												assign node2515 = (inp[1]) ? 3'b010 : 3'b110;
									assign node2519 = (inp[8]) ? node2525 : node2520;
										assign node2520 = (inp[1]) ? 3'b100 : node2521;
											assign node2521 = (inp[2]) ? 3'b100 : 3'b000;
										assign node2525 = (inp[1]) ? node2527 : 3'b010;
											assign node2527 = (inp[11]) ? 3'b100 : 3'b010;
				assign node2530 = (inp[0]) ? node2788 : node2531;
					assign node2531 = (inp[1]) ? node2649 : node2532;
						assign node2532 = (inp[7]) ? node2602 : node2533;
							assign node2533 = (inp[11]) ? node2575 : node2534;
								assign node2534 = (inp[8]) ? node2554 : node2535;
									assign node2535 = (inp[2]) ? node2547 : node2536;
										assign node2536 = (inp[4]) ? node2542 : node2537;
											assign node2537 = (inp[10]) ? node2539 : 3'b110;
												assign node2539 = (inp[5]) ? 3'b010 : 3'b110;
											assign node2542 = (inp[5]) ? node2544 : 3'b110;
												assign node2544 = (inp[10]) ? 3'b100 : 3'b110;
										assign node2547 = (inp[5]) ? node2551 : node2548;
											assign node2548 = (inp[10]) ? 3'b110 : 3'b010;
											assign node2551 = (inp[10]) ? 3'b010 : 3'b110;
									assign node2554 = (inp[4]) ? node2568 : node2555;
										assign node2555 = (inp[10]) ? node2563 : node2556;
											assign node2556 = (inp[5]) ? node2560 : node2557;
												assign node2557 = (inp[2]) ? 3'b000 : 3'b100;
												assign node2560 = (inp[2]) ? 3'b111 : 3'b001;
											assign node2563 = (inp[5]) ? 3'b110 : node2564;
												assign node2564 = (inp[2]) ? 3'b111 : 3'b011;
										assign node2568 = (inp[5]) ? node2572 : node2569;
											assign node2569 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2572 = (inp[10]) ? 3'b100 : 3'b010;
								assign node2575 = (inp[8]) ? node2585 : node2576;
									assign node2576 = (inp[4]) ? node2578 : 3'b010;
										assign node2578 = (inp[5]) ? node2582 : node2579;
											assign node2579 = (inp[10]) ? 3'b110 : 3'b010;
											assign node2582 = (inp[10]) ? 3'b000 : 3'b110;
									assign node2585 = (inp[10]) ? node2595 : node2586;
										assign node2586 = (inp[5]) ? node2592 : node2587;
											assign node2587 = (inp[4]) ? node2589 : 3'b001;
												assign node2589 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2592 = (inp[4]) ? 3'b010 : 3'b110;
										assign node2595 = (inp[5]) ? node2599 : node2596;
											assign node2596 = (inp[4]) ? 3'b010 : 3'b110;
											assign node2599 = (inp[4]) ? 3'b100 : 3'b010;
							assign node2602 = (inp[10]) ? node2624 : node2603;
								assign node2603 = (inp[11]) ? node2617 : node2604;
									assign node2604 = (inp[5]) ? node2610 : node2605;
										assign node2605 = (inp[4]) ? 3'b001 : node2606;
											assign node2606 = (inp[8]) ? 3'b011 : 3'b001;
										assign node2610 = (inp[4]) ? node2614 : node2611;
											assign node2611 = (inp[8]) ? 3'b101 : 3'b001;
											assign node2614 = (inp[8]) ? 3'b001 : 3'b110;
									assign node2617 = (inp[4]) ? node2619 : 3'b101;
										assign node2619 = (inp[8]) ? node2621 : 3'b110;
											assign node2621 = (inp[5]) ? 3'b110 : 3'b001;
								assign node2624 = (inp[4]) ? node2638 : node2625;
									assign node2625 = (inp[11]) ? node2633 : node2626;
										assign node2626 = (inp[8]) ? node2628 : 3'b110;
											assign node2628 = (inp[2]) ? 3'b011 : node2629;
												assign node2629 = (inp[5]) ? 3'b001 : 3'b101;
										assign node2633 = (inp[8]) ? node2635 : 3'b000;
											assign node2635 = (inp[2]) ? 3'b000 : 3'b001;
									assign node2638 = (inp[11]) ? node2644 : node2639;
										assign node2639 = (inp[2]) ? node2641 : 3'b110;
											assign node2641 = (inp[5]) ? 3'b010 : 3'b110;
										assign node2644 = (inp[8]) ? node2646 : 3'b010;
											assign node2646 = (inp[5]) ? 3'b010 : 3'b110;
						assign node2649 = (inp[7]) ? node2717 : node2650;
							assign node2650 = (inp[4]) ? node2688 : node2651;
								assign node2651 = (inp[8]) ? node2671 : node2652;
									assign node2652 = (inp[10]) ? node2662 : node2653;
										assign node2653 = (inp[2]) ? node2659 : node2654;
											assign node2654 = (inp[11]) ? node2656 : 3'b010;
												assign node2656 = (inp[5]) ? 3'b100 : 3'b110;
											assign node2659 = (inp[11]) ? 3'b010 : 3'b100;
										assign node2662 = (inp[11]) ? node2666 : node2663;
											assign node2663 = (inp[5]) ? 3'b100 : 3'b010;
											assign node2666 = (inp[5]) ? node2668 : 3'b100;
												assign node2668 = (inp[2]) ? 3'b000 : 3'b100;
									assign node2671 = (inp[10]) ? node2681 : node2672;
										assign node2672 = (inp[5]) ? node2678 : node2673;
											assign node2673 = (inp[11]) ? 3'b100 : node2674;
												assign node2674 = (inp[2]) ? 3'b100 : 3'b111;
											assign node2678 = (inp[11]) ? 3'b010 : 3'b000;
										assign node2681 = (inp[5]) ? node2685 : node2682;
											assign node2682 = (inp[11]) ? 3'b010 : 3'b000;
											assign node2685 = (inp[11]) ? 3'b100 : 3'b110;
								assign node2688 = (inp[11]) ? node2702 : node2689;
									assign node2689 = (inp[8]) ? node2695 : node2690;
										assign node2690 = (inp[5]) ? 3'b000 : node2691;
											assign node2691 = (inp[10]) ? 3'b000 : 3'b100;
										assign node2695 = (inp[5]) ? node2699 : node2696;
											assign node2696 = (inp[10]) ? 3'b100 : 3'b000;
											assign node2699 = (inp[10]) ? 3'b000 : 3'b100;
									assign node2702 = (inp[8]) ? node2704 : 3'b000;
										assign node2704 = (inp[2]) ? node2712 : node2705;
											assign node2705 = (inp[10]) ? node2709 : node2706;
												assign node2706 = (inp[5]) ? 3'b100 : 3'b000;
												assign node2709 = (inp[5]) ? 3'b000 : 3'b100;
											assign node2712 = (inp[5]) ? 3'b000 : node2713;
												assign node2713 = (inp[10]) ? 3'b000 : 3'b100;
							assign node2717 = (inp[4]) ? node2753 : node2718;
								assign node2718 = (inp[11]) ? node2734 : node2719;
									assign node2719 = (inp[5]) ? node2725 : node2720;
										assign node2720 = (inp[10]) ? 3'b001 : node2721;
											assign node2721 = (inp[8]) ? 3'b101 : 3'b001;
										assign node2725 = (inp[8]) ? node2731 : node2726;
											assign node2726 = (inp[10]) ? node2728 : 3'b110;
												assign node2728 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2731 = (inp[10]) ? 3'b110 : 3'b001;
									assign node2734 = (inp[8]) ? node2742 : node2735;
										assign node2735 = (inp[5]) ? 3'b110 : node2736;
											assign node2736 = (inp[2]) ? node2738 : 3'b010;
												assign node2738 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2742 = (inp[2]) ? node2748 : node2743;
											assign node2743 = (inp[10]) ? node2745 : 3'b001;
												assign node2745 = (inp[5]) ? 3'b110 : 3'b001;
											assign node2748 = (inp[5]) ? 3'b110 : node2749;
												assign node2749 = (inp[10]) ? 3'b110 : 3'b001;
								assign node2753 = (inp[10]) ? node2771 : node2754;
									assign node2754 = (inp[11]) ? node2764 : node2755;
										assign node2755 = (inp[8]) ? node2759 : node2756;
											assign node2756 = (inp[2]) ? 3'b010 : 3'b011;
											assign node2759 = (inp[5]) ? node2761 : 3'b110;
												assign node2761 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2764 = (inp[8]) ? node2768 : node2765;
											assign node2765 = (inp[5]) ? 3'b100 : 3'b110;
											assign node2768 = (inp[5]) ? 3'b010 : 3'b110;
									assign node2771 = (inp[8]) ? node2779 : node2772;
										assign node2772 = (inp[11]) ? node2774 : 3'b100;
											assign node2774 = (inp[5]) ? node2776 : 3'b100;
												assign node2776 = (inp[2]) ? 3'b000 : 3'b100;
										assign node2779 = (inp[5]) ? node2785 : node2780;
											assign node2780 = (inp[11]) ? 3'b010 : node2781;
												assign node2781 = (inp[2]) ? 3'b000 : 3'b110;
											assign node2785 = (inp[11]) ? 3'b100 : 3'b010;
					assign node2788 = (inp[4]) ? node2896 : node2789;
						assign node2789 = (inp[7]) ? node2835 : node2790;
							assign node2790 = (inp[10]) ? node2822 : node2791;
								assign node2791 = (inp[1]) ? node2811 : node2792;
									assign node2792 = (inp[8]) ? node2800 : node2793;
										assign node2793 = (inp[11]) ? node2797 : node2794;
											assign node2794 = (inp[2]) ? 3'b100 : 3'b110;
											assign node2797 = (inp[5]) ? 3'b000 : 3'b100;
										assign node2800 = (inp[5]) ? node2806 : node2801;
											assign node2801 = (inp[11]) ? 3'b010 : node2802;
												assign node2802 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2806 = (inp[11]) ? 3'b100 : node2807;
												assign node2807 = (inp[2]) ? 3'b100 : 3'b010;
									assign node2811 = (inp[11]) ? node2817 : node2812;
										assign node2812 = (inp[5]) ? node2814 : 3'b100;
											assign node2814 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2817 = (inp[2]) ? node2819 : 3'b000;
											assign node2819 = (inp[5]) ? 3'b000 : 3'b100;
								assign node2822 = (inp[1]) ? 3'b000 : node2823;
									assign node2823 = (inp[5]) ? node2829 : node2824;
										assign node2824 = (inp[11]) ? node2826 : 3'b100;
											assign node2826 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2829 = (inp[11]) ? 3'b000 : node2830;
											assign node2830 = (inp[8]) ? 3'b100 : 3'b000;
							assign node2835 = (inp[10]) ? node2875 : node2836;
								assign node2836 = (inp[2]) ? node2854 : node2837;
									assign node2837 = (inp[1]) ? node2845 : node2838;
										assign node2838 = (inp[5]) ? 3'b110 : node2839;
											assign node2839 = (inp[8]) ? 3'b001 : node2840;
												assign node2840 = (inp[11]) ? 3'b101 : 3'b010;
										assign node2845 = (inp[5]) ? node2851 : node2846;
											assign node2846 = (inp[11]) ? node2848 : 3'b110;
												assign node2848 = (inp[8]) ? 3'b110 : 3'b010;
											assign node2851 = (inp[8]) ? 3'b010 : 3'b100;
									assign node2854 = (inp[5]) ? node2866 : node2855;
										assign node2855 = (inp[1]) ? node2861 : node2856;
											assign node2856 = (inp[8]) ? node2858 : 3'b110;
												assign node2858 = (inp[11]) ? 3'b110 : 3'b001;
											assign node2861 = (inp[11]) ? 3'b010 : node2862;
												assign node2862 = (inp[8]) ? 3'b110 : 3'b010;
										assign node2866 = (inp[8]) ? node2870 : node2867;
											assign node2867 = (inp[1]) ? 3'b100 : 3'b010;
											assign node2870 = (inp[1]) ? 3'b010 : node2871;
												assign node2871 = (inp[11]) ? 3'b010 : 3'b110;
								assign node2875 = (inp[5]) ? node2887 : node2876;
									assign node2876 = (inp[1]) ? node2884 : node2877;
										assign node2877 = (inp[8]) ? node2879 : 3'b010;
											assign node2879 = (inp[11]) ? node2881 : 3'b110;
												assign node2881 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2884 = (inp[8]) ? 3'b010 : 3'b100;
									assign node2887 = (inp[1]) ? node2891 : node2888;
										assign node2888 = (inp[8]) ? 3'b010 : 3'b100;
										assign node2891 = (inp[8]) ? 3'b100 : node2892;
											assign node2892 = (inp[2]) ? 3'b000 : 3'b100;
						assign node2896 = (inp[7]) ? node2898 : 3'b000;
							assign node2898 = (inp[1]) ? node2924 : node2899;
								assign node2899 = (inp[5]) ? node2913 : node2900;
									assign node2900 = (inp[10]) ? node2906 : node2901;
										assign node2901 = (inp[11]) ? node2903 : 3'b010;
											assign node2903 = (inp[8]) ? 3'b010 : 3'b100;
										assign node2906 = (inp[11]) ? node2910 : node2907;
											assign node2907 = (inp[2]) ? 3'b100 : 3'b110;
											assign node2910 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2913 = (inp[8]) ? node2919 : node2914;
										assign node2914 = (inp[11]) ? 3'b000 : node2915;
											assign node2915 = (inp[10]) ? 3'b000 : 3'b100;
										assign node2919 = (inp[10]) ? node2921 : 3'b100;
											assign node2921 = (inp[11]) ? 3'b000 : 3'b100;
								assign node2924 = (inp[10]) ? 3'b000 : node2925;
									assign node2925 = (inp[11]) ? node2931 : node2926;
										assign node2926 = (inp[8]) ? 3'b100 : node2927;
											assign node2927 = (inp[2]) ? 3'b100 : 3'b000;
										assign node2931 = (inp[5]) ? 3'b000 : node2932;
											assign node2932 = (inp[2]) ? 3'b100 : 3'b000;

endmodule