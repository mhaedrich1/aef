module dtc_split66_bm7 (
	input  wire [12-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node11;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node35;
	wire [1-1:0] node37;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node53;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node69;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node84;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node96;
	wire [1-1:0] node97;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node107;
	wire [1-1:0] node108;
	wire [1-1:0] node112;
	wire [1-1:0] node114;
	wire [1-1:0] node117;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node133;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node158;
	wire [1-1:0] node162;
	wire [1-1:0] node164;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node174;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node187;
	wire [1-1:0] node189;
	wire [1-1:0] node193;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node216;
	wire [1-1:0] node218;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node247;
	wire [1-1:0] node250;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node257;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node264;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node272;
	wire [1-1:0] node273;
	wire [1-1:0] node276;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node285;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node295;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node300;
	wire [1-1:0] node302;
	wire [1-1:0] node305;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node314;
	wire [1-1:0] node316;
	wire [1-1:0] node318;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node324;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node329;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node337;
	wire [1-1:0] node341;
	wire [1-1:0] node342;
	wire [1-1:0] node346;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node352;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node369;
	wire [1-1:0] node371;
	wire [1-1:0] node374;
	wire [1-1:0] node375;
	wire [1-1:0] node377;
	wire [1-1:0] node380;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node390;
	wire [1-1:0] node391;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node403;
	wire [1-1:0] node404;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node418;
	wire [1-1:0] node421;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node431;
	wire [1-1:0] node433;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node443;
	wire [1-1:0] node445;
	wire [1-1:0] node447;
	wire [1-1:0] node448;
	wire [1-1:0] node452;
	wire [1-1:0] node454;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node467;
	wire [1-1:0] node470;
	wire [1-1:0] node472;
	wire [1-1:0] node475;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node481;
	wire [1-1:0] node483;
	wire [1-1:0] node485;
	wire [1-1:0] node488;
	wire [1-1:0] node489;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node507;
	wire [1-1:0] node508;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node516;
	wire [1-1:0] node520;
	wire [1-1:0] node521;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node527;
	wire [1-1:0] node528;
	wire [1-1:0] node532;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node538;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node545;
	wire [1-1:0] node548;
	wire [1-1:0] node550;
	wire [1-1:0] node553;
	wire [1-1:0] node555;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node564;
	wire [1-1:0] node565;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node568;
	wire [1-1:0] node573;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node578;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node584;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node592;
	wire [1-1:0] node594;
	wire [1-1:0] node597;
	wire [1-1:0] node598;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node605;
	wire [1-1:0] node608;
	wire [1-1:0] node609;
	wire [1-1:0] node611;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node622;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node631;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node638;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node645;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node658;
	wire [1-1:0] node663;
	wire [1-1:0] node664;
	wire [1-1:0] node665;
	wire [1-1:0] node666;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node674;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node683;
	wire [1-1:0] node686;
	wire [1-1:0] node688;
	wire [1-1:0] node691;
	wire [1-1:0] node692;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node701;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node718;
	wire [1-1:0] node723;
	wire [1-1:0] node724;
	wire [1-1:0] node725;
	wire [1-1:0] node728;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node735;
	wire [1-1:0] node738;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node754;
	wire [1-1:0] node756;
	wire [1-1:0] node759;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node763;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node767;
	wire [1-1:0] node771;
	wire [1-1:0] node772;
	wire [1-1:0] node774;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node782;
	wire [1-1:0] node784;
	wire [1-1:0] node785;
	wire [1-1:0] node788;
	wire [1-1:0] node790;
	wire [1-1:0] node793;
	wire [1-1:0] node794;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node806;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node818;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node827;
	wire [1-1:0] node829;
	wire [1-1:0] node832;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node841;
	wire [1-1:0] node844;
	wire [1-1:0] node846;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node851;
	wire [1-1:0] node852;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node864;
	wire [1-1:0] node866;
	wire [1-1:0] node867;
	wire [1-1:0] node868;
	wire [1-1:0] node872;
	wire [1-1:0] node874;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node882;
	wire [1-1:0] node885;
	wire [1-1:0] node886;
	wire [1-1:0] node887;
	wire [1-1:0] node891;
	wire [1-1:0] node894;
	wire [1-1:0] node895;
	wire [1-1:0] node897;
	wire [1-1:0] node900;
	wire [1-1:0] node902;
	wire [1-1:0] node904;
	wire [1-1:0] node907;
	wire [1-1:0] node908;
	wire [1-1:0] node909;
	wire [1-1:0] node911;
	wire [1-1:0] node915;
	wire [1-1:0] node916;
	wire [1-1:0] node917;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node926;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node933;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node949;
	wire [1-1:0] node951;
	wire [1-1:0] node954;
	wire [1-1:0] node955;
	wire [1-1:0] node956;
	wire [1-1:0] node960;
	wire [1-1:0] node961;
	wire [1-1:0] node963;
	wire [1-1:0] node966;
	wire [1-1:0] node968;
	wire [1-1:0] node970;
	wire [1-1:0] node973;
	wire [1-1:0] node974;
	wire [1-1:0] node975;
	wire [1-1:0] node977;
	wire [1-1:0] node978;
	wire [1-1:0] node979;
	wire [1-1:0] node984;
	wire [1-1:0] node985;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node993;
	wire [1-1:0] node994;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node999;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1006;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1011;
	wire [1-1:0] node1016;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1020;
	wire [1-1:0] node1022;
	wire [1-1:0] node1023;
	wire [1-1:0] node1026;
	wire [1-1:0] node1029;
	wire [1-1:0] node1030;
	wire [1-1:0] node1031;
	wire [1-1:0] node1034;
	wire [1-1:0] node1038;
	wire [1-1:0] node1039;
	wire [1-1:0] node1041;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1046;
	wire [1-1:0] node1050;
	wire [1-1:0] node1052;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1058;
	wire [1-1:0] node1059;
	wire [1-1:0] node1063;
	wire [1-1:0] node1064;
	wire [1-1:0] node1065;
	wire [1-1:0] node1069;
	wire [1-1:0] node1071;
	wire [1-1:0] node1074;
	wire [1-1:0] node1075;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1078;
	wire [1-1:0] node1080;
	wire [1-1:0] node1084;
	wire [1-1:0] node1085;
	wire [1-1:0] node1089;
	wire [1-1:0] node1090;
	wire [1-1:0] node1093;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1099;
	wire [1-1:0] node1102;
	wire [1-1:0] node1105;
	wire [1-1:0] node1107;
	wire [1-1:0] node1109;
	wire [1-1:0] node1113;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1116;
	wire [1-1:0] node1117;
	wire [1-1:0] node1118;
	wire [1-1:0] node1119;
	wire [1-1:0] node1121;
	wire [1-1:0] node1124;
	wire [1-1:0] node1127;
	wire [1-1:0] node1128;
	wire [1-1:0] node1129;
	wire [1-1:0] node1134;
	wire [1-1:0] node1135;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1154;
	wire [1-1:0] node1156;
	wire [1-1:0] node1159;
	wire [1-1:0] node1160;
	wire [1-1:0] node1161;
	wire [1-1:0] node1162;
	wire [1-1:0] node1164;
	wire [1-1:0] node1166;
	wire [1-1:0] node1169;
	wire [1-1:0] node1172;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1178;
	wire [1-1:0] node1181;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1188;
	wire [1-1:0] node1189;
	wire [1-1:0] node1190;
	wire [1-1:0] node1193;
	wire [1-1:0] node1196;
	wire [1-1:0] node1197;
	wire [1-1:0] node1200;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1205;
	wire [1-1:0] node1208;
	wire [1-1:0] node1212;
	wire [1-1:0] node1213;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1219;
	wire [1-1:0] node1222;
	wire [1-1:0] node1223;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1230;
	wire [1-1:0] node1233;
	wire [1-1:0] node1234;
	wire [1-1:0] node1235;
	wire [1-1:0] node1239;
	wire [1-1:0] node1240;
	wire [1-1:0] node1242;
	wire [1-1:0] node1246;
	wire [1-1:0] node1247;
	wire [1-1:0] node1248;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1260;
	wire [1-1:0] node1263;
	wire [1-1:0] node1264;
	wire [1-1:0] node1267;
	wire [1-1:0] node1268;
	wire [1-1:0] node1269;
	wire [1-1:0] node1274;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1278;
	wire [1-1:0] node1281;
	wire [1-1:0] node1282;
	wire [1-1:0] node1286;
	wire [1-1:0] node1288;
	wire [1-1:0] node1289;
	wire [1-1:0] node1292;
	wire [1-1:0] node1294;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1300;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1304;
	wire [1-1:0] node1307;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1313;
	wire [1-1:0] node1316;
	wire [1-1:0] node1318;
	wire [1-1:0] node1320;
	wire [1-1:0] node1323;
	wire [1-1:0] node1324;
	wire [1-1:0] node1325;
	wire [1-1:0] node1326;
	wire [1-1:0] node1330;
	wire [1-1:0] node1331;
	wire [1-1:0] node1332;
	wire [1-1:0] node1335;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1344;
	wire [1-1:0] node1346;
	wire [1-1:0] node1350;
	wire [1-1:0] node1351;
	wire [1-1:0] node1352;
	wire [1-1:0] node1353;
	wire [1-1:0] node1354;
	wire [1-1:0] node1357;
	wire [1-1:0] node1358;
	wire [1-1:0] node1362;
	wire [1-1:0] node1363;
	wire [1-1:0] node1367;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1374;
	wire [1-1:0] node1375;
	wire [1-1:0] node1376;
	wire [1-1:0] node1380;
	wire [1-1:0] node1381;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1388;
	wire [1-1:0] node1389;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1396;
	wire [1-1:0] node1397;
	wire [1-1:0] node1398;
	wire [1-1:0] node1399;
	wire [1-1:0] node1403;
	wire [1-1:0] node1405;
	wire [1-1:0] node1408;
	wire [1-1:0] node1410;
	wire [1-1:0] node1411;
	wire [1-1:0] node1415;
	wire [1-1:0] node1416;
	wire [1-1:0] node1417;
	wire [1-1:0] node1418;
	wire [1-1:0] node1424;
	wire [1-1:0] node1425;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1431;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1437;
	wire [1-1:0] node1440;
	wire [1-1:0] node1442;
	wire [1-1:0] node1445;
	wire [1-1:0] node1446;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1449;
	wire [1-1:0] node1451;
	wire [1-1:0] node1456;
	wire [1-1:0] node1457;
	wire [1-1:0] node1459;
	wire [1-1:0] node1462;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1468;
	wire [1-1:0] node1470;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1475;
	wire [1-1:0] node1478;
	wire [1-1:0] node1481;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1487;
	wire [1-1:0] node1490;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1493;
	wire [1-1:0] node1494;
	wire [1-1:0] node1495;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1499;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1506;
	wire [1-1:0] node1509;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1514;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1525;
	wire [1-1:0] node1526;
	wire [1-1:0] node1528;
	wire [1-1:0] node1531;
	wire [1-1:0] node1532;
	wire [1-1:0] node1536;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1551;
	wire [1-1:0] node1554;
	wire [1-1:0] node1556;
	wire [1-1:0] node1558;
	wire [1-1:0] node1561;
	wire [1-1:0] node1562;
	wire [1-1:0] node1563;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1570;
	wire [1-1:0] node1574;
	wire [1-1:0] node1575;
	wire [1-1:0] node1579;
	wire [1-1:0] node1580;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1586;
	wire [1-1:0] node1589;
	wire [1-1:0] node1590;
	wire [1-1:0] node1594;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1598;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1606;
	wire [1-1:0] node1607;
	wire [1-1:0] node1609;
	wire [1-1:0] node1610;
	wire [1-1:0] node1615;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1620;
	wire [1-1:0] node1621;
	wire [1-1:0] node1625;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1629;
	wire [1-1:0] node1633;
	wire [1-1:0] node1634;
	wire [1-1:0] node1638;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1641;
	wire [1-1:0] node1642;
	wire [1-1:0] node1644;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1651;
	wire [1-1:0] node1654;
	wire [1-1:0] node1655;
	wire [1-1:0] node1659;
	wire [1-1:0] node1661;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1668;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1674;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1681;
	wire [1-1:0] node1684;
	wire [1-1:0] node1685;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1692;
	wire [1-1:0] node1693;
	wire [1-1:0] node1694;
	wire [1-1:0] node1698;
	wire [1-1:0] node1699;
	wire [1-1:0] node1702;
	wire [1-1:0] node1704;
	wire [1-1:0] node1707;
	wire [1-1:0] node1708;
	wire [1-1:0] node1709;
	wire [1-1:0] node1711;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1722;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1725;
	wire [1-1:0] node1726;
	wire [1-1:0] node1727;
	wire [1-1:0] node1728;
	wire [1-1:0] node1733;
	wire [1-1:0] node1734;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1740;
	wire [1-1:0] node1744;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1754;
	wire [1-1:0] node1756;
	wire [1-1:0] node1757;
	wire [1-1:0] node1761;
	wire [1-1:0] node1763;
	wire [1-1:0] node1764;
	wire [1-1:0] node1767;
	wire [1-1:0] node1770;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1773;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1779;
	wire [1-1:0] node1783;
	wire [1-1:0] node1784;
	wire [1-1:0] node1788;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1791;
	wire [1-1:0] node1792;
	wire [1-1:0] node1798;
	wire [1-1:0] node1800;
	wire [1-1:0] node1801;
	wire [1-1:0] node1805;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1810;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1817;
	wire [1-1:0] node1818;
	wire [1-1:0] node1819;
	wire [1-1:0] node1820;
	wire [1-1:0] node1823;
	wire [1-1:0] node1824;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1831;
	wire [1-1:0] node1832;
	wire [1-1:0] node1837;
	wire [1-1:0] node1838;
	wire [1-1:0] node1840;
	wire [1-1:0] node1842;
	wire [1-1:0] node1846;
	wire [1-1:0] node1847;
	wire [1-1:0] node1848;
	wire [1-1:0] node1849;
	wire [1-1:0] node1850;
	wire [1-1:0] node1852;
	wire [1-1:0] node1855;
	wire [1-1:0] node1856;
	wire [1-1:0] node1858;
	wire [1-1:0] node1861;
	wire [1-1:0] node1864;
	wire [1-1:0] node1865;
	wire [1-1:0] node1867;
	wire [1-1:0] node1870;
	wire [1-1:0] node1872;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1879;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1888;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1893;
	wire [1-1:0] node1894;
	wire [1-1:0] node1900;
	wire [1-1:0] node1901;
	wire [1-1:0] node1902;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1907;
	wire [1-1:0] node1909;
	wire [1-1:0] node1913;
	wire [1-1:0] node1914;
	wire [1-1:0] node1916;
	wire [1-1:0] node1920;
	wire [1-1:0] node1922;
	wire [1-1:0] node1923;
	wire [1-1:0] node1925;
	wire [1-1:0] node1928;
	wire [1-1:0] node1930;
	wire [1-1:0] node1933;
	wire [1-1:0] node1934;
	wire [1-1:0] node1935;
	wire [1-1:0] node1936;
	wire [1-1:0] node1938;
	wire [1-1:0] node1941;
	wire [1-1:0] node1942;
	wire [1-1:0] node1944;
	wire [1-1:0] node1945;
	wire [1-1:0] node1947;
	wire [1-1:0] node1950;
	wire [1-1:0] node1952;
	wire [1-1:0] node1955;
	wire [1-1:0] node1957;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1962;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1965;
	wire [1-1:0] node1968;
	wire [1-1:0] node1972;
	wire [1-1:0] node1973;
	wire [1-1:0] node1977;
	wire [1-1:0] node1978;
	wire [1-1:0] node1979;
	wire [1-1:0] node1982;
	wire [1-1:0] node1985;
	wire [1-1:0] node1986;
	wire [1-1:0] node1990;
	wire [1-1:0] node1991;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1997;
	wire [1-1:0] node1999;
	wire [1-1:0] node2002;
	wire [1-1:0] node2003;
	wire [1-1:0] node2005;
	wire [1-1:0] node2008;
	wire [1-1:0] node2009;
	wire [1-1:0] node2010;
	wire [1-1:0] node2015;
	wire [1-1:0] node2016;
	wire [1-1:0] node2017;
	wire [1-1:0] node2018;
	wire [1-1:0] node2019;
	wire [1-1:0] node2020;
	wire [1-1:0] node2024;
	wire [1-1:0] node2026;
	wire [1-1:0] node2029;
	wire [1-1:0] node2030;
	wire [1-1:0] node2032;
	wire [1-1:0] node2034;
	wire [1-1:0] node2037;
	wire [1-1:0] node2039;
	wire [1-1:0] node2041;
	wire [1-1:0] node2044;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2047;
	wire [1-1:0] node2050;
	wire [1-1:0] node2052;
	wire [1-1:0] node2055;
	wire [1-1:0] node2058;
	wire [1-1:0] node2060;
	wire [1-1:0] node2062;
	wire [1-1:0] node2065;
	wire [1-1:0] node2066;
	wire [1-1:0] node2067;
	wire [1-1:0] node2068;
	wire [1-1:0] node2073;
	wire [1-1:0] node2074;
	wire [1-1:0] node2075;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2081;
	wire [1-1:0] node2082;
	wire [1-1:0] node2086;
	wire [1-1:0] node2087;
	wire [1-1:0] node2091;
	wire [1-1:0] node2092;
	wire [1-1:0] node2093;
	wire [1-1:0] node2094;
	wire [1-1:0] node2097;
	wire [1-1:0] node2101;
	wire [1-1:0] node2102;
	wire [1-1:0] node2106;
	wire [1-1:0] node2107;
	wire [1-1:0] node2108;
	wire [1-1:0] node2109;
	wire [1-1:0] node2110;
	wire [1-1:0] node2111;
	wire [1-1:0] node2112;
	wire [1-1:0] node2114;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2119;
	wire [1-1:0] node2124;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2127;
	wire [1-1:0] node2131;
	wire [1-1:0] node2132;
	wire [1-1:0] node2136;
	wire [1-1:0] node2137;
	wire [1-1:0] node2138;
	wire [1-1:0] node2142;
	wire [1-1:0] node2143;
	wire [1-1:0] node2147;
	wire [1-1:0] node2148;
	wire [1-1:0] node2149;
	wire [1-1:0] node2152;
	wire [1-1:0] node2153;
	wire [1-1:0] node2155;
	wire [1-1:0] node2158;
	wire [1-1:0] node2159;
	wire [1-1:0] node2161;
	wire [1-1:0] node2165;
	wire [1-1:0] node2166;
	wire [1-1:0] node2167;
	wire [1-1:0] node2168;
	wire [1-1:0] node2171;
	wire [1-1:0] node2173;
	wire [1-1:0] node2176;
	wire [1-1:0] node2178;
	wire [1-1:0] node2181;
	wire [1-1:0] node2183;
	wire [1-1:0] node2185;
	wire [1-1:0] node2188;
	wire [1-1:0] node2189;
	wire [1-1:0] node2190;
	wire [1-1:0] node2191;
	wire [1-1:0] node2192;
	wire [1-1:0] node2194;
	wire [1-1:0] node2197;
	wire [1-1:0] node2200;
	wire [1-1:0] node2201;
	wire [1-1:0] node2202;
	wire [1-1:0] node2207;
	wire [1-1:0] node2208;
	wire [1-1:0] node2209;
	wire [1-1:0] node2210;
	wire [1-1:0] node2213;
	wire [1-1:0] node2216;
	wire [1-1:0] node2218;
	wire [1-1:0] node2221;
	wire [1-1:0] node2222;
	wire [1-1:0] node2223;
	wire [1-1:0] node2224;
	wire [1-1:0] node2228;
	wire [1-1:0] node2231;
	wire [1-1:0] node2234;
	wire [1-1:0] node2235;
	wire [1-1:0] node2236;
	wire [1-1:0] node2238;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2244;
	wire [1-1:0] node2247;
	wire [1-1:0] node2249;
	wire [1-1:0] node2252;
	wire [1-1:0] node2253;
	wire [1-1:0] node2255;
	wire [1-1:0] node2256;
	wire [1-1:0] node2257;
	wire [1-1:0] node2260;
	wire [1-1:0] node2264;
	wire [1-1:0] node2265;
	wire [1-1:0] node2266;
	wire [1-1:0] node2269;
	wire [1-1:0] node2272;
	wire [1-1:0] node2273;
	wire [1-1:0] node2275;
	wire [1-1:0] node2278;
	wire [1-1:0] node2279;
	wire [1-1:0] node2283;
	wire [1-1:0] node2284;
	wire [1-1:0] node2285;
	wire [1-1:0] node2286;
	wire [1-1:0] node2287;
	wire [1-1:0] node2288;
	wire [1-1:0] node2290;
	wire [1-1:0] node2292;
	wire [1-1:0] node2295;
	wire [1-1:0] node2297;
	wire [1-1:0] node2299;
	wire [1-1:0] node2302;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2309;
	wire [1-1:0] node2310;
	wire [1-1:0] node2311;
	wire [1-1:0] node2312;
	wire [1-1:0] node2316;
	wire [1-1:0] node2318;
	wire [1-1:0] node2321;
	wire [1-1:0] node2322;
	wire [1-1:0] node2323;
	wire [1-1:0] node2327;
	wire [1-1:0] node2328;
	wire [1-1:0] node2331;
	wire [1-1:0] node2332;
	wire [1-1:0] node2336;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2339;
	wire [1-1:0] node2340;
	wire [1-1:0] node2341;
	wire [1-1:0] node2345;
	wire [1-1:0] node2346;
	wire [1-1:0] node2349;
	wire [1-1:0] node2353;
	wire [1-1:0] node2354;
	wire [1-1:0] node2355;
	wire [1-1:0] node2356;
	wire [1-1:0] node2359;
	wire [1-1:0] node2364;
	wire [1-1:0] node2365;
	wire [1-1:0] node2367;
	wire [1-1:0] node2368;
	wire [1-1:0] node2372;
	wire [1-1:0] node2373;
	wire [1-1:0] node2375;
	wire [1-1:0] node2378;
	wire [1-1:0] node2379;
	wire [1-1:0] node2383;
	wire [1-1:0] node2384;
	wire [1-1:0] node2385;
	wire [1-1:0] node2387;
	wire [1-1:0] node2388;
	wire [1-1:0] node2389;
	wire [1-1:0] node2393;
	wire [1-1:0] node2395;
	wire [1-1:0] node2396;
	wire [1-1:0] node2400;
	wire [1-1:0] node2401;
	wire [1-1:0] node2402;
	wire [1-1:0] node2404;
	wire [1-1:0] node2406;
	wire [1-1:0] node2409;
	wire [1-1:0] node2411;
	wire [1-1:0] node2414;
	wire [1-1:0] node2416;
	wire [1-1:0] node2419;
	wire [1-1:0] node2420;
	wire [1-1:0] node2422;
	wire [1-1:0] node2425;
	wire [1-1:0] node2426;
	wire [1-1:0] node2428;
	wire [1-1:0] node2430;
	wire [1-1:0] node2433;
	wire [1-1:0] node2434;
	wire [1-1:0] node2436;
	wire [1-1:0] node2438;
	wire [1-1:0] node2441;
	wire [1-1:0] node2443;
	wire [1-1:0] node2445;
	wire [1-1:0] node2448;
	wire [1-1:0] node2449;
	wire [1-1:0] node2450;
	wire [1-1:0] node2451;
	wire [1-1:0] node2452;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2455;
	wire [1-1:0] node2456;
	wire [1-1:0] node2459;
	wire [1-1:0] node2462;
	wire [1-1:0] node2463;
	wire [1-1:0] node2466;
	wire [1-1:0] node2469;
	wire [1-1:0] node2470;
	wire [1-1:0] node2474;
	wire [1-1:0] node2475;
	wire [1-1:0] node2476;
	wire [1-1:0] node2479;
	wire [1-1:0] node2482;
	wire [1-1:0] node2484;
	wire [1-1:0] node2486;
	wire [1-1:0] node2489;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2494;
	wire [1-1:0] node2498;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2501;
	wire [1-1:0] node2503;
	wire [1-1:0] node2506;
	wire [1-1:0] node2509;
	wire [1-1:0] node2510;
	wire [1-1:0] node2513;
	wire [1-1:0] node2515;
	wire [1-1:0] node2518;
	wire [1-1:0] node2519;
	wire [1-1:0] node2520;
	wire [1-1:0] node2524;
	wire [1-1:0] node2525;
	wire [1-1:0] node2526;
	wire [1-1:0] node2530;
	wire [1-1:0] node2531;
	wire [1-1:0] node2535;
	wire [1-1:0] node2536;
	wire [1-1:0] node2537;
	wire [1-1:0] node2538;
	wire [1-1:0] node2540;
	wire [1-1:0] node2541;
	wire [1-1:0] node2544;
	wire [1-1:0] node2547;
	wire [1-1:0] node2548;
	wire [1-1:0] node2550;
	wire [1-1:0] node2552;
	wire [1-1:0] node2555;
	wire [1-1:0] node2557;
	wire [1-1:0] node2560;
	wire [1-1:0] node2561;
	wire [1-1:0] node2562;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2567;
	wire [1-1:0] node2571;
	wire [1-1:0] node2572;
	wire [1-1:0] node2576;
	wire [1-1:0] node2578;
	wire [1-1:0] node2579;
	wire [1-1:0] node2583;
	wire [1-1:0] node2584;
	wire [1-1:0] node2585;
	wire [1-1:0] node2586;
	wire [1-1:0] node2588;
	wire [1-1:0] node2591;
	wire [1-1:0] node2593;
	wire [1-1:0] node2596;
	wire [1-1:0] node2598;
	wire [1-1:0] node2599;
	wire [1-1:0] node2603;
	wire [1-1:0] node2604;
	wire [1-1:0] node2605;
	wire [1-1:0] node2606;
	wire [1-1:0] node2607;
	wire [1-1:0] node2611;
	wire [1-1:0] node2614;
	wire [1-1:0] node2615;
	wire [1-1:0] node2617;
	wire [1-1:0] node2620;
	wire [1-1:0] node2621;
	wire [1-1:0] node2624;
	wire [1-1:0] node2627;
	wire [1-1:0] node2628;
	wire [1-1:0] node2630;
	wire [1-1:0] node2633;
	wire [1-1:0] node2634;
	wire [1-1:0] node2635;
	wire [1-1:0] node2638;
	wire [1-1:0] node2641;
	wire [1-1:0] node2642;
	wire [1-1:0] node2645;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2651;
	wire [1-1:0] node2652;
	wire [1-1:0] node2653;
	wire [1-1:0] node2654;
	wire [1-1:0] node2658;
	wire [1-1:0] node2659;
	wire [1-1:0] node2663;
	wire [1-1:0] node2664;
	wire [1-1:0] node2665;
	wire [1-1:0] node2669;
	wire [1-1:0] node2671;
	wire [1-1:0] node2672;
	wire [1-1:0] node2676;
	wire [1-1:0] node2677;
	wire [1-1:0] node2678;
	wire [1-1:0] node2679;
	wire [1-1:0] node2681;
	wire [1-1:0] node2684;
	wire [1-1:0] node2685;
	wire [1-1:0] node2689;
	wire [1-1:0] node2690;
	wire [1-1:0] node2694;
	wire [1-1:0] node2696;
	wire [1-1:0] node2697;
	wire [1-1:0] node2699;
	wire [1-1:0] node2703;
	wire [1-1:0] node2704;
	wire [1-1:0] node2705;
	wire [1-1:0] node2706;
	wire [1-1:0] node2707;
	wire [1-1:0] node2708;
	wire [1-1:0] node2711;
	wire [1-1:0] node2715;
	wire [1-1:0] node2716;
	wire [1-1:0] node2718;
	wire [1-1:0] node2722;
	wire [1-1:0] node2723;
	wire [1-1:0] node2725;
	wire [1-1:0] node2728;
	wire [1-1:0] node2731;
	wire [1-1:0] node2732;
	wire [1-1:0] node2733;
	wire [1-1:0] node2735;
	wire [1-1:0] node2738;
	wire [1-1:0] node2740;
	wire [1-1:0] node2741;
	wire [1-1:0] node2745;
	wire [1-1:0] node2746;
	wire [1-1:0] node2747;
	wire [1-1:0] node2749;
	wire [1-1:0] node2752;
	wire [1-1:0] node2755;
	wire [1-1:0] node2757;
	wire [1-1:0] node2758;
	wire [1-1:0] node2762;
	wire [1-1:0] node2763;
	wire [1-1:0] node2764;
	wire [1-1:0] node2765;
	wire [1-1:0] node2766;
	wire [1-1:0] node2768;
	wire [1-1:0] node2771;
	wire [1-1:0] node2773;
	wire [1-1:0] node2774;
	wire [1-1:0] node2778;
	wire [1-1:0] node2779;
	wire [1-1:0] node2783;
	wire [1-1:0] node2784;
	wire [1-1:0] node2786;
	wire [1-1:0] node2789;
	wire [1-1:0] node2791;
	wire [1-1:0] node2794;
	wire [1-1:0] node2795;
	wire [1-1:0] node2796;
	wire [1-1:0] node2797;
	wire [1-1:0] node2798;
	wire [1-1:0] node2799;
	wire [1-1:0] node2803;
	wire [1-1:0] node2807;
	wire [1-1:0] node2808;
	wire [1-1:0] node2809;
	wire [1-1:0] node2811;
	wire [1-1:0] node2815;
	wire [1-1:0] node2816;
	wire [1-1:0] node2820;
	wire [1-1:0] node2821;
	wire [1-1:0] node2822;
	wire [1-1:0] node2825;
	wire [1-1:0] node2826;
	wire [1-1:0] node2830;
	wire [1-1:0] node2832;
	wire [1-1:0] node2834;

	assign outp = (inp[9]) ? node1490 : node1;
		assign node1 = (inp[0]) ? node759 : node2;
			assign node2 = (inp[2]) ? node400 : node3;
				assign node3 = (inp[10]) ? node221 : node4;
					assign node4 = (inp[1]) ? node124 : node5;
						assign node5 = (inp[8]) ? node59 : node6;
							assign node6 = (inp[6]) ? node40 : node7;
								assign node7 = (inp[4]) ? node27 : node8;
									assign node8 = (inp[3]) ? node18 : node9;
										assign node9 = (inp[5]) ? node15 : node10;
											assign node10 = (inp[7]) ? 1'b1 : node11;
												assign node11 = (inp[11]) ? 1'b1 : 1'b0;
											assign node15 = (inp[11]) ? 1'b0 : 1'b1;
										assign node18 = (inp[11]) ? node22 : node19;
											assign node19 = (inp[7]) ? 1'b0 : 1'b1;
											assign node22 = (inp[5]) ? node24 : 1'b0;
												assign node24 = (inp[7]) ? 1'b1 : 1'b0;
									assign node27 = (inp[7]) ? node35 : node28;
										assign node28 = (inp[5]) ? 1'b1 : node29;
											assign node29 = (inp[3]) ? node31 : 1'b0;
												assign node31 = (inp[11]) ? 1'b0 : 1'b1;
										assign node35 = (inp[5]) ? node37 : 1'b1;
											assign node37 = (inp[11]) ? 1'b1 : 1'b0;
								assign node40 = (inp[5]) ? node46 : node41;
									assign node41 = (inp[4]) ? 1'b0 : node42;
										assign node42 = (inp[3]) ? 1'b1 : 1'b0;
									assign node46 = (inp[3]) ? node50 : node47;
										assign node47 = (inp[11]) ? 1'b1 : 1'b0;
										assign node50 = (inp[11]) ? node52 : 1'b1;
											assign node52 = (inp[4]) ? node56 : node53;
												assign node53 = (inp[7]) ? 1'b1 : 1'b0;
												assign node56 = (inp[7]) ? 1'b0 : 1'b1;
							assign node59 = (inp[3]) ? node87 : node60;
								assign node60 = (inp[7]) ? node76 : node61;
									assign node61 = (inp[5]) ? node69 : node62;
										assign node62 = (inp[4]) ? node64 : 1'b1;
											assign node64 = (inp[11]) ? 1'b0 : node65;
												assign node65 = (inp[6]) ? 1'b0 : 1'b1;
										assign node69 = (inp[6]) ? node71 : 1'b1;
											assign node71 = (inp[11]) ? node73 : 1'b1;
												assign node73 = (inp[4]) ? 1'b1 : 1'b0;
									assign node76 = (inp[5]) ? node78 : 1'b1;
										assign node78 = (inp[4]) ? node84 : node79;
											assign node79 = (inp[6]) ? 1'b1 : node80;
												assign node80 = (inp[11]) ? 1'b1 : 1'b0;
											assign node84 = (inp[11]) ? 1'b0 : 1'b1;
								assign node87 = (inp[4]) ? node105 : node88;
									assign node88 = (inp[6]) ? node96 : node89;
										assign node89 = (inp[7]) ? node91 : 1'b0;
											assign node91 = (inp[11]) ? 1'b0 : node92;
												assign node92 = (inp[5]) ? 1'b1 : 1'b0;
										assign node96 = (inp[5]) ? node100 : node97;
											assign node97 = (inp[11]) ? 1'b1 : 1'b0;
											assign node100 = (inp[7]) ? 1'b1 : node101;
												assign node101 = (inp[11]) ? 1'b0 : 1'b1;
									assign node105 = (inp[6]) ? node117 : node106;
										assign node106 = (inp[5]) ? node112 : node107;
											assign node107 = (inp[11]) ? 1'b1 : node108;
												assign node108 = (inp[7]) ? 1'b1 : 1'b0;
											assign node112 = (inp[7]) ? node114 : 1'b1;
												assign node114 = (inp[11]) ? 1'b0 : 1'b1;
										assign node117 = (inp[11]) ? node119 : 1'b0;
											assign node119 = (inp[5]) ? 1'b1 : node120;
												assign node120 = (inp[7]) ? 1'b1 : 1'b0;
						assign node124 = (inp[3]) ? node178 : node125;
							assign node125 = (inp[6]) ? node155 : node126;
								assign node126 = (inp[5]) ? node144 : node127;
									assign node127 = (inp[4]) ? node137 : node128;
										assign node128 = (inp[7]) ? 1'b1 : node129;
											assign node129 = (inp[11]) ? node133 : node130;
												assign node130 = (inp[8]) ? 1'b1 : 1'b0;
												assign node133 = (inp[8]) ? 1'b0 : 1'b1;
										assign node137 = (inp[7]) ? 1'b0 : node138;
											assign node138 = (inp[11]) ? node140 : 1'b0;
												assign node140 = (inp[8]) ? 1'b0 : 1'b1;
									assign node144 = (inp[4]) ? 1'b1 : node145;
										assign node145 = (inp[7]) ? node147 : 1'b0;
											assign node147 = (inp[8]) ? node151 : node148;
												assign node148 = (inp[11]) ? 1'b1 : 1'b0;
												assign node151 = (inp[11]) ? 1'b0 : 1'b1;
								assign node155 = (inp[8]) ? node167 : node156;
									assign node156 = (inp[5]) ? node162 : node157;
										assign node157 = (inp[4]) ? 1'b0 : node158;
											assign node158 = (inp[7]) ? 1'b1 : 1'b0;
										assign node162 = (inp[11]) ? node164 : 1'b1;
											assign node164 = (inp[7]) ? 1'b0 : 1'b1;
									assign node167 = (inp[11]) ? 1'b0 : node168;
										assign node168 = (inp[4]) ? node174 : node169;
											assign node169 = (inp[7]) ? 1'b0 : node170;
												assign node170 = (inp[5]) ? 1'b1 : 1'b0;
											assign node174 = (inp[5]) ? 1'b0 : 1'b1;
							assign node178 = (inp[7]) ? node200 : node179;
								assign node179 = (inp[6]) ? node193 : node180;
									assign node180 = (inp[5]) ? 1'b1 : node181;
										assign node181 = (inp[8]) ? node187 : node182;
											assign node182 = (inp[11]) ? 1'b1 : node183;
												assign node183 = (inp[4]) ? 1'b0 : 1'b1;
											assign node187 = (inp[4]) ? node189 : 1'b0;
												assign node189 = (inp[11]) ? 1'b0 : 1'b1;
									assign node193 = (inp[5]) ? node195 : 1'b1;
										assign node195 = (inp[4]) ? 1'b1 : node196;
											assign node196 = (inp[11]) ? 1'b0 : 1'b1;
								assign node200 = (inp[5]) ? node212 : node201;
									assign node201 = (inp[4]) ? node207 : node202;
										assign node202 = (inp[8]) ? node204 : 1'b1;
											assign node204 = (inp[6]) ? 1'b0 : 1'b1;
										assign node207 = (inp[8]) ? node209 : 1'b0;
											assign node209 = (inp[6]) ? 1'b1 : 1'b0;
									assign node212 = (inp[11]) ? node216 : node213;
										assign node213 = (inp[8]) ? 1'b0 : 1'b1;
										assign node216 = (inp[8]) ? node218 : 1'b0;
											assign node218 = (inp[4]) ? 1'b1 : 1'b0;
					assign node221 = (inp[5]) ? node321 : node222;
						assign node222 = (inp[7]) ? node268 : node223;
							assign node223 = (inp[8]) ? node243 : node224;
								assign node224 = (inp[3]) ? node232 : node225;
									assign node225 = (inp[6]) ? node227 : 1'b0;
										assign node227 = (inp[1]) ? 1'b1 : node228;
											assign node228 = (inp[4]) ? 1'b1 : 1'b0;
									assign node232 = (inp[6]) ? node238 : node233;
										assign node233 = (inp[4]) ? node235 : 1'b1;
											assign node235 = (inp[1]) ? 1'b0 : 1'b1;
										assign node238 = (inp[1]) ? 1'b0 : node239;
											assign node239 = (inp[4]) ? 1'b1 : 1'b0;
								assign node243 = (inp[11]) ? node253 : node244;
									assign node244 = (inp[3]) ? node250 : node245;
										assign node245 = (inp[6]) ? node247 : 1'b1;
											assign node247 = (inp[1]) ? 1'b0 : 1'b1;
										assign node250 = (inp[6]) ? 1'b1 : 1'b0;
									assign node253 = (inp[4]) ? 1'b0 : node254;
										assign node254 = (inp[1]) ? node260 : node255;
											assign node255 = (inp[3]) ? node257 : 1'b0;
												assign node257 = (inp[6]) ? 1'b0 : 1'b1;
											assign node260 = (inp[3]) ? node264 : node261;
												assign node261 = (inp[6]) ? 1'b1 : 1'b0;
												assign node264 = (inp[6]) ? 1'b0 : 1'b1;
							assign node268 = (inp[11]) ? node294 : node269;
								assign node269 = (inp[8]) ? node285 : node270;
									assign node270 = (inp[4]) ? node280 : node271;
										assign node271 = (inp[1]) ? 1'b0 : node272;
											assign node272 = (inp[3]) ? node276 : node273;
												assign node273 = (inp[6]) ? 1'b1 : 1'b0;
												assign node276 = (inp[6]) ? 1'b0 : 1'b1;
										assign node280 = (inp[6]) ? 1'b1 : node281;
											assign node281 = (inp[3]) ? 1'b0 : 1'b1;
									assign node285 = (inp[1]) ? node287 : 1'b0;
										assign node287 = (inp[6]) ? node291 : node288;
											assign node288 = (inp[4]) ? 1'b1 : 1'b0;
											assign node291 = (inp[4]) ? 1'b0 : 1'b1;
								assign node294 = (inp[8]) ? node308 : node295;
									assign node295 = (inp[4]) ? node305 : node296;
										assign node296 = (inp[3]) ? node300 : node297;
											assign node297 = (inp[1]) ? 1'b1 : 1'b0;
											assign node300 = (inp[1]) ? node302 : 1'b1;
												assign node302 = (inp[6]) ? 1'b1 : 1'b0;
										assign node305 = (inp[6]) ? 1'b0 : 1'b1;
									assign node308 = (inp[1]) ? node314 : node309;
										assign node309 = (inp[4]) ? 1'b1 : node310;
											assign node310 = (inp[3]) ? 1'b0 : 1'b1;
										assign node314 = (inp[3]) ? node316 : 1'b0;
											assign node316 = (inp[4]) ? node318 : 1'b1;
												assign node318 = (inp[6]) ? 1'b1 : 1'b0;
						assign node321 = (inp[7]) ? node355 : node322;
							assign node322 = (inp[4]) ? node346 : node323;
								assign node323 = (inp[8]) ? node333 : node324;
									assign node324 = (inp[6]) ? 1'b0 : node325;
										assign node325 = (inp[1]) ? node329 : node326;
											assign node326 = (inp[3]) ? 1'b0 : 1'b1;
											assign node329 = (inp[3]) ? 1'b1 : 1'b0;
									assign node333 = (inp[11]) ? node341 : node334;
										assign node334 = (inp[6]) ? 1'b1 : node335;
											assign node335 = (inp[1]) ? node337 : 1'b1;
												assign node337 = (inp[3]) ? 1'b1 : 1'b0;
										assign node341 = (inp[6]) ? 1'b0 : node342;
											assign node342 = (inp[1]) ? 1'b0 : 1'b1;
								assign node346 = (inp[8]) ? node348 : 1'b1;
									assign node348 = (inp[11]) ? node352 : node349;
										assign node349 = (inp[6]) ? 1'b0 : 1'b1;
										assign node352 = (inp[6]) ? 1'b1 : 1'b0;
							assign node355 = (inp[6]) ? node383 : node356;
								assign node356 = (inp[3]) ? node374 : node357;
									assign node357 = (inp[1]) ? node369 : node358;
										assign node358 = (inp[4]) ? node364 : node359;
											assign node359 = (inp[8]) ? 1'b0 : node360;
												assign node360 = (inp[11]) ? 1'b1 : 1'b0;
											assign node364 = (inp[11]) ? node366 : 1'b1;
												assign node366 = (inp[8]) ? 1'b1 : 1'b0;
										assign node369 = (inp[4]) ? node371 : 1'b1;
											assign node371 = (inp[8]) ? 1'b0 : 1'b1;
									assign node374 = (inp[8]) ? node380 : node375;
										assign node375 = (inp[1]) ? node377 : 1'b0;
											assign node377 = (inp[11]) ? 1'b1 : 1'b0;
										assign node380 = (inp[1]) ? 1'b0 : 1'b1;
								assign node383 = (inp[1]) ? node395 : node384;
									assign node384 = (inp[4]) ? node390 : node385;
										assign node385 = (inp[11]) ? 1'b1 : node386;
											assign node386 = (inp[8]) ? 1'b1 : 1'b0;
										assign node390 = (inp[8]) ? 1'b0 : node391;
											assign node391 = (inp[11]) ? 1'b0 : 1'b1;
									assign node395 = (inp[11]) ? 1'b0 : node396;
										assign node396 = (inp[8]) ? 1'b0 : 1'b1;
				assign node400 = (inp[10]) ? node562 : node401;
					assign node401 = (inp[3]) ? node463 : node402;
						assign node402 = (inp[11]) ? node436 : node403;
							assign node403 = (inp[5]) ? node413 : node404;
								assign node404 = (inp[8]) ? node406 : 1'b0;
									assign node406 = (inp[6]) ? node410 : node407;
										assign node407 = (inp[7]) ? 1'b0 : 1'b1;
										assign node410 = (inp[7]) ? 1'b1 : 1'b0;
								assign node413 = (inp[8]) ? node431 : node414;
									assign node414 = (inp[1]) ? node424 : node415;
										assign node415 = (inp[6]) ? node421 : node416;
											assign node416 = (inp[7]) ? node418 : 1'b0;
												assign node418 = (inp[4]) ? 1'b0 : 1'b1;
											assign node421 = (inp[7]) ? 1'b0 : 1'b1;
										assign node424 = (inp[7]) ? 1'b1 : node425;
											assign node425 = (inp[4]) ? 1'b1 : node426;
												assign node426 = (inp[6]) ? 1'b1 : 1'b0;
									assign node431 = (inp[6]) ? node433 : 1'b0;
										assign node433 = (inp[7]) ? 1'b0 : 1'b1;
							assign node436 = (inp[5]) ? node452 : node437;
								assign node437 = (inp[6]) ? node443 : node438;
									assign node438 = (inp[7]) ? 1'b0 : node439;
										assign node439 = (inp[8]) ? 1'b0 : 1'b1;
									assign node443 = (inp[7]) ? node445 : 1'b0;
										assign node445 = (inp[8]) ? node447 : 1'b0;
											assign node447 = (inp[1]) ? 1'b1 : node448;
												assign node448 = (inp[4]) ? 1'b0 : 1'b1;
								assign node452 = (inp[7]) ? node454 : 1'b0;
									assign node454 = (inp[8]) ? node460 : node455;
										assign node455 = (inp[1]) ? 1'b0 : node456;
											assign node456 = (inp[6]) ? 1'b1 : 1'b0;
										assign node460 = (inp[6]) ? 1'b0 : 1'b1;
						assign node463 = (inp[7]) ? node507 : node464;
							assign node464 = (inp[1]) ? node488 : node465;
								assign node465 = (inp[4]) ? node475 : node466;
									assign node466 = (inp[8]) ? node470 : node467;
										assign node467 = (inp[11]) ? 1'b0 : 1'b1;
										assign node470 = (inp[11]) ? node472 : 1'b0;
											assign node472 = (inp[5]) ? 1'b0 : 1'b1;
									assign node475 = (inp[11]) ? node481 : node476;
										assign node476 = (inp[6]) ? 1'b1 : node477;
											assign node477 = (inp[8]) ? 1'b0 : 1'b1;
										assign node481 = (inp[8]) ? node483 : 1'b0;
											assign node483 = (inp[6]) ? node485 : 1'b1;
												assign node485 = (inp[5]) ? 1'b0 : 1'b1;
								assign node488 = (inp[6]) ? node502 : node489;
									assign node489 = (inp[5]) ? 1'b0 : node490;
										assign node490 = (inp[8]) ? node496 : node491;
											assign node491 = (inp[4]) ? 1'b1 : node492;
												assign node492 = (inp[11]) ? 1'b0 : 1'b1;
											assign node496 = (inp[11]) ? node498 : 1'b0;
												assign node498 = (inp[4]) ? 1'b0 : 1'b1;
									assign node502 = (inp[11]) ? 1'b0 : node503;
										assign node503 = (inp[5]) ? 1'b1 : 1'b0;
							assign node507 = (inp[1]) ? node541 : node508;
								assign node508 = (inp[6]) ? node520 : node509;
									assign node509 = (inp[4]) ? 1'b0 : node510;
										assign node510 = (inp[5]) ? node512 : 1'b0;
											assign node512 = (inp[11]) ? node516 : node513;
												assign node513 = (inp[8]) ? 1'b0 : 1'b1;
												assign node516 = (inp[8]) ? 1'b1 : 1'b0;
									assign node520 = (inp[11]) ? node532 : node521;
										assign node521 = (inp[4]) ? node527 : node522;
											assign node522 = (inp[5]) ? 1'b1 : node523;
												assign node523 = (inp[8]) ? 1'b1 : 1'b0;
											assign node527 = (inp[8]) ? 1'b0 : node528;
												assign node528 = (inp[5]) ? 1'b0 : 1'b1;
										assign node532 = (inp[8]) ? node534 : 1'b0;
											assign node534 = (inp[5]) ? node538 : node535;
												assign node535 = (inp[4]) ? 1'b0 : 1'b1;
												assign node538 = (inp[4]) ? 1'b1 : 1'b0;
								assign node541 = (inp[4]) ? node553 : node542;
									assign node542 = (inp[8]) ? node548 : node543;
										assign node543 = (inp[5]) ? node545 : 1'b1;
											assign node545 = (inp[11]) ? 1'b1 : 1'b0;
										assign node548 = (inp[5]) ? node550 : 1'b0;
											assign node550 = (inp[6]) ? 1'b1 : 1'b0;
									assign node553 = (inp[6]) ? node555 : 1'b1;
										assign node555 = (inp[5]) ? node557 : 1'b0;
											assign node557 = (inp[11]) ? 1'b1 : node558;
												assign node558 = (inp[8]) ? 1'b1 : 1'b0;
					assign node562 = (inp[5]) ? node648 : node563;
						assign node563 = (inp[8]) ? node597 : node564;
							assign node564 = (inp[11]) ? node582 : node565;
								assign node565 = (inp[6]) ? node573 : node566;
									assign node566 = (inp[1]) ? 1'b0 : node567;
										assign node567 = (inp[7]) ? 1'b1 : node568;
											assign node568 = (inp[3]) ? 1'b1 : 1'b0;
									assign node573 = (inp[3]) ? node575 : 1'b1;
										assign node575 = (inp[7]) ? 1'b0 : node576;
											assign node576 = (inp[4]) ? node578 : 1'b1;
												assign node578 = (inp[1]) ? 1'b1 : 1'b0;
								assign node582 = (inp[3]) ? node592 : node583;
									assign node583 = (inp[4]) ? node587 : node584;
										assign node584 = (inp[7]) ? 1'b0 : 1'b1;
										assign node587 = (inp[7]) ? 1'b1 : node588;
											assign node588 = (inp[6]) ? 1'b1 : 1'b0;
									assign node592 = (inp[7]) ? node594 : 1'b1;
										assign node594 = (inp[6]) ? 1'b0 : 1'b1;
							assign node597 = (inp[3]) ? node615 : node598;
								assign node598 = (inp[6]) ? node602 : node599;
									assign node599 = (inp[11]) ? 1'b0 : 1'b1;
									assign node602 = (inp[11]) ? node608 : node603;
										assign node603 = (inp[7]) ? node605 : 1'b0;
											assign node605 = (inp[1]) ? 1'b0 : 1'b1;
										assign node608 = (inp[1]) ? 1'b1 : node609;
											assign node609 = (inp[4]) ? node611 : 1'b1;
												assign node611 = (inp[7]) ? 1'b0 : 1'b1;
								assign node615 = (inp[7]) ? node625 : node616;
									assign node616 = (inp[11]) ? node622 : node617;
										assign node617 = (inp[1]) ? 1'b0 : node618;
											assign node618 = (inp[6]) ? 1'b1 : 1'b0;
										assign node622 = (inp[4]) ? 1'b0 : 1'b1;
									assign node625 = (inp[4]) ? node641 : node626;
										assign node626 = (inp[11]) ? node634 : node627;
											assign node627 = (inp[6]) ? node631 : node628;
												assign node628 = (inp[1]) ? 1'b0 : 1'b1;
												assign node631 = (inp[1]) ? 1'b1 : 1'b0;
											assign node634 = (inp[1]) ? node638 : node635;
												assign node635 = (inp[6]) ? 1'b1 : 1'b0;
												assign node638 = (inp[6]) ? 1'b0 : 1'b1;
										assign node641 = (inp[11]) ? node645 : node642;
											assign node642 = (inp[1]) ? 1'b0 : 1'b1;
											assign node645 = (inp[1]) ? 1'b1 : 1'b0;
						assign node648 = (inp[8]) ? node696 : node649;
							assign node649 = (inp[7]) ? node663 : node650;
								assign node650 = (inp[6]) ? 1'b0 : node651;
									assign node651 = (inp[4]) ? node653 : 1'b0;
										assign node653 = (inp[11]) ? 1'b1 : node654;
											assign node654 = (inp[1]) ? node658 : node655;
												assign node655 = (inp[3]) ? 1'b1 : 1'b0;
												assign node658 = (inp[3]) ? 1'b0 : 1'b1;
								assign node663 = (inp[6]) ? node677 : node664;
									assign node664 = (inp[11]) ? node674 : node665;
										assign node665 = (inp[1]) ? node669 : node666;
											assign node666 = (inp[4]) ? 1'b1 : 1'b0;
											assign node669 = (inp[4]) ? 1'b0 : node670;
												assign node670 = (inp[3]) ? 1'b1 : 1'b0;
										assign node674 = (inp[1]) ? 1'b1 : 1'b0;
									assign node677 = (inp[4]) ? node691 : node678;
										assign node678 = (inp[3]) ? node686 : node679;
											assign node679 = (inp[1]) ? node683 : node680;
												assign node680 = (inp[11]) ? 1'b1 : 1'b0;
												assign node683 = (inp[11]) ? 1'b0 : 1'b1;
											assign node686 = (inp[1]) ? node688 : 1'b0;
												assign node688 = (inp[11]) ? 1'b1 : 1'b0;
										assign node691 = (inp[3]) ? 1'b0 : node692;
											assign node692 = (inp[11]) ? 1'b0 : 1'b1;
							assign node696 = (inp[4]) ? node732 : node697;
								assign node697 = (inp[1]) ? node715 : node698;
									assign node698 = (inp[7]) ? node710 : node699;
										assign node699 = (inp[3]) ? node705 : node700;
											assign node700 = (inp[11]) ? 1'b1 : node701;
												assign node701 = (inp[6]) ? 1'b1 : 1'b0;
											assign node705 = (inp[6]) ? 1'b0 : node706;
												assign node706 = (inp[11]) ? 1'b1 : 1'b0;
										assign node710 = (inp[3]) ? 1'b0 : node711;
											assign node711 = (inp[6]) ? 1'b1 : 1'b0;
									assign node715 = (inp[3]) ? node723 : node716;
										assign node716 = (inp[7]) ? 1'b0 : node717;
											assign node717 = (inp[11]) ? 1'b1 : node718;
												assign node718 = (inp[6]) ? 1'b1 : 1'b0;
										assign node723 = (inp[7]) ? 1'b1 : node724;
											assign node724 = (inp[6]) ? node728 : node725;
												assign node725 = (inp[11]) ? 1'b1 : 1'b0;
												assign node728 = (inp[11]) ? 1'b0 : 1'b1;
								assign node732 = (inp[1]) ? node746 : node733;
									assign node733 = (inp[7]) ? node741 : node734;
										assign node734 = (inp[11]) ? node738 : node735;
											assign node735 = (inp[6]) ? 1'b1 : 1'b0;
											assign node738 = (inp[3]) ? 1'b0 : 1'b1;
										assign node741 = (inp[3]) ? 1'b1 : node742;
											assign node742 = (inp[11]) ? 1'b1 : 1'b0;
									assign node746 = (inp[7]) ? node754 : node747;
										assign node747 = (inp[11]) ? node749 : 1'b1;
											assign node749 = (inp[6]) ? 1'b0 : node750;
												assign node750 = (inp[3]) ? 1'b1 : 1'b0;
										assign node754 = (inp[3]) ? node756 : 1'b0;
											assign node756 = (inp[6]) ? 1'b1 : 1'b0;
			assign node759 = (inp[8]) ? node1113 : node760;
				assign node760 = (inp[7]) ? node930 : node761;
					assign node761 = (inp[2]) ? node849 : node762;
						assign node762 = (inp[10]) ? node818 : node763;
							assign node763 = (inp[5]) ? node793 : node764;
								assign node764 = (inp[11]) ? node782 : node765;
									assign node765 = (inp[4]) ? node771 : node766;
										assign node766 = (inp[3]) ? 1'b0 : node767;
											assign node767 = (inp[6]) ? 1'b0 : 1'b1;
										assign node771 = (inp[1]) ? node777 : node772;
											assign node772 = (inp[3]) ? node774 : 1'b1;
												assign node774 = (inp[6]) ? 1'b0 : 1'b1;
											assign node777 = (inp[6]) ? 1'b1 : node778;
												assign node778 = (inp[3]) ? 1'b1 : 1'b0;
									assign node782 = (inp[1]) ? node784 : 1'b0;
										assign node784 = (inp[6]) ? node788 : node785;
											assign node785 = (inp[3]) ? 1'b0 : 1'b1;
											assign node788 = (inp[3]) ? node790 : 1'b0;
												assign node790 = (inp[4]) ? 1'b0 : 1'b1;
								assign node793 = (inp[11]) ? node809 : node794;
									assign node794 = (inp[6]) ? node800 : node795;
										assign node795 = (inp[3]) ? 1'b0 : node796;
											assign node796 = (inp[4]) ? 1'b0 : 1'b1;
										assign node800 = (inp[3]) ? node806 : node801;
											assign node801 = (inp[1]) ? 1'b0 : node802;
												assign node802 = (inp[4]) ? 1'b1 : 1'b0;
											assign node806 = (inp[1]) ? 1'b1 : 1'b0;
									assign node809 = (inp[6]) ? 1'b1 : node810;
										assign node810 = (inp[3]) ? 1'b0 : node811;
											assign node811 = (inp[1]) ? 1'b1 : node812;
												assign node812 = (inp[4]) ? 1'b0 : 1'b1;
							assign node818 = (inp[6]) ? node832 : node819;
								assign node819 = (inp[3]) ? node827 : node820;
									assign node820 = (inp[4]) ? node822 : 1'b1;
										assign node822 = (inp[1]) ? 1'b0 : node823;
											assign node823 = (inp[5]) ? 1'b0 : 1'b1;
									assign node827 = (inp[4]) ? node829 : 1'b0;
										assign node829 = (inp[5]) ? 1'b0 : 1'b1;
								assign node832 = (inp[1]) ? node838 : node833;
									assign node833 = (inp[3]) ? 1'b1 : node834;
										assign node834 = (inp[4]) ? 1'b0 : 1'b1;
									assign node838 = (inp[3]) ? node844 : node839;
										assign node839 = (inp[4]) ? node841 : 1'b1;
											assign node841 = (inp[5]) ? 1'b1 : 1'b0;
										assign node844 = (inp[4]) ? node846 : 1'b0;
											assign node846 = (inp[5]) ? 1'b0 : 1'b1;
						assign node849 = (inp[6]) ? node877 : node850;
							assign node850 = (inp[3]) ? node864 : node851;
								assign node851 = (inp[1]) ? node855 : node852;
									assign node852 = (inp[5]) ? 1'b0 : 1'b1;
									assign node855 = (inp[5]) ? 1'b1 : node856;
										assign node856 = (inp[4]) ? 1'b0 : node857;
											assign node857 = (inp[10]) ? 1'b1 : node858;
												assign node858 = (inp[11]) ? 1'b0 : 1'b1;
								assign node864 = (inp[11]) ? node866 : 1'b1;
									assign node866 = (inp[4]) ? node872 : node867;
										assign node867 = (inp[10]) ? 1'b1 : node868;
											assign node868 = (inp[5]) ? 1'b1 : 1'b0;
										assign node872 = (inp[10]) ? node874 : 1'b0;
											assign node874 = (inp[1]) ? 1'b0 : 1'b1;
							assign node877 = (inp[11]) ? node907 : node878;
								assign node878 = (inp[3]) ? node894 : node879;
									assign node879 = (inp[10]) ? node885 : node880;
										assign node880 = (inp[1]) ? node882 : 1'b1;
											assign node882 = (inp[4]) ? 1'b0 : 1'b1;
										assign node885 = (inp[4]) ? node891 : node886;
											assign node886 = (inp[1]) ? 1'b0 : node887;
												assign node887 = (inp[5]) ? 1'b1 : 1'b0;
											assign node891 = (inp[1]) ? 1'b1 : 1'b0;
									assign node894 = (inp[1]) ? node900 : node895;
										assign node895 = (inp[10]) ? node897 : 1'b0;
											assign node897 = (inp[5]) ? 1'b1 : 1'b0;
										assign node900 = (inp[10]) ? node902 : 1'b1;
											assign node902 = (inp[4]) ? node904 : 1'b0;
												assign node904 = (inp[5]) ? 1'b1 : 1'b0;
								assign node907 = (inp[1]) ? node915 : node908;
									assign node908 = (inp[3]) ? 1'b1 : node909;
										assign node909 = (inp[5]) ? node911 : 1'b1;
											assign node911 = (inp[4]) ? 1'b0 : 1'b1;
									assign node915 = (inp[4]) ? node921 : node916;
										assign node916 = (inp[5]) ? 1'b0 : node917;
											assign node917 = (inp[10]) ? 1'b1 : 1'b0;
										assign node921 = (inp[5]) ? 1'b1 : node922;
											assign node922 = (inp[10]) ? node926 : node923;
												assign node923 = (inp[3]) ? 1'b1 : 1'b0;
												assign node926 = (inp[3]) ? 1'b0 : 1'b1;
					assign node930 = (inp[11]) ? node1016 : node931;
						assign node931 = (inp[10]) ? node973 : node932;
							assign node932 = (inp[2]) ? node954 : node933;
								assign node933 = (inp[1]) ? node943 : node934;
									assign node934 = (inp[3]) ? 1'b1 : node935;
										assign node935 = (inp[6]) ? node937 : 1'b1;
											assign node937 = (inp[4]) ? 1'b1 : node938;
												assign node938 = (inp[5]) ? 1'b0 : 1'b1;
									assign node943 = (inp[5]) ? node949 : node944;
										assign node944 = (inp[6]) ? node946 : 1'b1;
											assign node946 = (inp[4]) ? 1'b0 : 1'b1;
										assign node949 = (inp[6]) ? node951 : 1'b0;
											assign node951 = (inp[4]) ? 1'b1 : 1'b0;
								assign node954 = (inp[3]) ? node960 : node955;
									assign node955 = (inp[1]) ? 1'b1 : node956;
										assign node956 = (inp[6]) ? 1'b1 : 1'b0;
									assign node960 = (inp[6]) ? node966 : node961;
										assign node961 = (inp[1]) ? node963 : 1'b1;
											assign node963 = (inp[4]) ? 1'b1 : 1'b0;
										assign node966 = (inp[5]) ? node968 : 1'b0;
											assign node968 = (inp[1]) ? node970 : 1'b0;
												assign node970 = (inp[4]) ? 1'b0 : 1'b1;
							assign node973 = (inp[4]) ? node993 : node974;
								assign node974 = (inp[3]) ? node984 : node975;
									assign node975 = (inp[2]) ? node977 : 1'b0;
										assign node977 = (inp[1]) ? 1'b0 : node978;
											assign node978 = (inp[6]) ? 1'b0 : node979;
												assign node979 = (inp[5]) ? 1'b0 : 1'b1;
									assign node984 = (inp[1]) ? node988 : node985;
										assign node985 = (inp[6]) ? 1'b1 : 1'b0;
										assign node988 = (inp[2]) ? 1'b1 : node989;
											assign node989 = (inp[6]) ? 1'b0 : 1'b1;
								assign node993 = (inp[2]) ? node1003 : node994;
									assign node994 = (inp[1]) ? 1'b1 : node995;
										assign node995 = (inp[5]) ? node999 : node996;
											assign node996 = (inp[3]) ? 1'b0 : 1'b1;
											assign node999 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1003 = (inp[3]) ? node1009 : node1004;
										assign node1004 = (inp[6]) ? node1006 : 1'b1;
											assign node1006 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1009 = (inp[1]) ? 1'b0 : node1010;
											assign node1010 = (inp[5]) ? 1'b1 : node1011;
												assign node1011 = (inp[6]) ? 1'b1 : 1'b0;
						assign node1016 = (inp[4]) ? node1074 : node1017;
							assign node1017 = (inp[10]) ? node1055 : node1018;
								assign node1018 = (inp[5]) ? node1038 : node1019;
									assign node1019 = (inp[1]) ? node1029 : node1020;
										assign node1020 = (inp[2]) ? node1022 : 1'b1;
											assign node1022 = (inp[3]) ? node1026 : node1023;
												assign node1023 = (inp[6]) ? 1'b1 : 1'b0;
												assign node1026 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1029 = (inp[3]) ? 1'b0 : node1030;
											assign node1030 = (inp[2]) ? node1034 : node1031;
												assign node1031 = (inp[6]) ? 1'b1 : 1'b0;
												assign node1034 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1038 = (inp[6]) ? node1044 : node1039;
										assign node1039 = (inp[1]) ? node1041 : 1'b0;
											assign node1041 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1044 = (inp[2]) ? node1050 : node1045;
											assign node1045 = (inp[1]) ? 1'b1 : node1046;
												assign node1046 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1050 = (inp[3]) ? node1052 : 1'b0;
												assign node1052 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1055 = (inp[3]) ? node1063 : node1056;
									assign node1056 = (inp[2]) ? node1058 : 1'b1;
										assign node1058 = (inp[5]) ? 1'b1 : node1059;
											assign node1059 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1063 = (inp[1]) ? node1069 : node1064;
										assign node1064 = (inp[6]) ? 1'b0 : node1065;
											assign node1065 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1069 = (inp[5]) ? node1071 : 1'b1;
											assign node1071 = (inp[6]) ? 1'b1 : 1'b0;
							assign node1074 = (inp[6]) ? node1096 : node1075;
								assign node1075 = (inp[1]) ? node1089 : node1076;
									assign node1076 = (inp[10]) ? node1084 : node1077;
										assign node1077 = (inp[5]) ? 1'b1 : node1078;
											assign node1078 = (inp[3]) ? node1080 : 1'b0;
												assign node1080 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1084 = (inp[5]) ? 1'b0 : node1085;
											assign node1085 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1089 = (inp[2]) ? node1093 : node1090;
										assign node1090 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1093 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1096 = (inp[10]) ? 1'b0 : node1097;
									assign node1097 = (inp[5]) ? node1105 : node1098;
										assign node1098 = (inp[3]) ? node1102 : node1099;
											assign node1099 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1102 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1105 = (inp[1]) ? node1107 : 1'b0;
											assign node1107 = (inp[2]) ? node1109 : 1'b0;
												assign node1109 = (inp[3]) ? 1'b1 : 1'b0;
				assign node1113 = (inp[11]) ? node1297 : node1114;
					assign node1114 = (inp[1]) ? node1212 : node1115;
						assign node1115 = (inp[2]) ? node1159 : node1116;
							assign node1116 = (inp[7]) ? node1134 : node1117;
								assign node1117 = (inp[3]) ? node1127 : node1118;
									assign node1118 = (inp[4]) ? node1124 : node1119;
										assign node1119 = (inp[5]) ? node1121 : 1'b0;
											assign node1121 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1124 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1127 = (inp[6]) ? 1'b0 : node1128;
										assign node1128 = (inp[4]) ? 1'b0 : node1129;
											assign node1129 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1134 = (inp[3]) ? node1146 : node1135;
									assign node1135 = (inp[6]) ? node1141 : node1136;
										assign node1136 = (inp[5]) ? 1'b0 : node1137;
											assign node1137 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1141 = (inp[5]) ? 1'b1 : node1142;
											assign node1142 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1146 = (inp[6]) ? node1154 : node1147;
										assign node1147 = (inp[5]) ? 1'b1 : node1148;
											assign node1148 = (inp[4]) ? 1'b0 : node1149;
												assign node1149 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1154 = (inp[10]) ? node1156 : 1'b0;
											assign node1156 = (inp[5]) ? 1'b0 : 1'b1;
							assign node1159 = (inp[4]) ? node1181 : node1160;
								assign node1160 = (inp[5]) ? node1172 : node1161;
									assign node1161 = (inp[6]) ? node1169 : node1162;
										assign node1162 = (inp[7]) ? node1164 : 1'b0;
											assign node1164 = (inp[3]) ? node1166 : 1'b1;
												assign node1166 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1169 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1172 = (inp[3]) ? node1174 : 1'b0;
										assign node1174 = (inp[6]) ? node1178 : node1175;
											assign node1175 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1178 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1181 = (inp[5]) ? node1203 : node1182;
									assign node1182 = (inp[7]) ? node1188 : node1183;
										assign node1183 = (inp[3]) ? 1'b0 : node1184;
											assign node1184 = (inp[6]) ? 1'b1 : 1'b0;
										assign node1188 = (inp[6]) ? node1196 : node1189;
											assign node1189 = (inp[3]) ? node1193 : node1190;
												assign node1190 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1193 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1196 = (inp[10]) ? node1200 : node1197;
												assign node1197 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1200 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1203 = (inp[3]) ? 1'b1 : node1204;
										assign node1204 = (inp[7]) ? node1208 : node1205;
											assign node1205 = (inp[6]) ? 1'b1 : 1'b0;
											assign node1208 = (inp[6]) ? 1'b0 : 1'b1;
						assign node1212 = (inp[2]) ? node1246 : node1213;
							assign node1213 = (inp[4]) ? node1227 : node1214;
								assign node1214 = (inp[7]) ? node1222 : node1215;
									assign node1215 = (inp[3]) ? node1219 : node1216;
										assign node1216 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1219 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1222 = (inp[10]) ? 1'b1 : node1223;
										assign node1223 = (inp[5]) ? 1'b1 : 1'b0;
								assign node1227 = (inp[3]) ? node1233 : node1228;
									assign node1228 = (inp[5]) ? node1230 : 1'b1;
										assign node1230 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1233 = (inp[10]) ? node1239 : node1234;
										assign node1234 = (inp[7]) ? 1'b1 : node1235;
											assign node1235 = (inp[6]) ? 1'b1 : 1'b0;
										assign node1239 = (inp[6]) ? 1'b0 : node1240;
											assign node1240 = (inp[5]) ? node1242 : 1'b0;
												assign node1242 = (inp[7]) ? 1'b1 : 1'b0;
							assign node1246 = (inp[10]) ? node1274 : node1247;
								assign node1247 = (inp[7]) ? node1263 : node1248;
									assign node1248 = (inp[3]) ? node1254 : node1249;
										assign node1249 = (inp[5]) ? 1'b1 : node1250;
											assign node1250 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1254 = (inp[6]) ? node1260 : node1255;
											assign node1255 = (inp[4]) ? 1'b0 : node1256;
												assign node1256 = (inp[5]) ? 1'b1 : 1'b0;
											assign node1260 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1263 = (inp[3]) ? node1267 : node1264;
										assign node1264 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1267 = (inp[4]) ? 1'b1 : node1268;
											assign node1268 = (inp[6]) ? 1'b0 : node1269;
												assign node1269 = (inp[5]) ? 1'b1 : 1'b0;
								assign node1274 = (inp[6]) ? node1286 : node1275;
									assign node1275 = (inp[7]) ? node1281 : node1276;
										assign node1276 = (inp[5]) ? node1278 : 1'b0;
											assign node1278 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1281 = (inp[3]) ? 1'b1 : node1282;
											assign node1282 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1286 = (inp[3]) ? node1288 : 1'b0;
										assign node1288 = (inp[4]) ? node1292 : node1289;
											assign node1289 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1292 = (inp[7]) ? node1294 : 1'b0;
												assign node1294 = (inp[5]) ? 1'b1 : 1'b0;
					assign node1297 = (inp[3]) ? node1393 : node1298;
						assign node1298 = (inp[2]) ? node1350 : node1299;
							assign node1299 = (inp[5]) ? node1323 : node1300;
								assign node1300 = (inp[6]) ? node1316 : node1301;
									assign node1301 = (inp[4]) ? node1307 : node1302;
										assign node1302 = (inp[1]) ? node1304 : 1'b1;
											assign node1304 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1307 = (inp[10]) ? node1309 : 1'b0;
											assign node1309 = (inp[1]) ? node1313 : node1310;
												assign node1310 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1313 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1316 = (inp[4]) ? node1318 : 1'b0;
										assign node1318 = (inp[10]) ? node1320 : 1'b1;
											assign node1320 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1323 = (inp[1]) ? node1339 : node1324;
									assign node1324 = (inp[4]) ? node1330 : node1325;
										assign node1325 = (inp[6]) ? 1'b1 : node1326;
											assign node1326 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1330 = (inp[6]) ? 1'b0 : node1331;
											assign node1331 = (inp[7]) ? node1335 : node1332;
												assign node1332 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1335 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1339 = (inp[6]) ? 1'b1 : node1340;
										assign node1340 = (inp[4]) ? node1344 : node1341;
											assign node1341 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1344 = (inp[7]) ? node1346 : 1'b1;
												assign node1346 = (inp[10]) ? 1'b1 : 1'b0;
							assign node1350 = (inp[6]) ? node1374 : node1351;
								assign node1351 = (inp[10]) ? node1367 : node1352;
									assign node1352 = (inp[1]) ? node1362 : node1353;
										assign node1353 = (inp[4]) ? node1357 : node1354;
											assign node1354 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1357 = (inp[5]) ? 1'b0 : node1358;
												assign node1358 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1362 = (inp[7]) ? 1'b1 : node1363;
											assign node1363 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1367 = (inp[1]) ? 1'b0 : node1368;
										assign node1368 = (inp[4]) ? 1'b1 : node1369;
											assign node1369 = (inp[5]) ? 1'b1 : 1'b0;
								assign node1374 = (inp[1]) ? node1380 : node1375;
									assign node1375 = (inp[7]) ? 1'b0 : node1376;
										assign node1376 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1380 = (inp[7]) ? node1388 : node1381;
										assign node1381 = (inp[4]) ? node1383 : 1'b0;
											assign node1383 = (inp[10]) ? 1'b1 : node1384;
												assign node1384 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1388 = (inp[5]) ? 1'b0 : node1389;
											assign node1389 = (inp[4]) ? 1'b0 : 1'b1;
						assign node1393 = (inp[2]) ? node1445 : node1394;
							assign node1394 = (inp[10]) ? node1424 : node1395;
								assign node1395 = (inp[5]) ? node1415 : node1396;
									assign node1396 = (inp[6]) ? node1408 : node1397;
										assign node1397 = (inp[4]) ? node1403 : node1398;
											assign node1398 = (inp[1]) ? 1'b0 : node1399;
												assign node1399 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1403 = (inp[7]) ? node1405 : 1'b1;
												assign node1405 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1408 = (inp[1]) ? node1410 : 1'b0;
											assign node1410 = (inp[4]) ? 1'b0 : node1411;
												assign node1411 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1415 = (inp[4]) ? 1'b0 : node1416;
										assign node1416 = (inp[1]) ? 1'b0 : node1417;
											assign node1417 = (inp[7]) ? 1'b1 : node1418;
												assign node1418 = (inp[6]) ? 1'b1 : 1'b0;
								assign node1424 = (inp[4]) ? node1440 : node1425;
									assign node1425 = (inp[5]) ? node1431 : node1426;
										assign node1426 = (inp[7]) ? 1'b0 : node1427;
											assign node1427 = (inp[6]) ? 1'b1 : 1'b0;
										assign node1431 = (inp[6]) ? node1437 : node1432;
											assign node1432 = (inp[1]) ? 1'b1 : node1433;
												assign node1433 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1437 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1440 = (inp[6]) ? node1442 : 1'b1;
										assign node1442 = (inp[5]) ? 1'b0 : 1'b1;
							assign node1445 = (inp[5]) ? node1465 : node1446;
								assign node1446 = (inp[1]) ? node1456 : node1447;
									assign node1447 = (inp[7]) ? 1'b1 : node1448;
										assign node1448 = (inp[10]) ? 1'b1 : node1449;
											assign node1449 = (inp[4]) ? node1451 : 1'b1;
												assign node1451 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1456 = (inp[7]) ? node1462 : node1457;
										assign node1457 = (inp[10]) ? node1459 : 1'b1;
											assign node1459 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1462 = (inp[6]) ? 1'b1 : 1'b0;
								assign node1465 = (inp[7]) ? node1473 : node1466;
									assign node1466 = (inp[10]) ? node1468 : 1'b1;
										assign node1468 = (inp[1]) ? node1470 : 1'b0;
											assign node1470 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1473 = (inp[1]) ? node1481 : node1474;
										assign node1474 = (inp[4]) ? node1478 : node1475;
											assign node1475 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1478 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1481 = (inp[10]) ? node1483 : 1'b0;
											assign node1483 = (inp[4]) ? node1487 : node1484;
												assign node1484 = (inp[6]) ? 1'b0 : 1'b1;
												assign node1487 = (inp[6]) ? 1'b1 : 1'b0;
		assign node1490 = (inp[0]) ? node2106 : node1491;
			assign node1491 = (inp[11]) ? node1805 : node1492;
				assign node1492 = (inp[10]) ? node1638 : node1493;
					assign node1493 = (inp[5]) ? node1561 : node1494;
						assign node1494 = (inp[6]) ? node1518 : node1495;
							assign node1495 = (inp[3]) ? node1503 : node1496;
								assign node1496 = (inp[2]) ? 1'b0 : node1497;
									assign node1497 = (inp[7]) ? node1499 : 1'b0;
										assign node1499 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1503 = (inp[7]) ? node1509 : node1504;
									assign node1504 = (inp[4]) ? node1506 : 1'b1;
										assign node1506 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1509 = (inp[2]) ? 1'b0 : node1510;
										assign node1510 = (inp[1]) ? node1514 : node1511;
											assign node1511 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1514 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1518 = (inp[3]) ? node1536 : node1519;
								assign node1519 = (inp[7]) ? node1521 : 1'b1;
									assign node1521 = (inp[8]) ? node1525 : node1522;
										assign node1522 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1525 = (inp[1]) ? node1531 : node1526;
											assign node1526 = (inp[2]) ? node1528 : 1'b1;
												assign node1528 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1531 = (inp[2]) ? 1'b1 : node1532;
												assign node1532 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1536 = (inp[8]) ? node1546 : node1537;
									assign node1537 = (inp[7]) ? 1'b1 : node1538;
										assign node1538 = (inp[2]) ? 1'b1 : node1539;
											assign node1539 = (inp[1]) ? 1'b0 : node1540;
												assign node1540 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1546 = (inp[1]) ? node1554 : node1547;
										assign node1547 = (inp[2]) ? node1551 : node1548;
											assign node1548 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1551 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1554 = (inp[4]) ? node1556 : 1'b0;
											assign node1556 = (inp[7]) ? node1558 : 1'b0;
												assign node1558 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1561 = (inp[6]) ? node1615 : node1562;
							assign node1562 = (inp[8]) ? node1594 : node1563;
								assign node1563 = (inp[1]) ? node1579 : node1564;
									assign node1564 = (inp[4]) ? node1574 : node1565;
										assign node1565 = (inp[2]) ? 1'b1 : node1566;
											assign node1566 = (inp[3]) ? node1570 : node1567;
												assign node1567 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1570 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1574 = (inp[7]) ? 1'b0 : node1575;
											assign node1575 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1579 = (inp[4]) ? node1589 : node1580;
										assign node1580 = (inp[7]) ? node1582 : 1'b1;
											assign node1582 = (inp[2]) ? node1586 : node1583;
												assign node1583 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1586 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1589 = (inp[7]) ? 1'b1 : node1590;
											assign node1590 = (inp[3]) ? 1'b1 : 1'b0;
								assign node1594 = (inp[1]) ? node1606 : node1595;
									assign node1595 = (inp[4]) ? node1601 : node1596;
										assign node1596 = (inp[3]) ? node1598 : 1'b0;
											assign node1598 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1601 = (inp[7]) ? 1'b1 : node1602;
											assign node1602 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1606 = (inp[4]) ? 1'b0 : node1607;
										assign node1607 = (inp[2]) ? node1609 : 1'b0;
											assign node1609 = (inp[3]) ? 1'b1 : node1610;
												assign node1610 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1615 = (inp[2]) ? node1625 : node1616;
								assign node1616 = (inp[7]) ? node1620 : node1617;
									assign node1617 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1620 = (inp[4]) ? 1'b0 : node1621;
										assign node1621 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1625 = (inp[7]) ? node1627 : 1'b0;
									assign node1627 = (inp[3]) ? node1633 : node1628;
										assign node1628 = (inp[1]) ? 1'b0 : node1629;
											assign node1629 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1633 = (inp[1]) ? 1'b1 : node1634;
											assign node1634 = (inp[8]) ? 1'b0 : 1'b1;
					assign node1638 = (inp[5]) ? node1722 : node1639;
						assign node1639 = (inp[2]) ? node1689 : node1640;
							assign node1640 = (inp[3]) ? node1664 : node1641;
								assign node1641 = (inp[4]) ? node1647 : node1642;
									assign node1642 = (inp[1]) ? node1644 : 1'b1;
										assign node1644 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1647 = (inp[8]) ? node1659 : node1648;
										assign node1648 = (inp[1]) ? node1654 : node1649;
											assign node1649 = (inp[6]) ? node1651 : 1'b1;
												assign node1651 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1654 = (inp[6]) ? 1'b1 : node1655;
												assign node1655 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1659 = (inp[7]) ? node1661 : 1'b0;
											assign node1661 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1664 = (inp[4]) ? node1684 : node1665;
									assign node1665 = (inp[1]) ? node1671 : node1666;
										assign node1666 = (inp[8]) ? node1668 : 1'b0;
											assign node1668 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1671 = (inp[8]) ? node1677 : node1672;
											assign node1672 = (inp[6]) ? node1674 : 1'b1;
												assign node1674 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1677 = (inp[7]) ? node1681 : node1678;
												assign node1678 = (inp[6]) ? 1'b1 : 1'b0;
												assign node1681 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1684 = (inp[6]) ? 1'b1 : node1685;
										assign node1685 = (inp[1]) ? 1'b0 : 1'b1;
							assign node1689 = (inp[1]) ? node1707 : node1690;
								assign node1690 = (inp[6]) ? node1692 : 1'b0;
									assign node1692 = (inp[3]) ? node1698 : node1693;
										assign node1693 = (inp[4]) ? 1'b0 : node1694;
											assign node1694 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1698 = (inp[8]) ? node1702 : node1699;
											assign node1699 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1702 = (inp[7]) ? node1704 : 1'b1;
												assign node1704 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1707 = (inp[6]) ? node1717 : node1708;
									assign node1708 = (inp[7]) ? node1714 : node1709;
										assign node1709 = (inp[3]) ? node1711 : 1'b1;
											assign node1711 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1714 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1717 = (inp[3]) ? 1'b0 : node1718;
										assign node1718 = (inp[7]) ? 1'b1 : 1'b0;
						assign node1722 = (inp[1]) ? node1770 : node1723;
							assign node1723 = (inp[2]) ? node1747 : node1724;
								assign node1724 = (inp[7]) ? node1738 : node1725;
									assign node1725 = (inp[4]) ? node1733 : node1726;
										assign node1726 = (inp[6]) ? 1'b1 : node1727;
											assign node1727 = (inp[8]) ? 1'b0 : node1728;
												assign node1728 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1733 = (inp[6]) ? 1'b0 : node1734;
											assign node1734 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1738 = (inp[4]) ? node1744 : node1739;
										assign node1739 = (inp[6]) ? 1'b0 : node1740;
											assign node1740 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1744 = (inp[6]) ? 1'b1 : 1'b0;
								assign node1747 = (inp[6]) ? node1761 : node1748;
									assign node1748 = (inp[4]) ? node1754 : node1749;
										assign node1749 = (inp[8]) ? 1'b1 : node1750;
											assign node1750 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1754 = (inp[3]) ? node1756 : 1'b0;
											assign node1756 = (inp[8]) ? 1'b0 : node1757;
												assign node1757 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1761 = (inp[7]) ? node1763 : 1'b1;
										assign node1763 = (inp[3]) ? node1767 : node1764;
											assign node1764 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1767 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1770 = (inp[7]) ? node1788 : node1771;
								assign node1771 = (inp[4]) ? node1777 : node1772;
									assign node1772 = (inp[8]) ? 1'b1 : node1773;
										assign node1773 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1777 = (inp[2]) ? node1783 : node1778;
										assign node1778 = (inp[6]) ? 1'b0 : node1779;
											assign node1779 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1783 = (inp[6]) ? 1'b1 : node1784;
											assign node1784 = (inp[3]) ? 1'b1 : 1'b0;
								assign node1788 = (inp[2]) ? node1798 : node1789;
									assign node1789 = (inp[8]) ? 1'b1 : node1790;
										assign node1790 = (inp[3]) ? 1'b1 : node1791;
											assign node1791 = (inp[4]) ? 1'b1 : node1792;
												assign node1792 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1798 = (inp[3]) ? node1800 : 1'b1;
										assign node1800 = (inp[6]) ? 1'b0 : node1801;
											assign node1801 = (inp[4]) ? 1'b1 : 1'b0;
				assign node1805 = (inp[3]) ? node1933 : node1806;
					assign node1806 = (inp[7]) ? node1846 : node1807;
						assign node1807 = (inp[5]) ? node1817 : node1808;
							assign node1808 = (inp[6]) ? node1810 : 1'b1;
								assign node1810 = (inp[1]) ? 1'b1 : node1811;
									assign node1811 = (inp[4]) ? 1'b1 : node1812;
										assign node1812 = (inp[2]) ? 1'b1 : 1'b0;
							assign node1817 = (inp[4]) ? node1829 : node1818;
								assign node1818 = (inp[6]) ? 1'b1 : node1819;
									assign node1819 = (inp[10]) ? node1823 : node1820;
										assign node1820 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1823 = (inp[8]) ? 1'b1 : node1824;
											assign node1824 = (inp[2]) ? 1'b1 : 1'b0;
								assign node1829 = (inp[2]) ? node1837 : node1830;
									assign node1830 = (inp[10]) ? 1'b0 : node1831;
										assign node1831 = (inp[6]) ? 1'b0 : node1832;
											assign node1832 = (inp[8]) ? 1'b1 : 1'b0;
									assign node1837 = (inp[6]) ? 1'b1 : node1838;
										assign node1838 = (inp[1]) ? node1840 : 1'b1;
											assign node1840 = (inp[8]) ? node1842 : 1'b0;
												assign node1842 = (inp[10]) ? 1'b0 : 1'b1;
						assign node1846 = (inp[8]) ? node1900 : node1847;
							assign node1847 = (inp[1]) ? node1875 : node1848;
								assign node1848 = (inp[2]) ? node1864 : node1849;
									assign node1849 = (inp[10]) ? node1855 : node1850;
										assign node1850 = (inp[5]) ? node1852 : 1'b0;
											assign node1852 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1855 = (inp[4]) ? node1861 : node1856;
											assign node1856 = (inp[6]) ? node1858 : 1'b1;
												assign node1858 = (inp[5]) ? 1'b1 : 1'b0;
											assign node1861 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1864 = (inp[4]) ? node1870 : node1865;
										assign node1865 = (inp[5]) ? node1867 : 1'b0;
											assign node1867 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1870 = (inp[10]) ? node1872 : 1'b1;
											assign node1872 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1875 = (inp[6]) ? node1891 : node1876;
									assign node1876 = (inp[2]) ? node1884 : node1877;
										assign node1877 = (inp[5]) ? 1'b0 : node1878;
											assign node1878 = (inp[4]) ? 1'b0 : node1879;
												assign node1879 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1884 = (inp[5]) ? node1888 : node1885;
											assign node1885 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1888 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1891 = (inp[10]) ? 1'b0 : node1892;
										assign node1892 = (inp[5]) ? 1'b1 : node1893;
											assign node1893 = (inp[2]) ? 1'b0 : node1894;
												assign node1894 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1900 = (inp[2]) ? node1920 : node1901;
								assign node1901 = (inp[4]) ? node1913 : node1902;
									assign node1902 = (inp[1]) ? 1'b0 : node1903;
										assign node1903 = (inp[6]) ? node1907 : node1904;
											assign node1904 = (inp[5]) ? 1'b1 : 1'b0;
											assign node1907 = (inp[10]) ? node1909 : 1'b1;
												assign node1909 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1913 = (inp[1]) ? 1'b1 : node1914;
										assign node1914 = (inp[6]) ? node1916 : 1'b0;
											assign node1916 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1920 = (inp[5]) ? node1922 : 1'b1;
									assign node1922 = (inp[6]) ? node1928 : node1923;
										assign node1923 = (inp[4]) ? node1925 : 1'b1;
											assign node1925 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1928 = (inp[10]) ? node1930 : 1'b0;
											assign node1930 = (inp[1]) ? 1'b1 : 1'b0;
					assign node1933 = (inp[6]) ? node2015 : node1934;
						assign node1934 = (inp[7]) ? node1960 : node1935;
							assign node1935 = (inp[5]) ? node1941 : node1936;
								assign node1936 = (inp[1]) ? node1938 : 1'b0;
									assign node1938 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1941 = (inp[4]) ? node1955 : node1942;
									assign node1942 = (inp[1]) ? node1944 : 1'b1;
										assign node1944 = (inp[2]) ? node1950 : node1945;
											assign node1945 = (inp[8]) ? node1947 : 1'b0;
												assign node1947 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1950 = (inp[8]) ? node1952 : 1'b1;
												assign node1952 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1955 = (inp[1]) ? node1957 : 1'b0;
										assign node1957 = (inp[2]) ? 1'b1 : 1'b0;
							assign node1960 = (inp[2]) ? node1990 : node1961;
								assign node1961 = (inp[1]) ? node1977 : node1962;
									assign node1962 = (inp[8]) ? node1972 : node1963;
										assign node1963 = (inp[5]) ? 1'b1 : node1964;
											assign node1964 = (inp[10]) ? node1968 : node1965;
												assign node1965 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1968 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1972 = (inp[5]) ? 1'b0 : node1973;
											assign node1973 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1977 = (inp[8]) ? node1985 : node1978;
										assign node1978 = (inp[10]) ? node1982 : node1979;
											assign node1979 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1982 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1985 = (inp[5]) ? 1'b1 : node1986;
											assign node1986 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1990 = (inp[1]) ? node2002 : node1991;
									assign node1991 = (inp[8]) ? node1997 : node1992;
										assign node1992 = (inp[10]) ? 1'b0 : node1993;
											assign node1993 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1997 = (inp[5]) ? node1999 : 1'b1;
											assign node1999 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2002 = (inp[5]) ? node2008 : node2003;
										assign node2003 = (inp[10]) ? node2005 : 1'b0;
											assign node2005 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2008 = (inp[4]) ? 1'b1 : node2009;
											assign node2009 = (inp[8]) ? 1'b0 : node2010;
												assign node2010 = (inp[10]) ? 1'b0 : 1'b1;
						assign node2015 = (inp[2]) ? node2065 : node2016;
							assign node2016 = (inp[1]) ? node2044 : node2017;
								assign node2017 = (inp[5]) ? node2029 : node2018;
									assign node2018 = (inp[4]) ? node2024 : node2019;
										assign node2019 = (inp[8]) ? 1'b0 : node2020;
											assign node2020 = (inp[7]) ? 1'b1 : 1'b0;
										assign node2024 = (inp[7]) ? node2026 : 1'b1;
											assign node2026 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2029 = (inp[4]) ? node2037 : node2030;
										assign node2030 = (inp[10]) ? node2032 : 1'b1;
											assign node2032 = (inp[7]) ? node2034 : 1'b1;
												assign node2034 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2037 = (inp[7]) ? node2039 : 1'b0;
											assign node2039 = (inp[10]) ? node2041 : 1'b1;
												assign node2041 = (inp[8]) ? 1'b1 : 1'b0;
								assign node2044 = (inp[4]) ? node2058 : node2045;
									assign node2045 = (inp[8]) ? node2055 : node2046;
										assign node2046 = (inp[7]) ? node2050 : node2047;
											assign node2047 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2050 = (inp[5]) ? node2052 : 1'b1;
												assign node2052 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2055 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2058 = (inp[7]) ? node2060 : 1'b0;
										assign node2060 = (inp[8]) ? node2062 : 1'b0;
											assign node2062 = (inp[10]) ? 1'b1 : 1'b0;
							assign node2065 = (inp[7]) ? node2073 : node2066;
								assign node2066 = (inp[1]) ? 1'b1 : node2067;
									assign node2067 = (inp[5]) ? 1'b1 : node2068;
										assign node2068 = (inp[4]) ? 1'b0 : 1'b1;
								assign node2073 = (inp[8]) ? node2091 : node2074;
									assign node2074 = (inp[10]) ? node2086 : node2075;
										assign node2075 = (inp[5]) ? node2081 : node2076;
											assign node2076 = (inp[4]) ? 1'b1 : node2077;
												assign node2077 = (inp[1]) ? 1'b1 : 1'b0;
											assign node2081 = (inp[4]) ? 1'b0 : node2082;
												assign node2082 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2086 = (inp[1]) ? 1'b1 : node2087;
											assign node2087 = (inp[4]) ? 1'b1 : 1'b0;
									assign node2091 = (inp[10]) ? node2101 : node2092;
										assign node2092 = (inp[4]) ? 1'b1 : node2093;
											assign node2093 = (inp[5]) ? node2097 : node2094;
												assign node2094 = (inp[1]) ? 1'b0 : 1'b1;
												assign node2097 = (inp[1]) ? 1'b1 : 1'b0;
										assign node2101 = (inp[1]) ? 1'b0 : node2102;
											assign node2102 = (inp[4]) ? 1'b0 : 1'b1;
			assign node2106 = (inp[7]) ? node2448 : node2107;
				assign node2107 = (inp[2]) ? node2283 : node2108;
					assign node2108 = (inp[10]) ? node2188 : node2109;
						assign node2109 = (inp[1]) ? node2147 : node2110;
							assign node2110 = (inp[11]) ? node2124 : node2111;
								assign node2111 = (inp[3]) ? node2117 : node2112;
									assign node2112 = (inp[4]) ? node2114 : 1'b1;
										assign node2114 = (inp[6]) ? 1'b0 : 1'b1;
									assign node2117 = (inp[6]) ? 1'b1 : node2118;
										assign node2118 = (inp[5]) ? 1'b1 : node2119;
											assign node2119 = (inp[4]) ? 1'b1 : 1'b0;
								assign node2124 = (inp[6]) ? node2136 : node2125;
									assign node2125 = (inp[8]) ? node2131 : node2126;
										assign node2126 = (inp[5]) ? 1'b1 : node2127;
											assign node2127 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2131 = (inp[3]) ? 1'b0 : node2132;
											assign node2132 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2136 = (inp[5]) ? node2142 : node2137;
										assign node2137 = (inp[3]) ? 1'b1 : node2138;
											assign node2138 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2142 = (inp[3]) ? 1'b0 : node2143;
											assign node2143 = (inp[4]) ? 1'b1 : 1'b0;
							assign node2147 = (inp[3]) ? node2165 : node2148;
								assign node2148 = (inp[6]) ? node2152 : node2149;
									assign node2149 = (inp[4]) ? 1'b1 : 1'b0;
									assign node2152 = (inp[4]) ? node2158 : node2153;
										assign node2153 = (inp[5]) ? node2155 : 1'b1;
											assign node2155 = (inp[8]) ? 1'b1 : 1'b0;
										assign node2158 = (inp[8]) ? 1'b0 : node2159;
											assign node2159 = (inp[5]) ? node2161 : 1'b0;
												assign node2161 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2165 = (inp[4]) ? node2181 : node2166;
									assign node2166 = (inp[6]) ? node2176 : node2167;
										assign node2167 = (inp[5]) ? node2171 : node2168;
											assign node2168 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2171 = (inp[8]) ? node2173 : 1'b1;
												assign node2173 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2176 = (inp[5]) ? node2178 : 1'b0;
											assign node2178 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2181 = (inp[5]) ? node2183 : 1'b1;
										assign node2183 = (inp[6]) ? node2185 : 1'b1;
											assign node2185 = (inp[11]) ? 1'b1 : 1'b0;
						assign node2188 = (inp[11]) ? node2234 : node2189;
							assign node2189 = (inp[1]) ? node2207 : node2190;
								assign node2190 = (inp[3]) ? node2200 : node2191;
									assign node2191 = (inp[4]) ? node2197 : node2192;
										assign node2192 = (inp[5]) ? node2194 : 1'b0;
											assign node2194 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2197 = (inp[6]) ? 1'b1 : 1'b0;
									assign node2200 = (inp[6]) ? 1'b0 : node2201;
										assign node2201 = (inp[4]) ? 1'b0 : node2202;
											assign node2202 = (inp[5]) ? 1'b0 : 1'b1;
								assign node2207 = (inp[5]) ? node2221 : node2208;
									assign node2208 = (inp[8]) ? node2216 : node2209;
										assign node2209 = (inp[4]) ? node2213 : node2210;
											assign node2210 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2213 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2216 = (inp[4]) ? node2218 : 1'b1;
											assign node2218 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2221 = (inp[8]) ? node2231 : node2222;
										assign node2222 = (inp[4]) ? node2228 : node2223;
											assign node2223 = (inp[3]) ? 1'b1 : node2224;
												assign node2224 = (inp[6]) ? 1'b0 : 1'b1;
											assign node2228 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2231 = (inp[3]) ? 1'b1 : 1'b0;
							assign node2234 = (inp[3]) ? node2252 : node2235;
								assign node2235 = (inp[4]) ? node2241 : node2236;
									assign node2236 = (inp[6]) ? node2238 : 1'b0;
										assign node2238 = (inp[5]) ? 1'b0 : 1'b1;
									assign node2241 = (inp[6]) ? node2247 : node2242;
										assign node2242 = (inp[5]) ? node2244 : 1'b1;
											assign node2244 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2247 = (inp[5]) ? node2249 : 1'b0;
											assign node2249 = (inp[1]) ? 1'b0 : 1'b1;
								assign node2252 = (inp[4]) ? node2264 : node2253;
									assign node2253 = (inp[6]) ? node2255 : 1'b1;
										assign node2255 = (inp[8]) ? 1'b1 : node2256;
											assign node2256 = (inp[5]) ? node2260 : node2257;
												assign node2257 = (inp[1]) ? 1'b0 : 1'b1;
												assign node2260 = (inp[1]) ? 1'b1 : 1'b0;
									assign node2264 = (inp[8]) ? node2272 : node2265;
										assign node2265 = (inp[6]) ? node2269 : node2266;
											assign node2266 = (inp[5]) ? 1'b1 : 1'b0;
											assign node2269 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2272 = (inp[1]) ? node2278 : node2273;
											assign node2273 = (inp[6]) ? node2275 : 1'b0;
												assign node2275 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2278 = (inp[6]) ? 1'b1 : node2279;
												assign node2279 = (inp[5]) ? 1'b1 : 1'b0;
					assign node2283 = (inp[11]) ? node2383 : node2284;
						assign node2284 = (inp[8]) ? node2336 : node2285;
							assign node2285 = (inp[5]) ? node2309 : node2286;
								assign node2286 = (inp[1]) ? node2302 : node2287;
									assign node2287 = (inp[10]) ? node2295 : node2288;
										assign node2288 = (inp[6]) ? node2290 : 1'b1;
											assign node2290 = (inp[3]) ? node2292 : 1'b0;
												assign node2292 = (inp[4]) ? 1'b1 : 1'b0;
										assign node2295 = (inp[6]) ? node2297 : 1'b0;
											assign node2297 = (inp[3]) ? node2299 : 1'b1;
												assign node2299 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2302 = (inp[10]) ? node2304 : 1'b1;
										assign node2304 = (inp[3]) ? 1'b1 : node2305;
											assign node2305 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2309 = (inp[10]) ? node2321 : node2310;
									assign node2310 = (inp[4]) ? node2316 : node2311;
										assign node2311 = (inp[1]) ? 1'b0 : node2312;
											assign node2312 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2316 = (inp[3]) ? node2318 : 1'b0;
											assign node2318 = (inp[6]) ? 1'b1 : 1'b0;
									assign node2321 = (inp[6]) ? node2327 : node2322;
										assign node2322 = (inp[1]) ? 1'b1 : node2323;
											assign node2323 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2327 = (inp[4]) ? node2331 : node2328;
											assign node2328 = (inp[1]) ? 1'b1 : 1'b0;
											assign node2331 = (inp[3]) ? 1'b0 : node2332;
												assign node2332 = (inp[1]) ? 1'b0 : 1'b1;
							assign node2336 = (inp[1]) ? node2364 : node2337;
								assign node2337 = (inp[3]) ? node2353 : node2338;
									assign node2338 = (inp[5]) ? 1'b1 : node2339;
										assign node2339 = (inp[4]) ? node2345 : node2340;
											assign node2340 = (inp[10]) ? 1'b0 : node2341;
												assign node2341 = (inp[6]) ? 1'b0 : 1'b1;
											assign node2345 = (inp[6]) ? node2349 : node2346;
												assign node2346 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2349 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2353 = (inp[10]) ? 1'b0 : node2354;
										assign node2354 = (inp[4]) ? 1'b1 : node2355;
											assign node2355 = (inp[5]) ? node2359 : node2356;
												assign node2356 = (inp[6]) ? 1'b0 : 1'b1;
												assign node2359 = (inp[6]) ? 1'b1 : 1'b0;
								assign node2364 = (inp[6]) ? node2372 : node2365;
									assign node2365 = (inp[3]) ? node2367 : 1'b0;
										assign node2367 = (inp[5]) ? 1'b0 : node2368;
											assign node2368 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2372 = (inp[10]) ? node2378 : node2373;
										assign node2373 = (inp[4]) ? node2375 : 1'b0;
											assign node2375 = (inp[5]) ? 1'b1 : 1'b0;
										assign node2378 = (inp[3]) ? 1'b1 : node2379;
											assign node2379 = (inp[5]) ? 1'b1 : 1'b0;
						assign node2383 = (inp[3]) ? node2419 : node2384;
							assign node2384 = (inp[1]) ? node2400 : node2385;
								assign node2385 = (inp[5]) ? node2387 : 1'b0;
									assign node2387 = (inp[4]) ? node2393 : node2388;
										assign node2388 = (inp[6]) ? 1'b0 : node2389;
											assign node2389 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2393 = (inp[8]) ? node2395 : 1'b1;
											assign node2395 = (inp[6]) ? 1'b1 : node2396;
												assign node2396 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2400 = (inp[6]) ? node2414 : node2401;
									assign node2401 = (inp[4]) ? node2409 : node2402;
										assign node2402 = (inp[5]) ? node2404 : 1'b0;
											assign node2404 = (inp[8]) ? node2406 : 1'b0;
												assign node2406 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2409 = (inp[5]) ? node2411 : 1'b1;
											assign node2411 = (inp[8]) ? 1'b1 : 1'b0;
									assign node2414 = (inp[4]) ? node2416 : 1'b1;
										assign node2416 = (inp[5]) ? 1'b0 : 1'b1;
							assign node2419 = (inp[5]) ? node2425 : node2420;
								assign node2420 = (inp[6]) ? node2422 : 1'b0;
									assign node2422 = (inp[4]) ? 1'b1 : 1'b0;
								assign node2425 = (inp[8]) ? node2433 : node2426;
									assign node2426 = (inp[6]) ? node2428 : 1'b0;
										assign node2428 = (inp[1]) ? node2430 : 1'b0;
											assign node2430 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2433 = (inp[10]) ? node2441 : node2434;
										assign node2434 = (inp[6]) ? node2436 : 1'b1;
											assign node2436 = (inp[1]) ? node2438 : 1'b0;
												assign node2438 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2441 = (inp[6]) ? node2443 : 1'b0;
											assign node2443 = (inp[1]) ? node2445 : 1'b0;
												assign node2445 = (inp[4]) ? 1'b0 : 1'b1;
				assign node2448 = (inp[4]) ? node2648 : node2449;
					assign node2449 = (inp[3]) ? node2535 : node2450;
						assign node2450 = (inp[6]) ? node2498 : node2451;
							assign node2451 = (inp[5]) ? node2489 : node2452;
								assign node2452 = (inp[8]) ? node2474 : node2453;
									assign node2453 = (inp[10]) ? node2469 : node2454;
										assign node2454 = (inp[2]) ? node2462 : node2455;
											assign node2455 = (inp[1]) ? node2459 : node2456;
												assign node2456 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2459 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2462 = (inp[11]) ? node2466 : node2463;
												assign node2463 = (inp[1]) ? 1'b1 : 1'b0;
												assign node2466 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2469 = (inp[1]) ? 1'b0 : node2470;
											assign node2470 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2474 = (inp[1]) ? node2482 : node2475;
										assign node2475 = (inp[11]) ? node2479 : node2476;
											assign node2476 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2479 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2482 = (inp[10]) ? node2484 : 1'b1;
											assign node2484 = (inp[11]) ? node2486 : 1'b1;
												assign node2486 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2489 = (inp[10]) ? 1'b1 : node2490;
									assign node2490 = (inp[8]) ? node2494 : node2491;
										assign node2491 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2494 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2498 = (inp[10]) ? node2518 : node2499;
								assign node2499 = (inp[5]) ? node2509 : node2500;
									assign node2500 = (inp[8]) ? node2506 : node2501;
										assign node2501 = (inp[1]) ? node2503 : 1'b1;
											assign node2503 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2506 = (inp[2]) ? 1'b1 : 1'b0;
									assign node2509 = (inp[2]) ? node2513 : node2510;
										assign node2510 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2513 = (inp[11]) ? node2515 : 1'b0;
											assign node2515 = (inp[8]) ? 1'b0 : 1'b1;
								assign node2518 = (inp[2]) ? node2524 : node2519;
									assign node2519 = (inp[8]) ? 1'b0 : node2520;
										assign node2520 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2524 = (inp[8]) ? node2530 : node2525;
										assign node2525 = (inp[5]) ? 1'b0 : node2526;
											assign node2526 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2530 = (inp[1]) ? 1'b1 : node2531;
											assign node2531 = (inp[5]) ? 1'b1 : 1'b0;
						assign node2535 = (inp[1]) ? node2583 : node2536;
							assign node2536 = (inp[5]) ? node2560 : node2537;
								assign node2537 = (inp[11]) ? node2547 : node2538;
									assign node2538 = (inp[6]) ? node2540 : 1'b1;
										assign node2540 = (inp[2]) ? node2544 : node2541;
											assign node2541 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2544 = (inp[8]) ? 1'b1 : 1'b0;
									assign node2547 = (inp[8]) ? node2555 : node2548;
										assign node2548 = (inp[2]) ? node2550 : 1'b1;
											assign node2550 = (inp[10]) ? node2552 : 1'b0;
												assign node2552 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2555 = (inp[2]) ? node2557 : 1'b0;
											assign node2557 = (inp[6]) ? 1'b1 : 1'b0;
								assign node2560 = (inp[10]) ? node2576 : node2561;
									assign node2561 = (inp[2]) ? node2571 : node2562;
										assign node2562 = (inp[6]) ? 1'b0 : node2563;
											assign node2563 = (inp[8]) ? node2567 : node2564;
												assign node2564 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2567 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2571 = (inp[6]) ? 1'b1 : node2572;
											assign node2572 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2576 = (inp[6]) ? node2578 : 1'b1;
										assign node2578 = (inp[11]) ? 1'b1 : node2579;
											assign node2579 = (inp[8]) ? 1'b1 : 1'b0;
							assign node2583 = (inp[6]) ? node2603 : node2584;
								assign node2584 = (inp[10]) ? node2596 : node2585;
									assign node2585 = (inp[11]) ? node2591 : node2586;
										assign node2586 = (inp[8]) ? node2588 : 1'b0;
											assign node2588 = (inp[5]) ? 1'b1 : 1'b0;
										assign node2591 = (inp[8]) ? node2593 : 1'b1;
											assign node2593 = (inp[5]) ? 1'b0 : 1'b1;
									assign node2596 = (inp[8]) ? node2598 : 1'b0;
										assign node2598 = (inp[5]) ? 1'b0 : node2599;
											assign node2599 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2603 = (inp[11]) ? node2627 : node2604;
									assign node2604 = (inp[5]) ? node2614 : node2605;
										assign node2605 = (inp[10]) ? node2611 : node2606;
											assign node2606 = (inp[8]) ? 1'b1 : node2607;
												assign node2607 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2611 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2614 = (inp[8]) ? node2620 : node2615;
											assign node2615 = (inp[2]) ? node2617 : 1'b1;
												assign node2617 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2620 = (inp[2]) ? node2624 : node2621;
												assign node2621 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2624 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2627 = (inp[5]) ? node2633 : node2628;
										assign node2628 = (inp[2]) ? node2630 : 1'b0;
											assign node2630 = (inp[8]) ? 1'b1 : 1'b0;
										assign node2633 = (inp[10]) ? node2641 : node2634;
											assign node2634 = (inp[2]) ? node2638 : node2635;
												assign node2635 = (inp[8]) ? 1'b1 : 1'b0;
												assign node2638 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2641 = (inp[8]) ? node2645 : node2642;
												assign node2642 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2645 = (inp[2]) ? 1'b1 : 1'b0;
					assign node2648 = (inp[8]) ? node2762 : node2649;
						assign node2649 = (inp[3]) ? node2703 : node2650;
							assign node2650 = (inp[1]) ? node2676 : node2651;
								assign node2651 = (inp[6]) ? node2663 : node2652;
									assign node2652 = (inp[2]) ? node2658 : node2653;
										assign node2653 = (inp[5]) ? 1'b1 : node2654;
											assign node2654 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2658 = (inp[10]) ? 1'b0 : node2659;
											assign node2659 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2663 = (inp[2]) ? node2669 : node2664;
										assign node2664 = (inp[11]) ? 1'b0 : node2665;
											assign node2665 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2669 = (inp[5]) ? node2671 : 1'b1;
											assign node2671 = (inp[11]) ? 1'b0 : node2672;
												assign node2672 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2676 = (inp[11]) ? node2694 : node2677;
									assign node2677 = (inp[10]) ? node2689 : node2678;
										assign node2678 = (inp[6]) ? node2684 : node2679;
											assign node2679 = (inp[2]) ? node2681 : 1'b1;
												assign node2681 = (inp[5]) ? 1'b1 : 1'b0;
											assign node2684 = (inp[5]) ? 1'b0 : node2685;
												assign node2685 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2689 = (inp[5]) ? 1'b1 : node2690;
											assign node2690 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2694 = (inp[10]) ? node2696 : 1'b1;
										assign node2696 = (inp[5]) ? 1'b0 : node2697;
											assign node2697 = (inp[2]) ? node2699 : 1'b1;
												assign node2699 = (inp[6]) ? 1'b1 : 1'b0;
							assign node2703 = (inp[1]) ? node2731 : node2704;
								assign node2704 = (inp[5]) ? node2722 : node2705;
									assign node2705 = (inp[10]) ? node2715 : node2706;
										assign node2706 = (inp[6]) ? 1'b0 : node2707;
											assign node2707 = (inp[2]) ? node2711 : node2708;
												assign node2708 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2711 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2715 = (inp[2]) ? 1'b1 : node2716;
											assign node2716 = (inp[6]) ? node2718 : 1'b0;
												assign node2718 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2722 = (inp[6]) ? node2728 : node2723;
										assign node2723 = (inp[11]) ? node2725 : 1'b0;
											assign node2725 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2728 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2731 = (inp[5]) ? node2745 : node2732;
									assign node2732 = (inp[10]) ? node2738 : node2733;
										assign node2733 = (inp[2]) ? node2735 : 1'b0;
											assign node2735 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2738 = (inp[2]) ? node2740 : 1'b1;
											assign node2740 = (inp[11]) ? 1'b0 : node2741;
												assign node2741 = (inp[6]) ? 1'b1 : 1'b0;
									assign node2745 = (inp[11]) ? node2755 : node2746;
										assign node2746 = (inp[2]) ? node2752 : node2747;
											assign node2747 = (inp[10]) ? node2749 : 1'b0;
												assign node2749 = (inp[6]) ? 1'b1 : 1'b0;
											assign node2752 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2755 = (inp[6]) ? node2757 : 1'b0;
											assign node2757 = (inp[2]) ? 1'b0 : node2758;
												assign node2758 = (inp[10]) ? 1'b0 : 1'b1;
						assign node2762 = (inp[10]) ? node2794 : node2763;
							assign node2763 = (inp[3]) ? node2783 : node2764;
								assign node2764 = (inp[1]) ? node2778 : node2765;
									assign node2765 = (inp[11]) ? node2771 : node2766;
										assign node2766 = (inp[2]) ? node2768 : 1'b0;
											assign node2768 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2771 = (inp[6]) ? node2773 : 1'b1;
											assign node2773 = (inp[2]) ? 1'b0 : node2774;
												assign node2774 = (inp[5]) ? 1'b0 : 1'b1;
									assign node2778 = (inp[5]) ? 1'b0 : node2779;
										assign node2779 = (inp[6]) ? 1'b1 : 1'b0;
								assign node2783 = (inp[11]) ? node2789 : node2784;
									assign node2784 = (inp[2]) ? node2786 : 1'b1;
										assign node2786 = (inp[1]) ? 1'b0 : 1'b1;
									assign node2789 = (inp[2]) ? node2791 : 1'b0;
										assign node2791 = (inp[1]) ? 1'b1 : 1'b0;
							assign node2794 = (inp[6]) ? node2820 : node2795;
								assign node2795 = (inp[2]) ? node2807 : node2796;
									assign node2796 = (inp[1]) ? 1'b0 : node2797;
										assign node2797 = (inp[11]) ? node2803 : node2798;
											assign node2798 = (inp[3]) ? 1'b0 : node2799;
												assign node2799 = (inp[5]) ? 1'b1 : 1'b0;
											assign node2803 = (inp[5]) ? 1'b0 : 1'b1;
									assign node2807 = (inp[1]) ? node2815 : node2808;
										assign node2808 = (inp[5]) ? 1'b0 : node2809;
											assign node2809 = (inp[3]) ? node2811 : 1'b0;
												assign node2811 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2815 = (inp[5]) ? 1'b1 : node2816;
											assign node2816 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2820 = (inp[5]) ? node2830 : node2821;
									assign node2821 = (inp[11]) ? node2825 : node2822;
										assign node2822 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2825 = (inp[1]) ? 1'b1 : node2826;
											assign node2826 = (inp[2]) ? 1'b1 : 1'b0;
									assign node2830 = (inp[2]) ? node2832 : 1'b1;
										assign node2832 = (inp[1]) ? node2834 : 1'b1;
											assign node2834 = (inp[3]) ? 1'b0 : 1'b1;

endmodule