module dtc_split66_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node11;
	wire [16-1:0] node14;
	wire [16-1:0] node17;
	wire [16-1:0] node18;
	wire [16-1:0] node21;
	wire [16-1:0] node24;
	wire [16-1:0] node25;
	wire [16-1:0] node26;
	wire [16-1:0] node29;
	wire [16-1:0] node32;
	wire [16-1:0] node33;
	wire [16-1:0] node36;
	wire [16-1:0] node39;
	wire [16-1:0] node40;
	wire [16-1:0] node41;
	wire [16-1:0] node42;
	wire [16-1:0] node45;
	wire [16-1:0] node48;
	wire [16-1:0] node49;
	wire [16-1:0] node52;
	wire [16-1:0] node55;
	wire [16-1:0] node56;
	wire [16-1:0] node57;
	wire [16-1:0] node60;
	wire [16-1:0] node63;
	wire [16-1:0] node64;
	wire [16-1:0] node67;
	wire [16-1:0] node70;
	wire [16-1:0] node71;
	wire [16-1:0] node72;
	wire [16-1:0] node73;
	wire [16-1:0] node74;
	wire [16-1:0] node77;
	wire [16-1:0] node80;
	wire [16-1:0] node81;
	wire [16-1:0] node84;
	wire [16-1:0] node87;
	wire [16-1:0] node88;
	wire [16-1:0] node89;
	wire [16-1:0] node92;
	wire [16-1:0] node95;
	wire [16-1:0] node96;
	wire [16-1:0] node99;
	wire [16-1:0] node102;
	wire [16-1:0] node103;
	wire [16-1:0] node104;
	wire [16-1:0] node105;
	wire [16-1:0] node108;
	wire [16-1:0] node111;
	wire [16-1:0] node112;
	wire [16-1:0] node115;
	wire [16-1:0] node118;
	wire [16-1:0] node119;
	wire [16-1:0] node120;
	wire [16-1:0] node123;
	wire [16-1:0] node126;
	wire [16-1:0] node127;
	wire [16-1:0] node130;
	wire [16-1:0] node133;
	wire [16-1:0] node134;
	wire [16-1:0] node135;
	wire [16-1:0] node136;
	wire [16-1:0] node137;
	wire [16-1:0] node138;
	wire [16-1:0] node141;
	wire [16-1:0] node144;
	wire [16-1:0] node145;
	wire [16-1:0] node148;
	wire [16-1:0] node151;
	wire [16-1:0] node152;
	wire [16-1:0] node153;
	wire [16-1:0] node156;
	wire [16-1:0] node159;
	wire [16-1:0] node160;
	wire [16-1:0] node163;
	wire [16-1:0] node166;
	wire [16-1:0] node167;
	wire [16-1:0] node168;
	wire [16-1:0] node169;
	wire [16-1:0] node172;
	wire [16-1:0] node175;
	wire [16-1:0] node176;
	wire [16-1:0] node179;
	wire [16-1:0] node182;
	wire [16-1:0] node183;
	wire [16-1:0] node184;
	wire [16-1:0] node187;
	wire [16-1:0] node190;
	wire [16-1:0] node191;
	wire [16-1:0] node194;
	wire [16-1:0] node197;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node200;
	wire [16-1:0] node201;
	wire [16-1:0] node204;
	wire [16-1:0] node207;
	wire [16-1:0] node208;
	wire [16-1:0] node211;
	wire [16-1:0] node214;
	wire [16-1:0] node215;
	wire [16-1:0] node216;
	wire [16-1:0] node219;
	wire [16-1:0] node222;
	wire [16-1:0] node223;
	wire [16-1:0] node226;
	wire [16-1:0] node229;
	wire [16-1:0] node230;
	wire [16-1:0] node231;
	wire [16-1:0] node232;
	wire [16-1:0] node235;
	wire [16-1:0] node238;
	wire [16-1:0] node239;
	wire [16-1:0] node242;
	wire [16-1:0] node245;
	wire [16-1:0] node246;
	wire [16-1:0] node247;
	wire [16-1:0] node250;
	wire [16-1:0] node253;
	wire [16-1:0] node254;
	wire [16-1:0] node257;
	wire [16-1:0] node260;
	wire [16-1:0] node261;
	wire [16-1:0] node262;
	wire [16-1:0] node263;
	wire [16-1:0] node264;
	wire [16-1:0] node265;
	wire [16-1:0] node266;
	wire [16-1:0] node269;
	wire [16-1:0] node272;
	wire [16-1:0] node273;
	wire [16-1:0] node276;
	wire [16-1:0] node279;
	wire [16-1:0] node280;
	wire [16-1:0] node281;
	wire [16-1:0] node284;
	wire [16-1:0] node287;
	wire [16-1:0] node288;
	wire [16-1:0] node291;
	wire [16-1:0] node294;
	wire [16-1:0] node295;
	wire [16-1:0] node296;
	wire [16-1:0] node297;
	wire [16-1:0] node300;
	wire [16-1:0] node303;
	wire [16-1:0] node304;
	wire [16-1:0] node307;
	wire [16-1:0] node310;
	wire [16-1:0] node311;
	wire [16-1:0] node312;
	wire [16-1:0] node315;
	wire [16-1:0] node318;
	wire [16-1:0] node319;
	wire [16-1:0] node322;
	wire [16-1:0] node325;
	wire [16-1:0] node326;
	wire [16-1:0] node327;
	wire [16-1:0] node328;
	wire [16-1:0] node329;
	wire [16-1:0] node332;
	wire [16-1:0] node335;
	wire [16-1:0] node336;
	wire [16-1:0] node339;
	wire [16-1:0] node342;
	wire [16-1:0] node343;
	wire [16-1:0] node344;
	wire [16-1:0] node347;
	wire [16-1:0] node350;
	wire [16-1:0] node351;
	wire [16-1:0] node354;
	wire [16-1:0] node357;
	wire [16-1:0] node358;
	wire [16-1:0] node359;
	wire [16-1:0] node360;
	wire [16-1:0] node363;
	wire [16-1:0] node366;
	wire [16-1:0] node367;
	wire [16-1:0] node370;
	wire [16-1:0] node373;
	wire [16-1:0] node374;
	wire [16-1:0] node375;
	wire [16-1:0] node378;
	wire [16-1:0] node381;
	wire [16-1:0] node382;
	wire [16-1:0] node385;
	wire [16-1:0] node388;
	wire [16-1:0] node389;
	wire [16-1:0] node390;
	wire [16-1:0] node391;
	wire [16-1:0] node392;
	wire [16-1:0] node393;
	wire [16-1:0] node396;
	wire [16-1:0] node399;
	wire [16-1:0] node400;
	wire [16-1:0] node403;
	wire [16-1:0] node406;
	wire [16-1:0] node407;
	wire [16-1:0] node408;
	wire [16-1:0] node411;
	wire [16-1:0] node414;
	wire [16-1:0] node415;
	wire [16-1:0] node418;
	wire [16-1:0] node421;
	wire [16-1:0] node422;
	wire [16-1:0] node423;
	wire [16-1:0] node424;
	wire [16-1:0] node427;
	wire [16-1:0] node430;
	wire [16-1:0] node431;
	wire [16-1:0] node434;
	wire [16-1:0] node437;
	wire [16-1:0] node438;
	wire [16-1:0] node439;
	wire [16-1:0] node442;
	wire [16-1:0] node445;
	wire [16-1:0] node446;
	wire [16-1:0] node449;
	wire [16-1:0] node452;
	wire [16-1:0] node453;
	wire [16-1:0] node454;
	wire [16-1:0] node455;
	wire [16-1:0] node456;
	wire [16-1:0] node459;
	wire [16-1:0] node462;
	wire [16-1:0] node463;
	wire [16-1:0] node466;
	wire [16-1:0] node469;
	wire [16-1:0] node470;
	wire [16-1:0] node471;
	wire [16-1:0] node474;
	wire [16-1:0] node477;
	wire [16-1:0] node478;
	wire [16-1:0] node481;
	wire [16-1:0] node484;
	wire [16-1:0] node485;
	wire [16-1:0] node486;
	wire [16-1:0] node487;
	wire [16-1:0] node490;
	wire [16-1:0] node493;
	wire [16-1:0] node494;
	wire [16-1:0] node497;
	wire [16-1:0] node500;
	wire [16-1:0] node501;
	wire [16-1:0] node502;
	wire [16-1:0] node505;
	wire [16-1:0] node508;
	wire [16-1:0] node509;
	wire [16-1:0] node512;
	wire [16-1:0] node515;
	wire [16-1:0] node516;
	wire [16-1:0] node517;
	wire [16-1:0] node518;
	wire [16-1:0] node519;
	wire [16-1:0] node520;
	wire [16-1:0] node521;
	wire [16-1:0] node522;
	wire [16-1:0] node525;
	wire [16-1:0] node528;
	wire [16-1:0] node529;
	wire [16-1:0] node532;
	wire [16-1:0] node535;
	wire [16-1:0] node536;
	wire [16-1:0] node537;
	wire [16-1:0] node540;
	wire [16-1:0] node543;
	wire [16-1:0] node544;
	wire [16-1:0] node547;
	wire [16-1:0] node550;
	wire [16-1:0] node551;
	wire [16-1:0] node552;
	wire [16-1:0] node553;
	wire [16-1:0] node556;
	wire [16-1:0] node559;
	wire [16-1:0] node560;
	wire [16-1:0] node563;
	wire [16-1:0] node566;
	wire [16-1:0] node567;
	wire [16-1:0] node568;
	wire [16-1:0] node571;
	wire [16-1:0] node574;
	wire [16-1:0] node575;
	wire [16-1:0] node578;
	wire [16-1:0] node581;
	wire [16-1:0] node582;
	wire [16-1:0] node583;
	wire [16-1:0] node584;
	wire [16-1:0] node585;
	wire [16-1:0] node588;
	wire [16-1:0] node591;
	wire [16-1:0] node592;
	wire [16-1:0] node595;
	wire [16-1:0] node598;
	wire [16-1:0] node599;
	wire [16-1:0] node600;
	wire [16-1:0] node603;
	wire [16-1:0] node606;
	wire [16-1:0] node607;
	wire [16-1:0] node610;
	wire [16-1:0] node613;
	wire [16-1:0] node614;
	wire [16-1:0] node615;
	wire [16-1:0] node616;
	wire [16-1:0] node619;
	wire [16-1:0] node622;
	wire [16-1:0] node623;
	wire [16-1:0] node626;
	wire [16-1:0] node629;
	wire [16-1:0] node630;
	wire [16-1:0] node631;
	wire [16-1:0] node634;
	wire [16-1:0] node637;
	wire [16-1:0] node638;
	wire [16-1:0] node641;
	wire [16-1:0] node644;
	wire [16-1:0] node645;
	wire [16-1:0] node646;
	wire [16-1:0] node647;
	wire [16-1:0] node648;
	wire [16-1:0] node649;
	wire [16-1:0] node652;
	wire [16-1:0] node655;
	wire [16-1:0] node656;
	wire [16-1:0] node659;
	wire [16-1:0] node662;
	wire [16-1:0] node663;
	wire [16-1:0] node664;
	wire [16-1:0] node667;
	wire [16-1:0] node670;
	wire [16-1:0] node671;
	wire [16-1:0] node674;
	wire [16-1:0] node677;
	wire [16-1:0] node678;
	wire [16-1:0] node679;
	wire [16-1:0] node680;
	wire [16-1:0] node683;
	wire [16-1:0] node686;
	wire [16-1:0] node687;
	wire [16-1:0] node690;
	wire [16-1:0] node693;
	wire [16-1:0] node694;
	wire [16-1:0] node695;
	wire [16-1:0] node698;
	wire [16-1:0] node701;
	wire [16-1:0] node702;
	wire [16-1:0] node705;
	wire [16-1:0] node708;
	wire [16-1:0] node709;
	wire [16-1:0] node710;
	wire [16-1:0] node711;
	wire [16-1:0] node712;
	wire [16-1:0] node715;
	wire [16-1:0] node718;
	wire [16-1:0] node719;
	wire [16-1:0] node722;
	wire [16-1:0] node725;
	wire [16-1:0] node726;
	wire [16-1:0] node727;
	wire [16-1:0] node730;
	wire [16-1:0] node733;
	wire [16-1:0] node734;
	wire [16-1:0] node737;
	wire [16-1:0] node740;
	wire [16-1:0] node741;
	wire [16-1:0] node742;
	wire [16-1:0] node743;
	wire [16-1:0] node746;
	wire [16-1:0] node749;
	wire [16-1:0] node750;
	wire [16-1:0] node753;
	wire [16-1:0] node756;
	wire [16-1:0] node757;
	wire [16-1:0] node758;
	wire [16-1:0] node761;
	wire [16-1:0] node764;
	wire [16-1:0] node765;
	wire [16-1:0] node768;
	wire [16-1:0] node771;
	wire [16-1:0] node772;
	wire [16-1:0] node773;
	wire [16-1:0] node774;
	wire [16-1:0] node775;
	wire [16-1:0] node776;
	wire [16-1:0] node777;
	wire [16-1:0] node780;
	wire [16-1:0] node783;
	wire [16-1:0] node784;
	wire [16-1:0] node787;
	wire [16-1:0] node790;
	wire [16-1:0] node791;
	wire [16-1:0] node792;
	wire [16-1:0] node795;
	wire [16-1:0] node798;
	wire [16-1:0] node799;
	wire [16-1:0] node802;
	wire [16-1:0] node805;
	wire [16-1:0] node806;
	wire [16-1:0] node807;
	wire [16-1:0] node808;
	wire [16-1:0] node811;
	wire [16-1:0] node814;
	wire [16-1:0] node815;
	wire [16-1:0] node818;
	wire [16-1:0] node821;
	wire [16-1:0] node822;
	wire [16-1:0] node823;
	wire [16-1:0] node826;
	wire [16-1:0] node829;
	wire [16-1:0] node830;
	wire [16-1:0] node833;
	wire [16-1:0] node836;
	wire [16-1:0] node837;
	wire [16-1:0] node838;
	wire [16-1:0] node839;
	wire [16-1:0] node840;
	wire [16-1:0] node843;
	wire [16-1:0] node846;
	wire [16-1:0] node847;
	wire [16-1:0] node850;
	wire [16-1:0] node853;
	wire [16-1:0] node854;
	wire [16-1:0] node855;
	wire [16-1:0] node858;
	wire [16-1:0] node861;
	wire [16-1:0] node862;
	wire [16-1:0] node865;
	wire [16-1:0] node868;
	wire [16-1:0] node869;
	wire [16-1:0] node870;
	wire [16-1:0] node871;
	wire [16-1:0] node874;
	wire [16-1:0] node877;
	wire [16-1:0] node878;
	wire [16-1:0] node881;
	wire [16-1:0] node884;
	wire [16-1:0] node885;
	wire [16-1:0] node886;
	wire [16-1:0] node889;
	wire [16-1:0] node892;
	wire [16-1:0] node893;
	wire [16-1:0] node896;
	wire [16-1:0] node899;
	wire [16-1:0] node900;
	wire [16-1:0] node901;
	wire [16-1:0] node902;
	wire [16-1:0] node903;
	wire [16-1:0] node904;
	wire [16-1:0] node907;
	wire [16-1:0] node910;
	wire [16-1:0] node911;
	wire [16-1:0] node914;
	wire [16-1:0] node917;
	wire [16-1:0] node918;
	wire [16-1:0] node919;
	wire [16-1:0] node922;
	wire [16-1:0] node925;
	wire [16-1:0] node926;
	wire [16-1:0] node929;
	wire [16-1:0] node932;
	wire [16-1:0] node933;
	wire [16-1:0] node934;
	wire [16-1:0] node935;
	wire [16-1:0] node938;
	wire [16-1:0] node941;
	wire [16-1:0] node942;
	wire [16-1:0] node945;
	wire [16-1:0] node948;
	wire [16-1:0] node949;
	wire [16-1:0] node950;
	wire [16-1:0] node953;
	wire [16-1:0] node956;
	wire [16-1:0] node957;
	wire [16-1:0] node960;
	wire [16-1:0] node963;
	wire [16-1:0] node964;
	wire [16-1:0] node965;
	wire [16-1:0] node966;
	wire [16-1:0] node967;
	wire [16-1:0] node970;
	wire [16-1:0] node973;
	wire [16-1:0] node974;
	wire [16-1:0] node977;
	wire [16-1:0] node980;
	wire [16-1:0] node981;
	wire [16-1:0] node982;
	wire [16-1:0] node985;
	wire [16-1:0] node988;
	wire [16-1:0] node989;
	wire [16-1:0] node992;
	wire [16-1:0] node995;
	wire [16-1:0] node996;
	wire [16-1:0] node997;
	wire [16-1:0] node998;
	wire [16-1:0] node1001;
	wire [16-1:0] node1004;
	wire [16-1:0] node1005;
	wire [16-1:0] node1008;
	wire [16-1:0] node1011;
	wire [16-1:0] node1012;
	wire [16-1:0] node1013;
	wire [16-1:0] node1016;
	wire [16-1:0] node1019;
	wire [16-1:0] node1020;
	wire [16-1:0] node1023;
	wire [16-1:0] node1026;
	wire [16-1:0] node1027;
	wire [16-1:0] node1028;
	wire [16-1:0] node1029;
	wire [16-1:0] node1030;
	wire [16-1:0] node1031;
	wire [16-1:0] node1032;
	wire [16-1:0] node1033;
	wire [16-1:0] node1034;
	wire [16-1:0] node1037;
	wire [16-1:0] node1040;
	wire [16-1:0] node1041;
	wire [16-1:0] node1044;
	wire [16-1:0] node1047;
	wire [16-1:0] node1048;
	wire [16-1:0] node1049;
	wire [16-1:0] node1052;
	wire [16-1:0] node1055;
	wire [16-1:0] node1056;
	wire [16-1:0] node1059;
	wire [16-1:0] node1062;
	wire [16-1:0] node1063;
	wire [16-1:0] node1064;
	wire [16-1:0] node1065;
	wire [16-1:0] node1068;
	wire [16-1:0] node1071;
	wire [16-1:0] node1072;
	wire [16-1:0] node1075;
	wire [16-1:0] node1078;
	wire [16-1:0] node1079;
	wire [16-1:0] node1080;
	wire [16-1:0] node1083;
	wire [16-1:0] node1086;
	wire [16-1:0] node1087;
	wire [16-1:0] node1090;
	wire [16-1:0] node1093;
	wire [16-1:0] node1094;
	wire [16-1:0] node1095;
	wire [16-1:0] node1096;
	wire [16-1:0] node1097;
	wire [16-1:0] node1100;
	wire [16-1:0] node1103;
	wire [16-1:0] node1104;
	wire [16-1:0] node1107;
	wire [16-1:0] node1110;
	wire [16-1:0] node1111;
	wire [16-1:0] node1112;
	wire [16-1:0] node1115;
	wire [16-1:0] node1118;
	wire [16-1:0] node1119;
	wire [16-1:0] node1122;
	wire [16-1:0] node1125;
	wire [16-1:0] node1126;
	wire [16-1:0] node1127;
	wire [16-1:0] node1128;
	wire [16-1:0] node1131;
	wire [16-1:0] node1134;
	wire [16-1:0] node1135;
	wire [16-1:0] node1138;
	wire [16-1:0] node1141;
	wire [16-1:0] node1142;
	wire [16-1:0] node1143;
	wire [16-1:0] node1146;
	wire [16-1:0] node1149;
	wire [16-1:0] node1150;
	wire [16-1:0] node1153;
	wire [16-1:0] node1156;
	wire [16-1:0] node1157;
	wire [16-1:0] node1158;
	wire [16-1:0] node1159;
	wire [16-1:0] node1160;
	wire [16-1:0] node1161;
	wire [16-1:0] node1164;
	wire [16-1:0] node1167;
	wire [16-1:0] node1168;
	wire [16-1:0] node1171;
	wire [16-1:0] node1174;
	wire [16-1:0] node1175;
	wire [16-1:0] node1176;
	wire [16-1:0] node1179;
	wire [16-1:0] node1182;
	wire [16-1:0] node1183;
	wire [16-1:0] node1186;
	wire [16-1:0] node1189;
	wire [16-1:0] node1190;
	wire [16-1:0] node1191;
	wire [16-1:0] node1192;
	wire [16-1:0] node1195;
	wire [16-1:0] node1198;
	wire [16-1:0] node1199;
	wire [16-1:0] node1202;
	wire [16-1:0] node1205;
	wire [16-1:0] node1206;
	wire [16-1:0] node1207;
	wire [16-1:0] node1210;
	wire [16-1:0] node1213;
	wire [16-1:0] node1214;
	wire [16-1:0] node1217;
	wire [16-1:0] node1220;
	wire [16-1:0] node1221;
	wire [16-1:0] node1222;
	wire [16-1:0] node1223;
	wire [16-1:0] node1224;
	wire [16-1:0] node1227;
	wire [16-1:0] node1230;
	wire [16-1:0] node1231;
	wire [16-1:0] node1234;
	wire [16-1:0] node1237;
	wire [16-1:0] node1238;
	wire [16-1:0] node1239;
	wire [16-1:0] node1242;
	wire [16-1:0] node1245;
	wire [16-1:0] node1246;
	wire [16-1:0] node1249;
	wire [16-1:0] node1252;
	wire [16-1:0] node1253;
	wire [16-1:0] node1254;
	wire [16-1:0] node1255;
	wire [16-1:0] node1258;
	wire [16-1:0] node1261;
	wire [16-1:0] node1262;
	wire [16-1:0] node1265;
	wire [16-1:0] node1268;
	wire [16-1:0] node1269;
	wire [16-1:0] node1270;
	wire [16-1:0] node1273;
	wire [16-1:0] node1276;
	wire [16-1:0] node1277;
	wire [16-1:0] node1280;
	wire [16-1:0] node1283;
	wire [16-1:0] node1284;
	wire [16-1:0] node1285;
	wire [16-1:0] node1286;
	wire [16-1:0] node1287;
	wire [16-1:0] node1288;
	wire [16-1:0] node1289;
	wire [16-1:0] node1292;
	wire [16-1:0] node1295;
	wire [16-1:0] node1296;
	wire [16-1:0] node1299;
	wire [16-1:0] node1302;
	wire [16-1:0] node1303;
	wire [16-1:0] node1304;
	wire [16-1:0] node1307;
	wire [16-1:0] node1310;
	wire [16-1:0] node1311;
	wire [16-1:0] node1314;
	wire [16-1:0] node1317;
	wire [16-1:0] node1318;
	wire [16-1:0] node1319;
	wire [16-1:0] node1320;
	wire [16-1:0] node1323;
	wire [16-1:0] node1326;
	wire [16-1:0] node1327;
	wire [16-1:0] node1330;
	wire [16-1:0] node1333;
	wire [16-1:0] node1334;
	wire [16-1:0] node1335;
	wire [16-1:0] node1338;
	wire [16-1:0] node1341;
	wire [16-1:0] node1342;
	wire [16-1:0] node1345;
	wire [16-1:0] node1348;
	wire [16-1:0] node1349;
	wire [16-1:0] node1350;
	wire [16-1:0] node1351;
	wire [16-1:0] node1352;
	wire [16-1:0] node1355;
	wire [16-1:0] node1358;
	wire [16-1:0] node1359;
	wire [16-1:0] node1362;
	wire [16-1:0] node1365;
	wire [16-1:0] node1366;
	wire [16-1:0] node1367;
	wire [16-1:0] node1370;
	wire [16-1:0] node1373;
	wire [16-1:0] node1374;
	wire [16-1:0] node1377;
	wire [16-1:0] node1380;
	wire [16-1:0] node1381;
	wire [16-1:0] node1382;
	wire [16-1:0] node1383;
	wire [16-1:0] node1386;
	wire [16-1:0] node1389;
	wire [16-1:0] node1390;
	wire [16-1:0] node1393;
	wire [16-1:0] node1396;
	wire [16-1:0] node1397;
	wire [16-1:0] node1398;
	wire [16-1:0] node1401;
	wire [16-1:0] node1404;
	wire [16-1:0] node1405;
	wire [16-1:0] node1408;
	wire [16-1:0] node1411;
	wire [16-1:0] node1412;
	wire [16-1:0] node1413;
	wire [16-1:0] node1414;
	wire [16-1:0] node1415;
	wire [16-1:0] node1416;
	wire [16-1:0] node1419;
	wire [16-1:0] node1422;
	wire [16-1:0] node1423;
	wire [16-1:0] node1426;
	wire [16-1:0] node1429;
	wire [16-1:0] node1430;
	wire [16-1:0] node1431;
	wire [16-1:0] node1434;
	wire [16-1:0] node1437;
	wire [16-1:0] node1438;
	wire [16-1:0] node1441;
	wire [16-1:0] node1444;
	wire [16-1:0] node1445;
	wire [16-1:0] node1446;
	wire [16-1:0] node1447;
	wire [16-1:0] node1450;
	wire [16-1:0] node1453;
	wire [16-1:0] node1454;
	wire [16-1:0] node1457;
	wire [16-1:0] node1460;
	wire [16-1:0] node1461;
	wire [16-1:0] node1462;
	wire [16-1:0] node1465;
	wire [16-1:0] node1468;
	wire [16-1:0] node1469;
	wire [16-1:0] node1472;
	wire [16-1:0] node1475;
	wire [16-1:0] node1476;
	wire [16-1:0] node1477;
	wire [16-1:0] node1478;
	wire [16-1:0] node1479;
	wire [16-1:0] node1482;
	wire [16-1:0] node1485;
	wire [16-1:0] node1486;
	wire [16-1:0] node1489;
	wire [16-1:0] node1492;
	wire [16-1:0] node1493;
	wire [16-1:0] node1494;
	wire [16-1:0] node1497;
	wire [16-1:0] node1500;
	wire [16-1:0] node1501;
	wire [16-1:0] node1504;
	wire [16-1:0] node1507;
	wire [16-1:0] node1508;
	wire [16-1:0] node1509;
	wire [16-1:0] node1510;
	wire [16-1:0] node1513;
	wire [16-1:0] node1516;
	wire [16-1:0] node1517;
	wire [16-1:0] node1520;
	wire [16-1:0] node1523;
	wire [16-1:0] node1524;
	wire [16-1:0] node1525;
	wire [16-1:0] node1528;
	wire [16-1:0] node1531;
	wire [16-1:0] node1532;
	wire [16-1:0] node1535;
	wire [16-1:0] node1538;
	wire [16-1:0] node1539;
	wire [16-1:0] node1540;
	wire [16-1:0] node1541;
	wire [16-1:0] node1542;
	wire [16-1:0] node1543;
	wire [16-1:0] node1544;
	wire [16-1:0] node1545;
	wire [16-1:0] node1548;
	wire [16-1:0] node1551;
	wire [16-1:0] node1552;
	wire [16-1:0] node1555;
	wire [16-1:0] node1558;
	wire [16-1:0] node1559;
	wire [16-1:0] node1560;
	wire [16-1:0] node1563;
	wire [16-1:0] node1566;
	wire [16-1:0] node1567;
	wire [16-1:0] node1570;
	wire [16-1:0] node1573;
	wire [16-1:0] node1574;
	wire [16-1:0] node1575;
	wire [16-1:0] node1576;
	wire [16-1:0] node1579;
	wire [16-1:0] node1582;
	wire [16-1:0] node1583;
	wire [16-1:0] node1586;
	wire [16-1:0] node1589;
	wire [16-1:0] node1590;
	wire [16-1:0] node1591;
	wire [16-1:0] node1594;
	wire [16-1:0] node1597;
	wire [16-1:0] node1598;
	wire [16-1:0] node1601;
	wire [16-1:0] node1604;
	wire [16-1:0] node1605;
	wire [16-1:0] node1606;
	wire [16-1:0] node1607;
	wire [16-1:0] node1608;
	wire [16-1:0] node1611;
	wire [16-1:0] node1614;
	wire [16-1:0] node1615;
	wire [16-1:0] node1618;
	wire [16-1:0] node1621;
	wire [16-1:0] node1622;
	wire [16-1:0] node1623;
	wire [16-1:0] node1626;
	wire [16-1:0] node1629;
	wire [16-1:0] node1630;
	wire [16-1:0] node1633;
	wire [16-1:0] node1636;
	wire [16-1:0] node1637;
	wire [16-1:0] node1638;
	wire [16-1:0] node1639;
	wire [16-1:0] node1642;
	wire [16-1:0] node1645;
	wire [16-1:0] node1646;
	wire [16-1:0] node1649;
	wire [16-1:0] node1652;
	wire [16-1:0] node1653;
	wire [16-1:0] node1654;
	wire [16-1:0] node1657;
	wire [16-1:0] node1660;
	wire [16-1:0] node1661;
	wire [16-1:0] node1664;
	wire [16-1:0] node1667;
	wire [16-1:0] node1668;
	wire [16-1:0] node1669;
	wire [16-1:0] node1670;
	wire [16-1:0] node1671;
	wire [16-1:0] node1672;
	wire [16-1:0] node1675;
	wire [16-1:0] node1678;
	wire [16-1:0] node1679;
	wire [16-1:0] node1682;
	wire [16-1:0] node1685;
	wire [16-1:0] node1686;
	wire [16-1:0] node1687;
	wire [16-1:0] node1690;
	wire [16-1:0] node1693;
	wire [16-1:0] node1694;
	wire [16-1:0] node1697;
	wire [16-1:0] node1700;
	wire [16-1:0] node1701;
	wire [16-1:0] node1702;
	wire [16-1:0] node1703;
	wire [16-1:0] node1706;
	wire [16-1:0] node1709;
	wire [16-1:0] node1710;
	wire [16-1:0] node1713;
	wire [16-1:0] node1716;
	wire [16-1:0] node1717;
	wire [16-1:0] node1718;
	wire [16-1:0] node1721;
	wire [16-1:0] node1724;
	wire [16-1:0] node1725;
	wire [16-1:0] node1728;
	wire [16-1:0] node1731;
	wire [16-1:0] node1732;
	wire [16-1:0] node1733;
	wire [16-1:0] node1734;
	wire [16-1:0] node1735;
	wire [16-1:0] node1738;
	wire [16-1:0] node1741;
	wire [16-1:0] node1742;
	wire [16-1:0] node1745;
	wire [16-1:0] node1748;
	wire [16-1:0] node1749;
	wire [16-1:0] node1750;
	wire [16-1:0] node1753;
	wire [16-1:0] node1756;
	wire [16-1:0] node1757;
	wire [16-1:0] node1760;
	wire [16-1:0] node1763;
	wire [16-1:0] node1764;
	wire [16-1:0] node1765;
	wire [16-1:0] node1766;
	wire [16-1:0] node1769;
	wire [16-1:0] node1772;
	wire [16-1:0] node1773;
	wire [16-1:0] node1776;
	wire [16-1:0] node1779;
	wire [16-1:0] node1780;
	wire [16-1:0] node1781;
	wire [16-1:0] node1784;
	wire [16-1:0] node1787;
	wire [16-1:0] node1788;
	wire [16-1:0] node1791;
	wire [16-1:0] node1794;
	wire [16-1:0] node1795;
	wire [16-1:0] node1796;
	wire [16-1:0] node1797;
	wire [16-1:0] node1798;
	wire [16-1:0] node1799;
	wire [16-1:0] node1800;
	wire [16-1:0] node1803;
	wire [16-1:0] node1806;
	wire [16-1:0] node1807;
	wire [16-1:0] node1810;
	wire [16-1:0] node1813;
	wire [16-1:0] node1814;
	wire [16-1:0] node1815;
	wire [16-1:0] node1818;
	wire [16-1:0] node1821;
	wire [16-1:0] node1822;
	wire [16-1:0] node1825;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1830;
	wire [16-1:0] node1831;
	wire [16-1:0] node1834;
	wire [16-1:0] node1837;
	wire [16-1:0] node1838;
	wire [16-1:0] node1841;
	wire [16-1:0] node1844;
	wire [16-1:0] node1845;
	wire [16-1:0] node1846;
	wire [16-1:0] node1849;
	wire [16-1:0] node1852;
	wire [16-1:0] node1853;
	wire [16-1:0] node1856;
	wire [16-1:0] node1859;
	wire [16-1:0] node1860;
	wire [16-1:0] node1861;
	wire [16-1:0] node1862;
	wire [16-1:0] node1863;
	wire [16-1:0] node1866;
	wire [16-1:0] node1869;
	wire [16-1:0] node1870;
	wire [16-1:0] node1873;
	wire [16-1:0] node1876;
	wire [16-1:0] node1877;
	wire [16-1:0] node1878;
	wire [16-1:0] node1881;
	wire [16-1:0] node1884;
	wire [16-1:0] node1885;
	wire [16-1:0] node1888;
	wire [16-1:0] node1891;
	wire [16-1:0] node1892;
	wire [16-1:0] node1893;
	wire [16-1:0] node1894;
	wire [16-1:0] node1897;
	wire [16-1:0] node1900;
	wire [16-1:0] node1901;
	wire [16-1:0] node1904;
	wire [16-1:0] node1907;
	wire [16-1:0] node1908;
	wire [16-1:0] node1909;
	wire [16-1:0] node1912;
	wire [16-1:0] node1915;
	wire [16-1:0] node1916;
	wire [16-1:0] node1919;
	wire [16-1:0] node1922;
	wire [16-1:0] node1923;
	wire [16-1:0] node1924;
	wire [16-1:0] node1925;
	wire [16-1:0] node1926;
	wire [16-1:0] node1927;
	wire [16-1:0] node1930;
	wire [16-1:0] node1933;
	wire [16-1:0] node1934;
	wire [16-1:0] node1937;
	wire [16-1:0] node1940;
	wire [16-1:0] node1941;
	wire [16-1:0] node1942;
	wire [16-1:0] node1945;
	wire [16-1:0] node1948;
	wire [16-1:0] node1949;
	wire [16-1:0] node1952;
	wire [16-1:0] node1955;
	wire [16-1:0] node1956;
	wire [16-1:0] node1957;
	wire [16-1:0] node1958;
	wire [16-1:0] node1961;
	wire [16-1:0] node1964;
	wire [16-1:0] node1965;
	wire [16-1:0] node1968;
	wire [16-1:0] node1971;
	wire [16-1:0] node1972;
	wire [16-1:0] node1973;
	wire [16-1:0] node1976;
	wire [16-1:0] node1979;
	wire [16-1:0] node1980;
	wire [16-1:0] node1983;
	wire [16-1:0] node1986;
	wire [16-1:0] node1987;
	wire [16-1:0] node1988;
	wire [16-1:0] node1989;
	wire [16-1:0] node1990;
	wire [16-1:0] node1993;
	wire [16-1:0] node1996;
	wire [16-1:0] node1997;
	wire [16-1:0] node2000;
	wire [16-1:0] node2003;
	wire [16-1:0] node2004;
	wire [16-1:0] node2005;
	wire [16-1:0] node2008;
	wire [16-1:0] node2011;
	wire [16-1:0] node2012;
	wire [16-1:0] node2015;
	wire [16-1:0] node2018;
	wire [16-1:0] node2019;
	wire [16-1:0] node2020;
	wire [16-1:0] node2021;
	wire [16-1:0] node2024;
	wire [16-1:0] node2027;
	wire [16-1:0] node2028;
	wire [16-1:0] node2031;
	wire [16-1:0] node2034;
	wire [16-1:0] node2035;
	wire [16-1:0] node2036;
	wire [16-1:0] node2039;
	wire [16-1:0] node2042;
	wire [16-1:0] node2043;
	wire [16-1:0] node2046;
	wire [16-1:0] node2049;
	wire [16-1:0] node2050;
	wire [16-1:0] node2051;
	wire [16-1:0] node2052;
	wire [16-1:0] node2053;
	wire [16-1:0] node2054;
	wire [16-1:0] node2055;
	wire [16-1:0] node2056;
	wire [16-1:0] node2057;
	wire [16-1:0] node2058;
	wire [16-1:0] node2061;
	wire [16-1:0] node2064;
	wire [16-1:0] node2065;
	wire [16-1:0] node2068;
	wire [16-1:0] node2071;
	wire [16-1:0] node2072;
	wire [16-1:0] node2073;
	wire [16-1:0] node2076;
	wire [16-1:0] node2079;
	wire [16-1:0] node2080;
	wire [16-1:0] node2083;
	wire [16-1:0] node2086;
	wire [16-1:0] node2087;
	wire [16-1:0] node2088;
	wire [16-1:0] node2089;
	wire [16-1:0] node2092;
	wire [16-1:0] node2095;
	wire [16-1:0] node2096;
	wire [16-1:0] node2099;
	wire [16-1:0] node2102;
	wire [16-1:0] node2103;
	wire [16-1:0] node2104;
	wire [16-1:0] node2107;
	wire [16-1:0] node2110;
	wire [16-1:0] node2111;
	wire [16-1:0] node2114;
	wire [16-1:0] node2117;
	wire [16-1:0] node2118;
	wire [16-1:0] node2119;
	wire [16-1:0] node2120;
	wire [16-1:0] node2121;
	wire [16-1:0] node2124;
	wire [16-1:0] node2127;
	wire [16-1:0] node2128;
	wire [16-1:0] node2131;
	wire [16-1:0] node2134;
	wire [16-1:0] node2135;
	wire [16-1:0] node2136;
	wire [16-1:0] node2139;
	wire [16-1:0] node2142;
	wire [16-1:0] node2143;
	wire [16-1:0] node2146;
	wire [16-1:0] node2149;
	wire [16-1:0] node2150;
	wire [16-1:0] node2151;
	wire [16-1:0] node2152;
	wire [16-1:0] node2155;
	wire [16-1:0] node2158;
	wire [16-1:0] node2159;
	wire [16-1:0] node2162;
	wire [16-1:0] node2165;
	wire [16-1:0] node2166;
	wire [16-1:0] node2167;
	wire [16-1:0] node2170;
	wire [16-1:0] node2173;
	wire [16-1:0] node2174;
	wire [16-1:0] node2177;
	wire [16-1:0] node2180;
	wire [16-1:0] node2181;
	wire [16-1:0] node2182;
	wire [16-1:0] node2183;
	wire [16-1:0] node2184;
	wire [16-1:0] node2185;
	wire [16-1:0] node2188;
	wire [16-1:0] node2191;
	wire [16-1:0] node2192;
	wire [16-1:0] node2195;
	wire [16-1:0] node2198;
	wire [16-1:0] node2199;
	wire [16-1:0] node2200;
	wire [16-1:0] node2203;
	wire [16-1:0] node2206;
	wire [16-1:0] node2207;
	wire [16-1:0] node2210;
	wire [16-1:0] node2213;
	wire [16-1:0] node2214;
	wire [16-1:0] node2215;
	wire [16-1:0] node2216;
	wire [16-1:0] node2219;
	wire [16-1:0] node2222;
	wire [16-1:0] node2223;
	wire [16-1:0] node2226;
	wire [16-1:0] node2229;
	wire [16-1:0] node2230;
	wire [16-1:0] node2231;
	wire [16-1:0] node2234;
	wire [16-1:0] node2237;
	wire [16-1:0] node2238;
	wire [16-1:0] node2241;
	wire [16-1:0] node2244;
	wire [16-1:0] node2245;
	wire [16-1:0] node2246;
	wire [16-1:0] node2247;
	wire [16-1:0] node2248;
	wire [16-1:0] node2251;
	wire [16-1:0] node2254;
	wire [16-1:0] node2255;
	wire [16-1:0] node2258;
	wire [16-1:0] node2261;
	wire [16-1:0] node2262;
	wire [16-1:0] node2263;
	wire [16-1:0] node2266;
	wire [16-1:0] node2269;
	wire [16-1:0] node2270;
	wire [16-1:0] node2273;
	wire [16-1:0] node2276;
	wire [16-1:0] node2277;
	wire [16-1:0] node2278;
	wire [16-1:0] node2279;
	wire [16-1:0] node2282;
	wire [16-1:0] node2285;
	wire [16-1:0] node2286;
	wire [16-1:0] node2289;
	wire [16-1:0] node2292;
	wire [16-1:0] node2293;
	wire [16-1:0] node2294;
	wire [16-1:0] node2297;
	wire [16-1:0] node2300;
	wire [16-1:0] node2301;
	wire [16-1:0] node2304;
	wire [16-1:0] node2307;
	wire [16-1:0] node2308;
	wire [16-1:0] node2309;
	wire [16-1:0] node2310;
	wire [16-1:0] node2311;
	wire [16-1:0] node2312;
	wire [16-1:0] node2313;
	wire [16-1:0] node2316;
	wire [16-1:0] node2319;
	wire [16-1:0] node2320;
	wire [16-1:0] node2323;
	wire [16-1:0] node2326;
	wire [16-1:0] node2327;
	wire [16-1:0] node2328;
	wire [16-1:0] node2331;
	wire [16-1:0] node2334;
	wire [16-1:0] node2335;
	wire [16-1:0] node2338;
	wire [16-1:0] node2341;
	wire [16-1:0] node2342;
	wire [16-1:0] node2343;
	wire [16-1:0] node2344;
	wire [16-1:0] node2347;
	wire [16-1:0] node2350;
	wire [16-1:0] node2351;
	wire [16-1:0] node2354;
	wire [16-1:0] node2357;
	wire [16-1:0] node2358;
	wire [16-1:0] node2359;
	wire [16-1:0] node2362;
	wire [16-1:0] node2365;
	wire [16-1:0] node2366;
	wire [16-1:0] node2369;
	wire [16-1:0] node2372;
	wire [16-1:0] node2373;
	wire [16-1:0] node2374;
	wire [16-1:0] node2375;
	wire [16-1:0] node2376;
	wire [16-1:0] node2379;
	wire [16-1:0] node2382;
	wire [16-1:0] node2383;
	wire [16-1:0] node2386;
	wire [16-1:0] node2389;
	wire [16-1:0] node2390;
	wire [16-1:0] node2391;
	wire [16-1:0] node2394;
	wire [16-1:0] node2397;
	wire [16-1:0] node2398;
	wire [16-1:0] node2401;
	wire [16-1:0] node2404;
	wire [16-1:0] node2405;
	wire [16-1:0] node2406;
	wire [16-1:0] node2407;
	wire [16-1:0] node2410;
	wire [16-1:0] node2413;
	wire [16-1:0] node2414;
	wire [16-1:0] node2417;
	wire [16-1:0] node2420;
	wire [16-1:0] node2421;
	wire [16-1:0] node2422;
	wire [16-1:0] node2425;
	wire [16-1:0] node2428;
	wire [16-1:0] node2429;
	wire [16-1:0] node2432;
	wire [16-1:0] node2435;
	wire [16-1:0] node2436;
	wire [16-1:0] node2437;
	wire [16-1:0] node2438;
	wire [16-1:0] node2439;
	wire [16-1:0] node2440;
	wire [16-1:0] node2443;
	wire [16-1:0] node2446;
	wire [16-1:0] node2447;
	wire [16-1:0] node2450;
	wire [16-1:0] node2453;
	wire [16-1:0] node2454;
	wire [16-1:0] node2455;
	wire [16-1:0] node2458;
	wire [16-1:0] node2461;
	wire [16-1:0] node2462;
	wire [16-1:0] node2465;
	wire [16-1:0] node2468;
	wire [16-1:0] node2469;
	wire [16-1:0] node2470;
	wire [16-1:0] node2471;
	wire [16-1:0] node2474;
	wire [16-1:0] node2477;
	wire [16-1:0] node2478;
	wire [16-1:0] node2481;
	wire [16-1:0] node2484;
	wire [16-1:0] node2485;
	wire [16-1:0] node2486;
	wire [16-1:0] node2489;
	wire [16-1:0] node2492;
	wire [16-1:0] node2493;
	wire [16-1:0] node2496;
	wire [16-1:0] node2499;
	wire [16-1:0] node2500;
	wire [16-1:0] node2501;
	wire [16-1:0] node2502;
	wire [16-1:0] node2503;
	wire [16-1:0] node2506;
	wire [16-1:0] node2509;
	wire [16-1:0] node2510;
	wire [16-1:0] node2513;
	wire [16-1:0] node2516;
	wire [16-1:0] node2517;
	wire [16-1:0] node2518;
	wire [16-1:0] node2521;
	wire [16-1:0] node2524;
	wire [16-1:0] node2525;
	wire [16-1:0] node2528;
	wire [16-1:0] node2531;
	wire [16-1:0] node2532;
	wire [16-1:0] node2533;
	wire [16-1:0] node2534;
	wire [16-1:0] node2537;
	wire [16-1:0] node2540;
	wire [16-1:0] node2541;
	wire [16-1:0] node2544;
	wire [16-1:0] node2547;
	wire [16-1:0] node2548;
	wire [16-1:0] node2549;
	wire [16-1:0] node2552;
	wire [16-1:0] node2555;
	wire [16-1:0] node2556;
	wire [16-1:0] node2559;
	wire [16-1:0] node2562;
	wire [16-1:0] node2563;
	wire [16-1:0] node2564;
	wire [16-1:0] node2565;
	wire [16-1:0] node2566;
	wire [16-1:0] node2567;
	wire [16-1:0] node2568;
	wire [16-1:0] node2569;
	wire [16-1:0] node2572;
	wire [16-1:0] node2575;
	wire [16-1:0] node2576;
	wire [16-1:0] node2579;
	wire [16-1:0] node2582;
	wire [16-1:0] node2583;
	wire [16-1:0] node2584;
	wire [16-1:0] node2587;
	wire [16-1:0] node2590;
	wire [16-1:0] node2591;
	wire [16-1:0] node2594;
	wire [16-1:0] node2597;
	wire [16-1:0] node2598;
	wire [16-1:0] node2599;
	wire [16-1:0] node2600;
	wire [16-1:0] node2603;
	wire [16-1:0] node2606;
	wire [16-1:0] node2607;
	wire [16-1:0] node2610;
	wire [16-1:0] node2613;
	wire [16-1:0] node2614;
	wire [16-1:0] node2615;
	wire [16-1:0] node2618;
	wire [16-1:0] node2621;
	wire [16-1:0] node2622;
	wire [16-1:0] node2625;
	wire [16-1:0] node2628;
	wire [16-1:0] node2629;
	wire [16-1:0] node2630;
	wire [16-1:0] node2631;
	wire [16-1:0] node2632;
	wire [16-1:0] node2635;
	wire [16-1:0] node2638;
	wire [16-1:0] node2639;
	wire [16-1:0] node2642;
	wire [16-1:0] node2645;
	wire [16-1:0] node2646;
	wire [16-1:0] node2647;
	wire [16-1:0] node2650;
	wire [16-1:0] node2653;
	wire [16-1:0] node2654;
	wire [16-1:0] node2657;
	wire [16-1:0] node2660;
	wire [16-1:0] node2661;
	wire [16-1:0] node2662;
	wire [16-1:0] node2663;
	wire [16-1:0] node2666;
	wire [16-1:0] node2669;
	wire [16-1:0] node2670;
	wire [16-1:0] node2673;
	wire [16-1:0] node2676;
	wire [16-1:0] node2677;
	wire [16-1:0] node2678;
	wire [16-1:0] node2681;
	wire [16-1:0] node2684;
	wire [16-1:0] node2685;
	wire [16-1:0] node2688;
	wire [16-1:0] node2691;
	wire [16-1:0] node2692;
	wire [16-1:0] node2693;
	wire [16-1:0] node2694;
	wire [16-1:0] node2695;
	wire [16-1:0] node2696;
	wire [16-1:0] node2699;
	wire [16-1:0] node2702;
	wire [16-1:0] node2703;
	wire [16-1:0] node2706;
	wire [16-1:0] node2709;
	wire [16-1:0] node2710;
	wire [16-1:0] node2711;
	wire [16-1:0] node2714;
	wire [16-1:0] node2717;
	wire [16-1:0] node2718;
	wire [16-1:0] node2721;
	wire [16-1:0] node2724;
	wire [16-1:0] node2725;
	wire [16-1:0] node2726;
	wire [16-1:0] node2727;
	wire [16-1:0] node2730;
	wire [16-1:0] node2733;
	wire [16-1:0] node2734;
	wire [16-1:0] node2737;
	wire [16-1:0] node2740;
	wire [16-1:0] node2741;
	wire [16-1:0] node2742;
	wire [16-1:0] node2745;
	wire [16-1:0] node2748;
	wire [16-1:0] node2749;
	wire [16-1:0] node2752;
	wire [16-1:0] node2755;
	wire [16-1:0] node2756;
	wire [16-1:0] node2757;
	wire [16-1:0] node2758;
	wire [16-1:0] node2759;
	wire [16-1:0] node2762;
	wire [16-1:0] node2765;
	wire [16-1:0] node2766;
	wire [16-1:0] node2769;
	wire [16-1:0] node2772;
	wire [16-1:0] node2773;
	wire [16-1:0] node2774;
	wire [16-1:0] node2777;
	wire [16-1:0] node2780;
	wire [16-1:0] node2781;
	wire [16-1:0] node2784;
	wire [16-1:0] node2787;
	wire [16-1:0] node2788;
	wire [16-1:0] node2789;
	wire [16-1:0] node2790;
	wire [16-1:0] node2793;
	wire [16-1:0] node2796;
	wire [16-1:0] node2797;
	wire [16-1:0] node2800;
	wire [16-1:0] node2803;
	wire [16-1:0] node2804;
	wire [16-1:0] node2805;
	wire [16-1:0] node2808;
	wire [16-1:0] node2811;
	wire [16-1:0] node2812;
	wire [16-1:0] node2815;
	wire [16-1:0] node2818;
	wire [16-1:0] node2819;
	wire [16-1:0] node2820;
	wire [16-1:0] node2821;
	wire [16-1:0] node2822;
	wire [16-1:0] node2823;
	wire [16-1:0] node2824;
	wire [16-1:0] node2827;
	wire [16-1:0] node2830;
	wire [16-1:0] node2831;
	wire [16-1:0] node2834;
	wire [16-1:0] node2837;
	wire [16-1:0] node2838;
	wire [16-1:0] node2839;
	wire [16-1:0] node2842;
	wire [16-1:0] node2845;
	wire [16-1:0] node2846;
	wire [16-1:0] node2849;
	wire [16-1:0] node2852;
	wire [16-1:0] node2853;
	wire [16-1:0] node2854;
	wire [16-1:0] node2855;
	wire [16-1:0] node2858;
	wire [16-1:0] node2861;
	wire [16-1:0] node2862;
	wire [16-1:0] node2865;
	wire [16-1:0] node2868;
	wire [16-1:0] node2869;
	wire [16-1:0] node2870;
	wire [16-1:0] node2873;
	wire [16-1:0] node2876;
	wire [16-1:0] node2877;
	wire [16-1:0] node2880;
	wire [16-1:0] node2883;
	wire [16-1:0] node2884;
	wire [16-1:0] node2885;
	wire [16-1:0] node2886;
	wire [16-1:0] node2887;
	wire [16-1:0] node2890;
	wire [16-1:0] node2893;
	wire [16-1:0] node2894;
	wire [16-1:0] node2897;
	wire [16-1:0] node2900;
	wire [16-1:0] node2901;
	wire [16-1:0] node2902;
	wire [16-1:0] node2905;
	wire [16-1:0] node2908;
	wire [16-1:0] node2909;
	wire [16-1:0] node2912;
	wire [16-1:0] node2915;
	wire [16-1:0] node2916;
	wire [16-1:0] node2917;
	wire [16-1:0] node2918;
	wire [16-1:0] node2921;
	wire [16-1:0] node2924;
	wire [16-1:0] node2925;
	wire [16-1:0] node2928;
	wire [16-1:0] node2931;
	wire [16-1:0] node2932;
	wire [16-1:0] node2933;
	wire [16-1:0] node2936;
	wire [16-1:0] node2939;
	wire [16-1:0] node2940;
	wire [16-1:0] node2943;
	wire [16-1:0] node2946;
	wire [16-1:0] node2947;
	wire [16-1:0] node2948;
	wire [16-1:0] node2949;
	wire [16-1:0] node2950;
	wire [16-1:0] node2951;
	wire [16-1:0] node2954;
	wire [16-1:0] node2957;
	wire [16-1:0] node2958;
	wire [16-1:0] node2961;
	wire [16-1:0] node2964;
	wire [16-1:0] node2965;
	wire [16-1:0] node2966;
	wire [16-1:0] node2969;
	wire [16-1:0] node2972;
	wire [16-1:0] node2973;
	wire [16-1:0] node2976;
	wire [16-1:0] node2979;
	wire [16-1:0] node2980;
	wire [16-1:0] node2981;
	wire [16-1:0] node2982;
	wire [16-1:0] node2985;
	wire [16-1:0] node2988;
	wire [16-1:0] node2989;
	wire [16-1:0] node2992;
	wire [16-1:0] node2995;
	wire [16-1:0] node2996;
	wire [16-1:0] node2997;
	wire [16-1:0] node3000;
	wire [16-1:0] node3003;
	wire [16-1:0] node3004;
	wire [16-1:0] node3007;
	wire [16-1:0] node3010;
	wire [16-1:0] node3011;
	wire [16-1:0] node3012;
	wire [16-1:0] node3013;
	wire [16-1:0] node3014;
	wire [16-1:0] node3017;
	wire [16-1:0] node3020;
	wire [16-1:0] node3021;
	wire [16-1:0] node3024;
	wire [16-1:0] node3027;
	wire [16-1:0] node3028;
	wire [16-1:0] node3029;
	wire [16-1:0] node3032;
	wire [16-1:0] node3035;
	wire [16-1:0] node3036;
	wire [16-1:0] node3039;
	wire [16-1:0] node3042;
	wire [16-1:0] node3043;
	wire [16-1:0] node3044;
	wire [16-1:0] node3045;
	wire [16-1:0] node3048;
	wire [16-1:0] node3051;
	wire [16-1:0] node3052;
	wire [16-1:0] node3055;
	wire [16-1:0] node3058;
	wire [16-1:0] node3059;
	wire [16-1:0] node3060;
	wire [16-1:0] node3063;
	wire [16-1:0] node3066;
	wire [16-1:0] node3067;
	wire [16-1:0] node3070;
	wire [16-1:0] node3073;
	wire [16-1:0] node3074;
	wire [16-1:0] node3075;
	wire [16-1:0] node3076;
	wire [16-1:0] node3077;
	wire [16-1:0] node3078;
	wire [16-1:0] node3079;
	wire [16-1:0] node3080;
	wire [16-1:0] node3081;
	wire [16-1:0] node3084;
	wire [16-1:0] node3087;
	wire [16-1:0] node3088;
	wire [16-1:0] node3091;
	wire [16-1:0] node3094;
	wire [16-1:0] node3095;
	wire [16-1:0] node3096;
	wire [16-1:0] node3099;
	wire [16-1:0] node3102;
	wire [16-1:0] node3103;
	wire [16-1:0] node3106;
	wire [16-1:0] node3109;
	wire [16-1:0] node3110;
	wire [16-1:0] node3111;
	wire [16-1:0] node3112;
	wire [16-1:0] node3115;
	wire [16-1:0] node3118;
	wire [16-1:0] node3119;
	wire [16-1:0] node3122;
	wire [16-1:0] node3125;
	wire [16-1:0] node3126;
	wire [16-1:0] node3127;
	wire [16-1:0] node3130;
	wire [16-1:0] node3133;
	wire [16-1:0] node3134;
	wire [16-1:0] node3137;
	wire [16-1:0] node3140;
	wire [16-1:0] node3141;
	wire [16-1:0] node3142;
	wire [16-1:0] node3143;
	wire [16-1:0] node3144;
	wire [16-1:0] node3147;
	wire [16-1:0] node3150;
	wire [16-1:0] node3151;
	wire [16-1:0] node3154;
	wire [16-1:0] node3157;
	wire [16-1:0] node3158;
	wire [16-1:0] node3159;
	wire [16-1:0] node3162;
	wire [16-1:0] node3165;
	wire [16-1:0] node3166;
	wire [16-1:0] node3169;
	wire [16-1:0] node3172;
	wire [16-1:0] node3173;
	wire [16-1:0] node3174;
	wire [16-1:0] node3175;
	wire [16-1:0] node3178;
	wire [16-1:0] node3181;
	wire [16-1:0] node3182;
	wire [16-1:0] node3185;
	wire [16-1:0] node3188;
	wire [16-1:0] node3189;
	wire [16-1:0] node3190;
	wire [16-1:0] node3193;
	wire [16-1:0] node3196;
	wire [16-1:0] node3197;
	wire [16-1:0] node3200;
	wire [16-1:0] node3203;
	wire [16-1:0] node3204;
	wire [16-1:0] node3205;
	wire [16-1:0] node3206;
	wire [16-1:0] node3207;
	wire [16-1:0] node3208;
	wire [16-1:0] node3211;
	wire [16-1:0] node3214;
	wire [16-1:0] node3215;
	wire [16-1:0] node3218;
	wire [16-1:0] node3221;
	wire [16-1:0] node3222;
	wire [16-1:0] node3223;
	wire [16-1:0] node3226;
	wire [16-1:0] node3229;
	wire [16-1:0] node3230;
	wire [16-1:0] node3233;
	wire [16-1:0] node3236;
	wire [16-1:0] node3237;
	wire [16-1:0] node3238;
	wire [16-1:0] node3239;
	wire [16-1:0] node3242;
	wire [16-1:0] node3245;
	wire [16-1:0] node3246;
	wire [16-1:0] node3249;
	wire [16-1:0] node3252;
	wire [16-1:0] node3253;
	wire [16-1:0] node3254;
	wire [16-1:0] node3257;
	wire [16-1:0] node3260;
	wire [16-1:0] node3261;
	wire [16-1:0] node3264;
	wire [16-1:0] node3267;
	wire [16-1:0] node3268;
	wire [16-1:0] node3269;
	wire [16-1:0] node3270;
	wire [16-1:0] node3271;
	wire [16-1:0] node3274;
	wire [16-1:0] node3277;
	wire [16-1:0] node3278;
	wire [16-1:0] node3281;
	wire [16-1:0] node3284;
	wire [16-1:0] node3285;
	wire [16-1:0] node3286;
	wire [16-1:0] node3289;
	wire [16-1:0] node3292;
	wire [16-1:0] node3293;
	wire [16-1:0] node3296;
	wire [16-1:0] node3299;
	wire [16-1:0] node3300;
	wire [16-1:0] node3301;
	wire [16-1:0] node3302;
	wire [16-1:0] node3305;
	wire [16-1:0] node3308;
	wire [16-1:0] node3309;
	wire [16-1:0] node3312;
	wire [16-1:0] node3315;
	wire [16-1:0] node3316;
	wire [16-1:0] node3317;
	wire [16-1:0] node3320;
	wire [16-1:0] node3323;
	wire [16-1:0] node3324;
	wire [16-1:0] node3327;
	wire [16-1:0] node3330;
	wire [16-1:0] node3331;
	wire [16-1:0] node3332;
	wire [16-1:0] node3333;
	wire [16-1:0] node3334;
	wire [16-1:0] node3335;
	wire [16-1:0] node3336;
	wire [16-1:0] node3339;
	wire [16-1:0] node3342;
	wire [16-1:0] node3343;
	wire [16-1:0] node3346;
	wire [16-1:0] node3349;
	wire [16-1:0] node3350;
	wire [16-1:0] node3351;
	wire [16-1:0] node3354;
	wire [16-1:0] node3357;
	wire [16-1:0] node3358;
	wire [16-1:0] node3361;
	wire [16-1:0] node3364;
	wire [16-1:0] node3365;
	wire [16-1:0] node3366;
	wire [16-1:0] node3367;
	wire [16-1:0] node3370;
	wire [16-1:0] node3373;
	wire [16-1:0] node3374;
	wire [16-1:0] node3377;
	wire [16-1:0] node3380;
	wire [16-1:0] node3381;
	wire [16-1:0] node3382;
	wire [16-1:0] node3385;
	wire [16-1:0] node3388;
	wire [16-1:0] node3389;
	wire [16-1:0] node3392;
	wire [16-1:0] node3395;
	wire [16-1:0] node3396;
	wire [16-1:0] node3397;
	wire [16-1:0] node3398;
	wire [16-1:0] node3399;
	wire [16-1:0] node3402;
	wire [16-1:0] node3405;
	wire [16-1:0] node3406;
	wire [16-1:0] node3409;
	wire [16-1:0] node3412;
	wire [16-1:0] node3413;
	wire [16-1:0] node3414;
	wire [16-1:0] node3417;
	wire [16-1:0] node3420;
	wire [16-1:0] node3421;
	wire [16-1:0] node3424;
	wire [16-1:0] node3427;
	wire [16-1:0] node3428;
	wire [16-1:0] node3429;
	wire [16-1:0] node3430;
	wire [16-1:0] node3433;
	wire [16-1:0] node3436;
	wire [16-1:0] node3437;
	wire [16-1:0] node3440;
	wire [16-1:0] node3443;
	wire [16-1:0] node3444;
	wire [16-1:0] node3445;
	wire [16-1:0] node3448;
	wire [16-1:0] node3451;
	wire [16-1:0] node3452;
	wire [16-1:0] node3455;
	wire [16-1:0] node3458;
	wire [16-1:0] node3459;
	wire [16-1:0] node3460;
	wire [16-1:0] node3461;
	wire [16-1:0] node3462;
	wire [16-1:0] node3463;
	wire [16-1:0] node3466;
	wire [16-1:0] node3469;
	wire [16-1:0] node3470;
	wire [16-1:0] node3473;
	wire [16-1:0] node3476;
	wire [16-1:0] node3477;
	wire [16-1:0] node3478;
	wire [16-1:0] node3481;
	wire [16-1:0] node3484;
	wire [16-1:0] node3485;
	wire [16-1:0] node3488;
	wire [16-1:0] node3491;
	wire [16-1:0] node3492;
	wire [16-1:0] node3493;
	wire [16-1:0] node3494;
	wire [16-1:0] node3497;
	wire [16-1:0] node3500;
	wire [16-1:0] node3501;
	wire [16-1:0] node3504;
	wire [16-1:0] node3507;
	wire [16-1:0] node3508;
	wire [16-1:0] node3509;
	wire [16-1:0] node3512;
	wire [16-1:0] node3515;
	wire [16-1:0] node3516;
	wire [16-1:0] node3519;
	wire [16-1:0] node3522;
	wire [16-1:0] node3523;
	wire [16-1:0] node3524;
	wire [16-1:0] node3525;
	wire [16-1:0] node3526;
	wire [16-1:0] node3529;
	wire [16-1:0] node3532;
	wire [16-1:0] node3533;
	wire [16-1:0] node3536;
	wire [16-1:0] node3539;
	wire [16-1:0] node3540;
	wire [16-1:0] node3541;
	wire [16-1:0] node3544;
	wire [16-1:0] node3547;
	wire [16-1:0] node3548;
	wire [16-1:0] node3551;
	wire [16-1:0] node3554;
	wire [16-1:0] node3555;
	wire [16-1:0] node3556;
	wire [16-1:0] node3557;
	wire [16-1:0] node3560;
	wire [16-1:0] node3563;
	wire [16-1:0] node3564;
	wire [16-1:0] node3567;
	wire [16-1:0] node3570;
	wire [16-1:0] node3571;
	wire [16-1:0] node3572;
	wire [16-1:0] node3575;
	wire [16-1:0] node3578;
	wire [16-1:0] node3579;
	wire [16-1:0] node3582;
	wire [16-1:0] node3585;
	wire [16-1:0] node3586;
	wire [16-1:0] node3587;
	wire [16-1:0] node3588;
	wire [16-1:0] node3589;
	wire [16-1:0] node3590;
	wire [16-1:0] node3591;
	wire [16-1:0] node3592;
	wire [16-1:0] node3595;
	wire [16-1:0] node3598;
	wire [16-1:0] node3599;
	wire [16-1:0] node3602;
	wire [16-1:0] node3605;
	wire [16-1:0] node3606;
	wire [16-1:0] node3607;
	wire [16-1:0] node3610;
	wire [16-1:0] node3613;
	wire [16-1:0] node3614;
	wire [16-1:0] node3617;
	wire [16-1:0] node3620;
	wire [16-1:0] node3621;
	wire [16-1:0] node3622;
	wire [16-1:0] node3623;
	wire [16-1:0] node3626;
	wire [16-1:0] node3629;
	wire [16-1:0] node3630;
	wire [16-1:0] node3633;
	wire [16-1:0] node3636;
	wire [16-1:0] node3637;
	wire [16-1:0] node3638;
	wire [16-1:0] node3641;
	wire [16-1:0] node3644;
	wire [16-1:0] node3645;
	wire [16-1:0] node3648;
	wire [16-1:0] node3651;
	wire [16-1:0] node3652;
	wire [16-1:0] node3653;
	wire [16-1:0] node3654;
	wire [16-1:0] node3655;
	wire [16-1:0] node3658;
	wire [16-1:0] node3661;
	wire [16-1:0] node3662;
	wire [16-1:0] node3665;
	wire [16-1:0] node3668;
	wire [16-1:0] node3669;
	wire [16-1:0] node3670;
	wire [16-1:0] node3673;
	wire [16-1:0] node3676;
	wire [16-1:0] node3677;
	wire [16-1:0] node3680;
	wire [16-1:0] node3683;
	wire [16-1:0] node3684;
	wire [16-1:0] node3685;
	wire [16-1:0] node3686;
	wire [16-1:0] node3689;
	wire [16-1:0] node3692;
	wire [16-1:0] node3693;
	wire [16-1:0] node3696;
	wire [16-1:0] node3699;
	wire [16-1:0] node3700;
	wire [16-1:0] node3701;
	wire [16-1:0] node3704;
	wire [16-1:0] node3707;
	wire [16-1:0] node3708;
	wire [16-1:0] node3711;
	wire [16-1:0] node3714;
	wire [16-1:0] node3715;
	wire [16-1:0] node3716;
	wire [16-1:0] node3717;
	wire [16-1:0] node3718;
	wire [16-1:0] node3719;
	wire [16-1:0] node3722;
	wire [16-1:0] node3725;
	wire [16-1:0] node3726;
	wire [16-1:0] node3729;
	wire [16-1:0] node3732;
	wire [16-1:0] node3733;
	wire [16-1:0] node3734;
	wire [16-1:0] node3737;
	wire [16-1:0] node3740;
	wire [16-1:0] node3741;
	wire [16-1:0] node3744;
	wire [16-1:0] node3747;
	wire [16-1:0] node3748;
	wire [16-1:0] node3749;
	wire [16-1:0] node3750;
	wire [16-1:0] node3753;
	wire [16-1:0] node3756;
	wire [16-1:0] node3757;
	wire [16-1:0] node3760;
	wire [16-1:0] node3763;
	wire [16-1:0] node3764;
	wire [16-1:0] node3765;
	wire [16-1:0] node3768;
	wire [16-1:0] node3771;
	wire [16-1:0] node3772;
	wire [16-1:0] node3775;
	wire [16-1:0] node3778;
	wire [16-1:0] node3779;
	wire [16-1:0] node3780;
	wire [16-1:0] node3781;
	wire [16-1:0] node3782;
	wire [16-1:0] node3785;
	wire [16-1:0] node3788;
	wire [16-1:0] node3789;
	wire [16-1:0] node3792;
	wire [16-1:0] node3795;
	wire [16-1:0] node3796;
	wire [16-1:0] node3797;
	wire [16-1:0] node3800;
	wire [16-1:0] node3803;
	wire [16-1:0] node3804;
	wire [16-1:0] node3807;
	wire [16-1:0] node3810;
	wire [16-1:0] node3811;
	wire [16-1:0] node3812;
	wire [16-1:0] node3813;
	wire [16-1:0] node3816;
	wire [16-1:0] node3819;
	wire [16-1:0] node3820;
	wire [16-1:0] node3823;
	wire [16-1:0] node3826;
	wire [16-1:0] node3827;
	wire [16-1:0] node3828;
	wire [16-1:0] node3831;
	wire [16-1:0] node3834;
	wire [16-1:0] node3835;
	wire [16-1:0] node3838;
	wire [16-1:0] node3841;
	wire [16-1:0] node3842;
	wire [16-1:0] node3843;
	wire [16-1:0] node3844;
	wire [16-1:0] node3845;
	wire [16-1:0] node3846;
	wire [16-1:0] node3847;
	wire [16-1:0] node3850;
	wire [16-1:0] node3853;
	wire [16-1:0] node3854;
	wire [16-1:0] node3857;
	wire [16-1:0] node3860;
	wire [16-1:0] node3861;
	wire [16-1:0] node3862;
	wire [16-1:0] node3865;
	wire [16-1:0] node3868;
	wire [16-1:0] node3869;
	wire [16-1:0] node3872;
	wire [16-1:0] node3875;
	wire [16-1:0] node3876;
	wire [16-1:0] node3877;
	wire [16-1:0] node3878;
	wire [16-1:0] node3881;
	wire [16-1:0] node3884;
	wire [16-1:0] node3885;
	wire [16-1:0] node3888;
	wire [16-1:0] node3891;
	wire [16-1:0] node3892;
	wire [16-1:0] node3893;
	wire [16-1:0] node3896;
	wire [16-1:0] node3899;
	wire [16-1:0] node3900;
	wire [16-1:0] node3903;
	wire [16-1:0] node3906;
	wire [16-1:0] node3907;
	wire [16-1:0] node3908;
	wire [16-1:0] node3909;
	wire [16-1:0] node3910;
	wire [16-1:0] node3913;
	wire [16-1:0] node3916;
	wire [16-1:0] node3917;
	wire [16-1:0] node3920;
	wire [16-1:0] node3923;
	wire [16-1:0] node3924;
	wire [16-1:0] node3925;
	wire [16-1:0] node3928;
	wire [16-1:0] node3931;
	wire [16-1:0] node3932;
	wire [16-1:0] node3935;
	wire [16-1:0] node3938;
	wire [16-1:0] node3939;
	wire [16-1:0] node3940;
	wire [16-1:0] node3941;
	wire [16-1:0] node3944;
	wire [16-1:0] node3947;
	wire [16-1:0] node3948;
	wire [16-1:0] node3951;
	wire [16-1:0] node3954;
	wire [16-1:0] node3955;
	wire [16-1:0] node3956;
	wire [16-1:0] node3959;
	wire [16-1:0] node3962;
	wire [16-1:0] node3963;
	wire [16-1:0] node3966;
	wire [16-1:0] node3969;
	wire [16-1:0] node3970;
	wire [16-1:0] node3971;
	wire [16-1:0] node3972;
	wire [16-1:0] node3973;
	wire [16-1:0] node3974;
	wire [16-1:0] node3977;
	wire [16-1:0] node3980;
	wire [16-1:0] node3981;
	wire [16-1:0] node3984;
	wire [16-1:0] node3987;
	wire [16-1:0] node3988;
	wire [16-1:0] node3989;
	wire [16-1:0] node3992;
	wire [16-1:0] node3995;
	wire [16-1:0] node3996;
	wire [16-1:0] node3999;
	wire [16-1:0] node4002;
	wire [16-1:0] node4003;
	wire [16-1:0] node4004;
	wire [16-1:0] node4005;
	wire [16-1:0] node4008;
	wire [16-1:0] node4011;
	wire [16-1:0] node4012;
	wire [16-1:0] node4015;
	wire [16-1:0] node4018;
	wire [16-1:0] node4019;
	wire [16-1:0] node4020;
	wire [16-1:0] node4023;
	wire [16-1:0] node4026;
	wire [16-1:0] node4027;
	wire [16-1:0] node4030;
	wire [16-1:0] node4033;
	wire [16-1:0] node4034;
	wire [16-1:0] node4035;
	wire [16-1:0] node4036;
	wire [16-1:0] node4037;
	wire [16-1:0] node4040;
	wire [16-1:0] node4043;
	wire [16-1:0] node4044;
	wire [16-1:0] node4047;
	wire [16-1:0] node4050;
	wire [16-1:0] node4051;
	wire [16-1:0] node4052;
	wire [16-1:0] node4055;
	wire [16-1:0] node4058;
	wire [16-1:0] node4059;
	wire [16-1:0] node4062;
	wire [16-1:0] node4065;
	wire [16-1:0] node4066;
	wire [16-1:0] node4067;
	wire [16-1:0] node4068;
	wire [16-1:0] node4071;
	wire [16-1:0] node4074;
	wire [16-1:0] node4075;
	wire [16-1:0] node4078;
	wire [16-1:0] node4081;
	wire [16-1:0] node4082;
	wire [16-1:0] node4083;
	wire [16-1:0] node4086;
	wire [16-1:0] node4089;
	wire [16-1:0] node4090;
	wire [16-1:0] node4093;
	wire [16-1:0] node4096;
	wire [16-1:0] node4097;
	wire [16-1:0] node4098;
	wire [16-1:0] node4099;
	wire [16-1:0] node4100;
	wire [16-1:0] node4101;
	wire [16-1:0] node4102;
	wire [16-1:0] node4103;
	wire [16-1:0] node4104;
	wire [16-1:0] node4105;
	wire [16-1:0] node4106;
	wire [16-1:0] node4109;
	wire [16-1:0] node4112;
	wire [16-1:0] node4113;
	wire [16-1:0] node4116;
	wire [16-1:0] node4119;
	wire [16-1:0] node4120;
	wire [16-1:0] node4121;
	wire [16-1:0] node4124;
	wire [16-1:0] node4127;
	wire [16-1:0] node4128;
	wire [16-1:0] node4131;
	wire [16-1:0] node4134;
	wire [16-1:0] node4135;
	wire [16-1:0] node4136;
	wire [16-1:0] node4137;
	wire [16-1:0] node4140;
	wire [16-1:0] node4143;
	wire [16-1:0] node4144;
	wire [16-1:0] node4147;
	wire [16-1:0] node4150;
	wire [16-1:0] node4151;
	wire [16-1:0] node4152;
	wire [16-1:0] node4155;
	wire [16-1:0] node4158;
	wire [16-1:0] node4159;
	wire [16-1:0] node4162;
	wire [16-1:0] node4165;
	wire [16-1:0] node4166;
	wire [16-1:0] node4167;
	wire [16-1:0] node4168;
	wire [16-1:0] node4169;
	wire [16-1:0] node4172;
	wire [16-1:0] node4175;
	wire [16-1:0] node4176;
	wire [16-1:0] node4179;
	wire [16-1:0] node4182;
	wire [16-1:0] node4183;
	wire [16-1:0] node4184;
	wire [16-1:0] node4187;
	wire [16-1:0] node4190;
	wire [16-1:0] node4191;
	wire [16-1:0] node4194;
	wire [16-1:0] node4197;
	wire [16-1:0] node4198;
	wire [16-1:0] node4199;
	wire [16-1:0] node4200;
	wire [16-1:0] node4203;
	wire [16-1:0] node4206;
	wire [16-1:0] node4207;
	wire [16-1:0] node4210;
	wire [16-1:0] node4213;
	wire [16-1:0] node4214;
	wire [16-1:0] node4215;
	wire [16-1:0] node4218;
	wire [16-1:0] node4221;
	wire [16-1:0] node4222;
	wire [16-1:0] node4225;
	wire [16-1:0] node4228;
	wire [16-1:0] node4229;
	wire [16-1:0] node4230;
	wire [16-1:0] node4231;
	wire [16-1:0] node4232;
	wire [16-1:0] node4233;
	wire [16-1:0] node4236;
	wire [16-1:0] node4239;
	wire [16-1:0] node4240;
	wire [16-1:0] node4243;
	wire [16-1:0] node4246;
	wire [16-1:0] node4247;
	wire [16-1:0] node4248;
	wire [16-1:0] node4251;
	wire [16-1:0] node4254;
	wire [16-1:0] node4255;
	wire [16-1:0] node4258;
	wire [16-1:0] node4261;
	wire [16-1:0] node4262;
	wire [16-1:0] node4263;
	wire [16-1:0] node4264;
	wire [16-1:0] node4267;
	wire [16-1:0] node4270;
	wire [16-1:0] node4271;
	wire [16-1:0] node4274;
	wire [16-1:0] node4277;
	wire [16-1:0] node4278;
	wire [16-1:0] node4279;
	wire [16-1:0] node4282;
	wire [16-1:0] node4285;
	wire [16-1:0] node4286;
	wire [16-1:0] node4289;
	wire [16-1:0] node4292;
	wire [16-1:0] node4293;
	wire [16-1:0] node4294;
	wire [16-1:0] node4295;
	wire [16-1:0] node4296;
	wire [16-1:0] node4299;
	wire [16-1:0] node4302;
	wire [16-1:0] node4303;
	wire [16-1:0] node4306;
	wire [16-1:0] node4309;
	wire [16-1:0] node4310;
	wire [16-1:0] node4311;
	wire [16-1:0] node4314;
	wire [16-1:0] node4317;
	wire [16-1:0] node4318;
	wire [16-1:0] node4321;
	wire [16-1:0] node4324;
	wire [16-1:0] node4325;
	wire [16-1:0] node4326;
	wire [16-1:0] node4327;
	wire [16-1:0] node4330;
	wire [16-1:0] node4333;
	wire [16-1:0] node4334;
	wire [16-1:0] node4337;
	wire [16-1:0] node4340;
	wire [16-1:0] node4341;
	wire [16-1:0] node4342;
	wire [16-1:0] node4345;
	wire [16-1:0] node4348;
	wire [16-1:0] node4349;
	wire [16-1:0] node4352;
	wire [16-1:0] node4355;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4358;
	wire [16-1:0] node4359;
	wire [16-1:0] node4360;
	wire [16-1:0] node4361;
	wire [16-1:0] node4364;
	wire [16-1:0] node4367;
	wire [16-1:0] node4368;
	wire [16-1:0] node4371;
	wire [16-1:0] node4374;
	wire [16-1:0] node4375;
	wire [16-1:0] node4376;
	wire [16-1:0] node4379;
	wire [16-1:0] node4382;
	wire [16-1:0] node4383;
	wire [16-1:0] node4386;
	wire [16-1:0] node4389;
	wire [16-1:0] node4390;
	wire [16-1:0] node4391;
	wire [16-1:0] node4392;
	wire [16-1:0] node4395;
	wire [16-1:0] node4398;
	wire [16-1:0] node4399;
	wire [16-1:0] node4402;
	wire [16-1:0] node4405;
	wire [16-1:0] node4406;
	wire [16-1:0] node4407;
	wire [16-1:0] node4410;
	wire [16-1:0] node4413;
	wire [16-1:0] node4414;
	wire [16-1:0] node4417;
	wire [16-1:0] node4420;
	wire [16-1:0] node4421;
	wire [16-1:0] node4422;
	wire [16-1:0] node4423;
	wire [16-1:0] node4424;
	wire [16-1:0] node4427;
	wire [16-1:0] node4430;
	wire [16-1:0] node4431;
	wire [16-1:0] node4434;
	wire [16-1:0] node4437;
	wire [16-1:0] node4438;
	wire [16-1:0] node4439;
	wire [16-1:0] node4442;
	wire [16-1:0] node4445;
	wire [16-1:0] node4446;
	wire [16-1:0] node4449;
	wire [16-1:0] node4452;
	wire [16-1:0] node4453;
	wire [16-1:0] node4454;
	wire [16-1:0] node4455;
	wire [16-1:0] node4458;
	wire [16-1:0] node4461;
	wire [16-1:0] node4462;
	wire [16-1:0] node4465;
	wire [16-1:0] node4468;
	wire [16-1:0] node4469;
	wire [16-1:0] node4470;
	wire [16-1:0] node4473;
	wire [16-1:0] node4476;
	wire [16-1:0] node4477;
	wire [16-1:0] node4480;
	wire [16-1:0] node4483;
	wire [16-1:0] node4484;
	wire [16-1:0] node4485;
	wire [16-1:0] node4486;
	wire [16-1:0] node4487;
	wire [16-1:0] node4488;
	wire [16-1:0] node4491;
	wire [16-1:0] node4494;
	wire [16-1:0] node4495;
	wire [16-1:0] node4498;
	wire [16-1:0] node4501;
	wire [16-1:0] node4502;
	wire [16-1:0] node4503;
	wire [16-1:0] node4506;
	wire [16-1:0] node4509;
	wire [16-1:0] node4510;
	wire [16-1:0] node4513;
	wire [16-1:0] node4516;
	wire [16-1:0] node4517;
	wire [16-1:0] node4518;
	wire [16-1:0] node4519;
	wire [16-1:0] node4522;
	wire [16-1:0] node4525;
	wire [16-1:0] node4526;
	wire [16-1:0] node4529;
	wire [16-1:0] node4532;
	wire [16-1:0] node4533;
	wire [16-1:0] node4534;
	wire [16-1:0] node4537;
	wire [16-1:0] node4540;
	wire [16-1:0] node4541;
	wire [16-1:0] node4544;
	wire [16-1:0] node4547;
	wire [16-1:0] node4548;
	wire [16-1:0] node4549;
	wire [16-1:0] node4550;
	wire [16-1:0] node4551;
	wire [16-1:0] node4554;
	wire [16-1:0] node4557;
	wire [16-1:0] node4558;
	wire [16-1:0] node4561;
	wire [16-1:0] node4564;
	wire [16-1:0] node4565;
	wire [16-1:0] node4566;
	wire [16-1:0] node4569;
	wire [16-1:0] node4572;
	wire [16-1:0] node4573;
	wire [16-1:0] node4576;
	wire [16-1:0] node4579;
	wire [16-1:0] node4580;
	wire [16-1:0] node4581;
	wire [16-1:0] node4582;
	wire [16-1:0] node4585;
	wire [16-1:0] node4588;
	wire [16-1:0] node4589;
	wire [16-1:0] node4592;
	wire [16-1:0] node4595;
	wire [16-1:0] node4596;
	wire [16-1:0] node4597;
	wire [16-1:0] node4600;
	wire [16-1:0] node4603;
	wire [16-1:0] node4604;
	wire [16-1:0] node4607;
	wire [16-1:0] node4610;
	wire [16-1:0] node4611;
	wire [16-1:0] node4612;
	wire [16-1:0] node4613;
	wire [16-1:0] node4614;
	wire [16-1:0] node4615;
	wire [16-1:0] node4616;
	wire [16-1:0] node4617;
	wire [16-1:0] node4620;
	wire [16-1:0] node4623;
	wire [16-1:0] node4624;
	wire [16-1:0] node4627;
	wire [16-1:0] node4630;
	wire [16-1:0] node4631;
	wire [16-1:0] node4632;
	wire [16-1:0] node4635;
	wire [16-1:0] node4638;
	wire [16-1:0] node4639;
	wire [16-1:0] node4642;
	wire [16-1:0] node4645;
	wire [16-1:0] node4646;
	wire [16-1:0] node4647;
	wire [16-1:0] node4648;
	wire [16-1:0] node4651;
	wire [16-1:0] node4654;
	wire [16-1:0] node4655;
	wire [16-1:0] node4658;
	wire [16-1:0] node4661;
	wire [16-1:0] node4662;
	wire [16-1:0] node4663;
	wire [16-1:0] node4666;
	wire [16-1:0] node4669;
	wire [16-1:0] node4670;
	wire [16-1:0] node4673;
	wire [16-1:0] node4676;
	wire [16-1:0] node4677;
	wire [16-1:0] node4678;
	wire [16-1:0] node4679;
	wire [16-1:0] node4680;
	wire [16-1:0] node4683;
	wire [16-1:0] node4686;
	wire [16-1:0] node4687;
	wire [16-1:0] node4690;
	wire [16-1:0] node4693;
	wire [16-1:0] node4694;
	wire [16-1:0] node4695;
	wire [16-1:0] node4698;
	wire [16-1:0] node4701;
	wire [16-1:0] node4702;
	wire [16-1:0] node4705;
	wire [16-1:0] node4708;
	wire [16-1:0] node4709;
	wire [16-1:0] node4710;
	wire [16-1:0] node4711;
	wire [16-1:0] node4714;
	wire [16-1:0] node4717;
	wire [16-1:0] node4718;
	wire [16-1:0] node4721;
	wire [16-1:0] node4724;
	wire [16-1:0] node4725;
	wire [16-1:0] node4726;
	wire [16-1:0] node4729;
	wire [16-1:0] node4732;
	wire [16-1:0] node4733;
	wire [16-1:0] node4736;
	wire [16-1:0] node4739;
	wire [16-1:0] node4740;
	wire [16-1:0] node4741;
	wire [16-1:0] node4742;
	wire [16-1:0] node4743;
	wire [16-1:0] node4744;
	wire [16-1:0] node4747;
	wire [16-1:0] node4750;
	wire [16-1:0] node4751;
	wire [16-1:0] node4754;
	wire [16-1:0] node4757;
	wire [16-1:0] node4758;
	wire [16-1:0] node4759;
	wire [16-1:0] node4762;
	wire [16-1:0] node4765;
	wire [16-1:0] node4766;
	wire [16-1:0] node4769;
	wire [16-1:0] node4772;
	wire [16-1:0] node4773;
	wire [16-1:0] node4774;
	wire [16-1:0] node4775;
	wire [16-1:0] node4778;
	wire [16-1:0] node4781;
	wire [16-1:0] node4782;
	wire [16-1:0] node4785;
	wire [16-1:0] node4788;
	wire [16-1:0] node4789;
	wire [16-1:0] node4790;
	wire [16-1:0] node4793;
	wire [16-1:0] node4796;
	wire [16-1:0] node4797;
	wire [16-1:0] node4800;
	wire [16-1:0] node4803;
	wire [16-1:0] node4804;
	wire [16-1:0] node4805;
	wire [16-1:0] node4806;
	wire [16-1:0] node4807;
	wire [16-1:0] node4810;
	wire [16-1:0] node4813;
	wire [16-1:0] node4814;
	wire [16-1:0] node4817;
	wire [16-1:0] node4820;
	wire [16-1:0] node4821;
	wire [16-1:0] node4822;
	wire [16-1:0] node4825;
	wire [16-1:0] node4828;
	wire [16-1:0] node4829;
	wire [16-1:0] node4832;
	wire [16-1:0] node4835;
	wire [16-1:0] node4836;
	wire [16-1:0] node4837;
	wire [16-1:0] node4838;
	wire [16-1:0] node4841;
	wire [16-1:0] node4844;
	wire [16-1:0] node4845;
	wire [16-1:0] node4848;
	wire [16-1:0] node4851;
	wire [16-1:0] node4852;
	wire [16-1:0] node4853;
	wire [16-1:0] node4856;
	wire [16-1:0] node4859;
	wire [16-1:0] node4860;
	wire [16-1:0] node4863;
	wire [16-1:0] node4866;
	wire [16-1:0] node4867;
	wire [16-1:0] node4868;
	wire [16-1:0] node4869;
	wire [16-1:0] node4870;
	wire [16-1:0] node4871;
	wire [16-1:0] node4872;
	wire [16-1:0] node4875;
	wire [16-1:0] node4878;
	wire [16-1:0] node4879;
	wire [16-1:0] node4882;
	wire [16-1:0] node4885;
	wire [16-1:0] node4886;
	wire [16-1:0] node4887;
	wire [16-1:0] node4890;
	wire [16-1:0] node4893;
	wire [16-1:0] node4894;
	wire [16-1:0] node4897;
	wire [16-1:0] node4900;
	wire [16-1:0] node4901;
	wire [16-1:0] node4902;
	wire [16-1:0] node4903;
	wire [16-1:0] node4906;
	wire [16-1:0] node4909;
	wire [16-1:0] node4910;
	wire [16-1:0] node4913;
	wire [16-1:0] node4916;
	wire [16-1:0] node4917;
	wire [16-1:0] node4918;
	wire [16-1:0] node4921;
	wire [16-1:0] node4924;
	wire [16-1:0] node4925;
	wire [16-1:0] node4928;
	wire [16-1:0] node4931;
	wire [16-1:0] node4932;
	wire [16-1:0] node4933;
	wire [16-1:0] node4934;
	wire [16-1:0] node4935;
	wire [16-1:0] node4938;
	wire [16-1:0] node4941;
	wire [16-1:0] node4942;
	wire [16-1:0] node4945;
	wire [16-1:0] node4948;
	wire [16-1:0] node4949;
	wire [16-1:0] node4950;
	wire [16-1:0] node4953;
	wire [16-1:0] node4956;
	wire [16-1:0] node4957;
	wire [16-1:0] node4960;
	wire [16-1:0] node4963;
	wire [16-1:0] node4964;
	wire [16-1:0] node4965;
	wire [16-1:0] node4966;
	wire [16-1:0] node4969;
	wire [16-1:0] node4972;
	wire [16-1:0] node4973;
	wire [16-1:0] node4976;
	wire [16-1:0] node4979;
	wire [16-1:0] node4980;
	wire [16-1:0] node4981;
	wire [16-1:0] node4984;
	wire [16-1:0] node4987;
	wire [16-1:0] node4988;
	wire [16-1:0] node4991;
	wire [16-1:0] node4994;
	wire [16-1:0] node4995;
	wire [16-1:0] node4996;
	wire [16-1:0] node4997;
	wire [16-1:0] node4998;
	wire [16-1:0] node4999;
	wire [16-1:0] node5002;
	wire [16-1:0] node5005;
	wire [16-1:0] node5006;
	wire [16-1:0] node5009;
	wire [16-1:0] node5012;
	wire [16-1:0] node5013;
	wire [16-1:0] node5014;
	wire [16-1:0] node5017;
	wire [16-1:0] node5020;
	wire [16-1:0] node5021;
	wire [16-1:0] node5024;
	wire [16-1:0] node5027;
	wire [16-1:0] node5028;
	wire [16-1:0] node5029;
	wire [16-1:0] node5030;
	wire [16-1:0] node5033;
	wire [16-1:0] node5036;
	wire [16-1:0] node5037;
	wire [16-1:0] node5040;
	wire [16-1:0] node5043;
	wire [16-1:0] node5044;
	wire [16-1:0] node5045;
	wire [16-1:0] node5048;
	wire [16-1:0] node5051;
	wire [16-1:0] node5052;
	wire [16-1:0] node5055;
	wire [16-1:0] node5058;
	wire [16-1:0] node5059;
	wire [16-1:0] node5060;
	wire [16-1:0] node5061;
	wire [16-1:0] node5062;
	wire [16-1:0] node5065;
	wire [16-1:0] node5068;
	wire [16-1:0] node5069;
	wire [16-1:0] node5072;
	wire [16-1:0] node5075;
	wire [16-1:0] node5076;
	wire [16-1:0] node5077;
	wire [16-1:0] node5080;
	wire [16-1:0] node5083;
	wire [16-1:0] node5084;
	wire [16-1:0] node5087;
	wire [16-1:0] node5090;
	wire [16-1:0] node5091;
	wire [16-1:0] node5092;
	wire [16-1:0] node5093;
	wire [16-1:0] node5096;
	wire [16-1:0] node5099;
	wire [16-1:0] node5100;
	wire [16-1:0] node5103;
	wire [16-1:0] node5106;
	wire [16-1:0] node5107;
	wire [16-1:0] node5108;
	wire [16-1:0] node5111;
	wire [16-1:0] node5114;
	wire [16-1:0] node5115;
	wire [16-1:0] node5118;
	wire [16-1:0] node5121;
	wire [16-1:0] node5122;
	wire [16-1:0] node5123;
	wire [16-1:0] node5124;
	wire [16-1:0] node5125;
	wire [16-1:0] node5126;
	wire [16-1:0] node5127;
	wire [16-1:0] node5128;
	wire [16-1:0] node5129;
	wire [16-1:0] node5132;
	wire [16-1:0] node5135;
	wire [16-1:0] node5136;
	wire [16-1:0] node5139;
	wire [16-1:0] node5142;
	wire [16-1:0] node5143;
	wire [16-1:0] node5144;
	wire [16-1:0] node5147;
	wire [16-1:0] node5150;
	wire [16-1:0] node5151;
	wire [16-1:0] node5154;
	wire [16-1:0] node5157;
	wire [16-1:0] node5158;
	wire [16-1:0] node5159;
	wire [16-1:0] node5160;
	wire [16-1:0] node5163;
	wire [16-1:0] node5166;
	wire [16-1:0] node5167;
	wire [16-1:0] node5170;
	wire [16-1:0] node5173;
	wire [16-1:0] node5174;
	wire [16-1:0] node5175;
	wire [16-1:0] node5178;
	wire [16-1:0] node5181;
	wire [16-1:0] node5182;
	wire [16-1:0] node5185;
	wire [16-1:0] node5188;
	wire [16-1:0] node5189;
	wire [16-1:0] node5190;
	wire [16-1:0] node5191;
	wire [16-1:0] node5192;
	wire [16-1:0] node5195;
	wire [16-1:0] node5198;
	wire [16-1:0] node5199;
	wire [16-1:0] node5202;
	wire [16-1:0] node5205;
	wire [16-1:0] node5206;
	wire [16-1:0] node5207;
	wire [16-1:0] node5210;
	wire [16-1:0] node5213;
	wire [16-1:0] node5214;
	wire [16-1:0] node5217;
	wire [16-1:0] node5220;
	wire [16-1:0] node5221;
	wire [16-1:0] node5222;
	wire [16-1:0] node5223;
	wire [16-1:0] node5226;
	wire [16-1:0] node5229;
	wire [16-1:0] node5230;
	wire [16-1:0] node5233;
	wire [16-1:0] node5236;
	wire [16-1:0] node5237;
	wire [16-1:0] node5238;
	wire [16-1:0] node5241;
	wire [16-1:0] node5244;
	wire [16-1:0] node5245;
	wire [16-1:0] node5248;
	wire [16-1:0] node5251;
	wire [16-1:0] node5252;
	wire [16-1:0] node5253;
	wire [16-1:0] node5254;
	wire [16-1:0] node5255;
	wire [16-1:0] node5256;
	wire [16-1:0] node5259;
	wire [16-1:0] node5262;
	wire [16-1:0] node5263;
	wire [16-1:0] node5266;
	wire [16-1:0] node5269;
	wire [16-1:0] node5270;
	wire [16-1:0] node5271;
	wire [16-1:0] node5274;
	wire [16-1:0] node5277;
	wire [16-1:0] node5278;
	wire [16-1:0] node5281;
	wire [16-1:0] node5284;
	wire [16-1:0] node5285;
	wire [16-1:0] node5286;
	wire [16-1:0] node5287;
	wire [16-1:0] node5290;
	wire [16-1:0] node5293;
	wire [16-1:0] node5294;
	wire [16-1:0] node5297;
	wire [16-1:0] node5300;
	wire [16-1:0] node5301;
	wire [16-1:0] node5302;
	wire [16-1:0] node5305;
	wire [16-1:0] node5308;
	wire [16-1:0] node5309;
	wire [16-1:0] node5312;
	wire [16-1:0] node5315;
	wire [16-1:0] node5316;
	wire [16-1:0] node5317;
	wire [16-1:0] node5318;
	wire [16-1:0] node5319;
	wire [16-1:0] node5322;
	wire [16-1:0] node5325;
	wire [16-1:0] node5326;
	wire [16-1:0] node5329;
	wire [16-1:0] node5332;
	wire [16-1:0] node5333;
	wire [16-1:0] node5334;
	wire [16-1:0] node5337;
	wire [16-1:0] node5340;
	wire [16-1:0] node5341;
	wire [16-1:0] node5344;
	wire [16-1:0] node5347;
	wire [16-1:0] node5348;
	wire [16-1:0] node5349;
	wire [16-1:0] node5350;
	wire [16-1:0] node5353;
	wire [16-1:0] node5356;
	wire [16-1:0] node5357;
	wire [16-1:0] node5360;
	wire [16-1:0] node5363;
	wire [16-1:0] node5364;
	wire [16-1:0] node5365;
	wire [16-1:0] node5368;
	wire [16-1:0] node5371;
	wire [16-1:0] node5372;
	wire [16-1:0] node5375;
	wire [16-1:0] node5378;
	wire [16-1:0] node5379;
	wire [16-1:0] node5380;
	wire [16-1:0] node5381;
	wire [16-1:0] node5382;
	wire [16-1:0] node5383;
	wire [16-1:0] node5384;
	wire [16-1:0] node5387;
	wire [16-1:0] node5390;
	wire [16-1:0] node5391;
	wire [16-1:0] node5394;
	wire [16-1:0] node5397;
	wire [16-1:0] node5398;
	wire [16-1:0] node5399;
	wire [16-1:0] node5402;
	wire [16-1:0] node5405;
	wire [16-1:0] node5406;
	wire [16-1:0] node5409;
	wire [16-1:0] node5412;
	wire [16-1:0] node5413;
	wire [16-1:0] node5414;
	wire [16-1:0] node5415;
	wire [16-1:0] node5418;
	wire [16-1:0] node5421;
	wire [16-1:0] node5422;
	wire [16-1:0] node5425;
	wire [16-1:0] node5428;
	wire [16-1:0] node5429;
	wire [16-1:0] node5430;
	wire [16-1:0] node5433;
	wire [16-1:0] node5436;
	wire [16-1:0] node5437;
	wire [16-1:0] node5440;
	wire [16-1:0] node5443;
	wire [16-1:0] node5444;
	wire [16-1:0] node5445;
	wire [16-1:0] node5446;
	wire [16-1:0] node5447;
	wire [16-1:0] node5450;
	wire [16-1:0] node5453;
	wire [16-1:0] node5454;
	wire [16-1:0] node5457;
	wire [16-1:0] node5460;
	wire [16-1:0] node5461;
	wire [16-1:0] node5462;
	wire [16-1:0] node5465;
	wire [16-1:0] node5468;
	wire [16-1:0] node5469;
	wire [16-1:0] node5472;
	wire [16-1:0] node5475;
	wire [16-1:0] node5476;
	wire [16-1:0] node5477;
	wire [16-1:0] node5478;
	wire [16-1:0] node5481;
	wire [16-1:0] node5484;
	wire [16-1:0] node5485;
	wire [16-1:0] node5488;
	wire [16-1:0] node5491;
	wire [16-1:0] node5492;
	wire [16-1:0] node5493;
	wire [16-1:0] node5496;
	wire [16-1:0] node5499;
	wire [16-1:0] node5500;
	wire [16-1:0] node5503;
	wire [16-1:0] node5506;
	wire [16-1:0] node5507;
	wire [16-1:0] node5508;
	wire [16-1:0] node5509;
	wire [16-1:0] node5510;
	wire [16-1:0] node5511;
	wire [16-1:0] node5514;
	wire [16-1:0] node5517;
	wire [16-1:0] node5518;
	wire [16-1:0] node5521;
	wire [16-1:0] node5524;
	wire [16-1:0] node5525;
	wire [16-1:0] node5526;
	wire [16-1:0] node5529;
	wire [16-1:0] node5532;
	wire [16-1:0] node5533;
	wire [16-1:0] node5536;
	wire [16-1:0] node5539;
	wire [16-1:0] node5540;
	wire [16-1:0] node5541;
	wire [16-1:0] node5542;
	wire [16-1:0] node5545;
	wire [16-1:0] node5548;
	wire [16-1:0] node5549;
	wire [16-1:0] node5552;
	wire [16-1:0] node5555;
	wire [16-1:0] node5556;
	wire [16-1:0] node5557;
	wire [16-1:0] node5560;
	wire [16-1:0] node5563;
	wire [16-1:0] node5564;
	wire [16-1:0] node5567;
	wire [16-1:0] node5570;
	wire [16-1:0] node5571;
	wire [16-1:0] node5572;
	wire [16-1:0] node5573;
	wire [16-1:0] node5574;
	wire [16-1:0] node5577;
	wire [16-1:0] node5580;
	wire [16-1:0] node5581;
	wire [16-1:0] node5584;
	wire [16-1:0] node5587;
	wire [16-1:0] node5588;
	wire [16-1:0] node5589;
	wire [16-1:0] node5592;
	wire [16-1:0] node5595;
	wire [16-1:0] node5596;
	wire [16-1:0] node5599;
	wire [16-1:0] node5602;
	wire [16-1:0] node5603;
	wire [16-1:0] node5604;
	wire [16-1:0] node5605;
	wire [16-1:0] node5608;
	wire [16-1:0] node5611;
	wire [16-1:0] node5612;
	wire [16-1:0] node5615;
	wire [16-1:0] node5618;
	wire [16-1:0] node5619;
	wire [16-1:0] node5620;
	wire [16-1:0] node5623;
	wire [16-1:0] node5626;
	wire [16-1:0] node5627;
	wire [16-1:0] node5630;
	wire [16-1:0] node5633;
	wire [16-1:0] node5634;
	wire [16-1:0] node5635;
	wire [16-1:0] node5636;
	wire [16-1:0] node5637;
	wire [16-1:0] node5638;
	wire [16-1:0] node5639;
	wire [16-1:0] node5640;
	wire [16-1:0] node5643;
	wire [16-1:0] node5646;
	wire [16-1:0] node5647;
	wire [16-1:0] node5650;
	wire [16-1:0] node5653;
	wire [16-1:0] node5654;
	wire [16-1:0] node5655;
	wire [16-1:0] node5658;
	wire [16-1:0] node5661;
	wire [16-1:0] node5662;
	wire [16-1:0] node5665;
	wire [16-1:0] node5668;
	wire [16-1:0] node5669;
	wire [16-1:0] node5670;
	wire [16-1:0] node5671;
	wire [16-1:0] node5674;
	wire [16-1:0] node5677;
	wire [16-1:0] node5678;
	wire [16-1:0] node5681;
	wire [16-1:0] node5684;
	wire [16-1:0] node5685;
	wire [16-1:0] node5686;
	wire [16-1:0] node5689;
	wire [16-1:0] node5692;
	wire [16-1:0] node5693;
	wire [16-1:0] node5696;
	wire [16-1:0] node5699;
	wire [16-1:0] node5700;
	wire [16-1:0] node5701;
	wire [16-1:0] node5702;
	wire [16-1:0] node5703;
	wire [16-1:0] node5706;
	wire [16-1:0] node5709;
	wire [16-1:0] node5710;
	wire [16-1:0] node5713;
	wire [16-1:0] node5716;
	wire [16-1:0] node5717;
	wire [16-1:0] node5718;
	wire [16-1:0] node5721;
	wire [16-1:0] node5724;
	wire [16-1:0] node5725;
	wire [16-1:0] node5728;
	wire [16-1:0] node5731;
	wire [16-1:0] node5732;
	wire [16-1:0] node5733;
	wire [16-1:0] node5734;
	wire [16-1:0] node5737;
	wire [16-1:0] node5740;
	wire [16-1:0] node5741;
	wire [16-1:0] node5744;
	wire [16-1:0] node5747;
	wire [16-1:0] node5748;
	wire [16-1:0] node5749;
	wire [16-1:0] node5752;
	wire [16-1:0] node5755;
	wire [16-1:0] node5756;
	wire [16-1:0] node5759;
	wire [16-1:0] node5762;
	wire [16-1:0] node5763;
	wire [16-1:0] node5764;
	wire [16-1:0] node5765;
	wire [16-1:0] node5766;
	wire [16-1:0] node5767;
	wire [16-1:0] node5770;
	wire [16-1:0] node5773;
	wire [16-1:0] node5774;
	wire [16-1:0] node5777;
	wire [16-1:0] node5780;
	wire [16-1:0] node5781;
	wire [16-1:0] node5782;
	wire [16-1:0] node5785;
	wire [16-1:0] node5788;
	wire [16-1:0] node5789;
	wire [16-1:0] node5792;
	wire [16-1:0] node5795;
	wire [16-1:0] node5796;
	wire [16-1:0] node5797;
	wire [16-1:0] node5798;
	wire [16-1:0] node5801;
	wire [16-1:0] node5804;
	wire [16-1:0] node5805;
	wire [16-1:0] node5808;
	wire [16-1:0] node5811;
	wire [16-1:0] node5812;
	wire [16-1:0] node5813;
	wire [16-1:0] node5816;
	wire [16-1:0] node5819;
	wire [16-1:0] node5820;
	wire [16-1:0] node5823;
	wire [16-1:0] node5826;
	wire [16-1:0] node5827;
	wire [16-1:0] node5828;
	wire [16-1:0] node5829;
	wire [16-1:0] node5830;
	wire [16-1:0] node5833;
	wire [16-1:0] node5836;
	wire [16-1:0] node5837;
	wire [16-1:0] node5840;
	wire [16-1:0] node5843;
	wire [16-1:0] node5844;
	wire [16-1:0] node5845;
	wire [16-1:0] node5848;
	wire [16-1:0] node5851;
	wire [16-1:0] node5852;
	wire [16-1:0] node5855;
	wire [16-1:0] node5858;
	wire [16-1:0] node5859;
	wire [16-1:0] node5860;
	wire [16-1:0] node5861;
	wire [16-1:0] node5864;
	wire [16-1:0] node5867;
	wire [16-1:0] node5868;
	wire [16-1:0] node5871;
	wire [16-1:0] node5874;
	wire [16-1:0] node5875;
	wire [16-1:0] node5876;
	wire [16-1:0] node5879;
	wire [16-1:0] node5882;
	wire [16-1:0] node5883;
	wire [16-1:0] node5886;
	wire [16-1:0] node5889;
	wire [16-1:0] node5890;
	wire [16-1:0] node5891;
	wire [16-1:0] node5892;
	wire [16-1:0] node5893;
	wire [16-1:0] node5894;
	wire [16-1:0] node5895;
	wire [16-1:0] node5898;
	wire [16-1:0] node5901;
	wire [16-1:0] node5902;
	wire [16-1:0] node5905;
	wire [16-1:0] node5908;
	wire [16-1:0] node5909;
	wire [16-1:0] node5910;
	wire [16-1:0] node5913;
	wire [16-1:0] node5916;
	wire [16-1:0] node5917;
	wire [16-1:0] node5920;
	wire [16-1:0] node5923;
	wire [16-1:0] node5924;
	wire [16-1:0] node5925;
	wire [16-1:0] node5926;
	wire [16-1:0] node5929;
	wire [16-1:0] node5932;
	wire [16-1:0] node5933;
	wire [16-1:0] node5936;
	wire [16-1:0] node5939;
	wire [16-1:0] node5940;
	wire [16-1:0] node5941;
	wire [16-1:0] node5944;
	wire [16-1:0] node5947;
	wire [16-1:0] node5948;
	wire [16-1:0] node5951;
	wire [16-1:0] node5954;
	wire [16-1:0] node5955;
	wire [16-1:0] node5956;
	wire [16-1:0] node5957;
	wire [16-1:0] node5958;
	wire [16-1:0] node5961;
	wire [16-1:0] node5964;
	wire [16-1:0] node5965;
	wire [16-1:0] node5968;
	wire [16-1:0] node5971;
	wire [16-1:0] node5972;
	wire [16-1:0] node5973;
	wire [16-1:0] node5976;
	wire [16-1:0] node5979;
	wire [16-1:0] node5980;
	wire [16-1:0] node5983;
	wire [16-1:0] node5986;
	wire [16-1:0] node5987;
	wire [16-1:0] node5988;
	wire [16-1:0] node5989;
	wire [16-1:0] node5992;
	wire [16-1:0] node5995;
	wire [16-1:0] node5996;
	wire [16-1:0] node5999;
	wire [16-1:0] node6002;
	wire [16-1:0] node6003;
	wire [16-1:0] node6004;
	wire [16-1:0] node6007;
	wire [16-1:0] node6010;
	wire [16-1:0] node6011;
	wire [16-1:0] node6014;
	wire [16-1:0] node6017;
	wire [16-1:0] node6018;
	wire [16-1:0] node6019;
	wire [16-1:0] node6020;
	wire [16-1:0] node6021;
	wire [16-1:0] node6022;
	wire [16-1:0] node6025;
	wire [16-1:0] node6028;
	wire [16-1:0] node6029;
	wire [16-1:0] node6032;
	wire [16-1:0] node6035;
	wire [16-1:0] node6036;
	wire [16-1:0] node6037;
	wire [16-1:0] node6040;
	wire [16-1:0] node6043;
	wire [16-1:0] node6044;
	wire [16-1:0] node6047;
	wire [16-1:0] node6050;
	wire [16-1:0] node6051;
	wire [16-1:0] node6052;
	wire [16-1:0] node6053;
	wire [16-1:0] node6056;
	wire [16-1:0] node6059;
	wire [16-1:0] node6060;
	wire [16-1:0] node6063;
	wire [16-1:0] node6066;
	wire [16-1:0] node6067;
	wire [16-1:0] node6068;
	wire [16-1:0] node6071;
	wire [16-1:0] node6074;
	wire [16-1:0] node6075;
	wire [16-1:0] node6078;
	wire [16-1:0] node6081;
	wire [16-1:0] node6082;
	wire [16-1:0] node6083;
	wire [16-1:0] node6084;
	wire [16-1:0] node6085;
	wire [16-1:0] node6088;
	wire [16-1:0] node6091;
	wire [16-1:0] node6092;
	wire [16-1:0] node6095;
	wire [16-1:0] node6098;
	wire [16-1:0] node6099;
	wire [16-1:0] node6100;
	wire [16-1:0] node6103;
	wire [16-1:0] node6106;
	wire [16-1:0] node6107;
	wire [16-1:0] node6110;
	wire [16-1:0] node6113;
	wire [16-1:0] node6114;
	wire [16-1:0] node6115;
	wire [16-1:0] node6116;
	wire [16-1:0] node6119;
	wire [16-1:0] node6122;
	wire [16-1:0] node6123;
	wire [16-1:0] node6126;
	wire [16-1:0] node6129;
	wire [16-1:0] node6130;
	wire [16-1:0] node6131;
	wire [16-1:0] node6134;
	wire [16-1:0] node6137;
	wire [16-1:0] node6138;
	wire [16-1:0] node6141;
	wire [16-1:0] node6144;
	wire [16-1:0] node6145;
	wire [16-1:0] node6146;
	wire [16-1:0] node6147;
	wire [16-1:0] node6148;
	wire [16-1:0] node6149;
	wire [16-1:0] node6150;
	wire [16-1:0] node6151;
	wire [16-1:0] node6152;
	wire [16-1:0] node6153;
	wire [16-1:0] node6156;
	wire [16-1:0] node6159;
	wire [16-1:0] node6160;
	wire [16-1:0] node6163;
	wire [16-1:0] node6166;
	wire [16-1:0] node6167;
	wire [16-1:0] node6168;
	wire [16-1:0] node6171;
	wire [16-1:0] node6174;
	wire [16-1:0] node6175;
	wire [16-1:0] node6178;
	wire [16-1:0] node6181;
	wire [16-1:0] node6182;
	wire [16-1:0] node6183;
	wire [16-1:0] node6184;
	wire [16-1:0] node6187;
	wire [16-1:0] node6190;
	wire [16-1:0] node6191;
	wire [16-1:0] node6194;
	wire [16-1:0] node6197;
	wire [16-1:0] node6198;
	wire [16-1:0] node6199;
	wire [16-1:0] node6202;
	wire [16-1:0] node6205;
	wire [16-1:0] node6206;
	wire [16-1:0] node6209;
	wire [16-1:0] node6212;
	wire [16-1:0] node6213;
	wire [16-1:0] node6214;
	wire [16-1:0] node6215;
	wire [16-1:0] node6216;
	wire [16-1:0] node6219;
	wire [16-1:0] node6222;
	wire [16-1:0] node6223;
	wire [16-1:0] node6226;
	wire [16-1:0] node6229;
	wire [16-1:0] node6230;
	wire [16-1:0] node6231;
	wire [16-1:0] node6234;
	wire [16-1:0] node6237;
	wire [16-1:0] node6238;
	wire [16-1:0] node6241;
	wire [16-1:0] node6244;
	wire [16-1:0] node6245;
	wire [16-1:0] node6246;
	wire [16-1:0] node6247;
	wire [16-1:0] node6250;
	wire [16-1:0] node6253;
	wire [16-1:0] node6254;
	wire [16-1:0] node6257;
	wire [16-1:0] node6260;
	wire [16-1:0] node6261;
	wire [16-1:0] node6262;
	wire [16-1:0] node6265;
	wire [16-1:0] node6268;
	wire [16-1:0] node6269;
	wire [16-1:0] node6272;
	wire [16-1:0] node6275;
	wire [16-1:0] node6276;
	wire [16-1:0] node6277;
	wire [16-1:0] node6278;
	wire [16-1:0] node6279;
	wire [16-1:0] node6280;
	wire [16-1:0] node6283;
	wire [16-1:0] node6286;
	wire [16-1:0] node6287;
	wire [16-1:0] node6290;
	wire [16-1:0] node6293;
	wire [16-1:0] node6294;
	wire [16-1:0] node6295;
	wire [16-1:0] node6298;
	wire [16-1:0] node6301;
	wire [16-1:0] node6302;
	wire [16-1:0] node6305;
	wire [16-1:0] node6308;
	wire [16-1:0] node6309;
	wire [16-1:0] node6310;
	wire [16-1:0] node6311;
	wire [16-1:0] node6314;
	wire [16-1:0] node6317;
	wire [16-1:0] node6318;
	wire [16-1:0] node6321;
	wire [16-1:0] node6324;
	wire [16-1:0] node6325;
	wire [16-1:0] node6326;
	wire [16-1:0] node6329;
	wire [16-1:0] node6332;
	wire [16-1:0] node6333;
	wire [16-1:0] node6336;
	wire [16-1:0] node6339;
	wire [16-1:0] node6340;
	wire [16-1:0] node6341;
	wire [16-1:0] node6342;
	wire [16-1:0] node6343;
	wire [16-1:0] node6346;
	wire [16-1:0] node6349;
	wire [16-1:0] node6350;
	wire [16-1:0] node6353;
	wire [16-1:0] node6356;
	wire [16-1:0] node6357;
	wire [16-1:0] node6358;
	wire [16-1:0] node6361;
	wire [16-1:0] node6364;
	wire [16-1:0] node6365;
	wire [16-1:0] node6368;
	wire [16-1:0] node6371;
	wire [16-1:0] node6372;
	wire [16-1:0] node6373;
	wire [16-1:0] node6374;
	wire [16-1:0] node6377;
	wire [16-1:0] node6380;
	wire [16-1:0] node6381;
	wire [16-1:0] node6384;
	wire [16-1:0] node6387;
	wire [16-1:0] node6388;
	wire [16-1:0] node6389;
	wire [16-1:0] node6392;
	wire [16-1:0] node6395;
	wire [16-1:0] node6396;
	wire [16-1:0] node6399;
	wire [16-1:0] node6402;
	wire [16-1:0] node6403;
	wire [16-1:0] node6404;
	wire [16-1:0] node6405;
	wire [16-1:0] node6406;
	wire [16-1:0] node6407;
	wire [16-1:0] node6408;
	wire [16-1:0] node6411;
	wire [16-1:0] node6414;
	wire [16-1:0] node6415;
	wire [16-1:0] node6418;
	wire [16-1:0] node6421;
	wire [16-1:0] node6422;
	wire [16-1:0] node6423;
	wire [16-1:0] node6426;
	wire [16-1:0] node6429;
	wire [16-1:0] node6430;
	wire [16-1:0] node6433;
	wire [16-1:0] node6436;
	wire [16-1:0] node6437;
	wire [16-1:0] node6438;
	wire [16-1:0] node6439;
	wire [16-1:0] node6442;
	wire [16-1:0] node6445;
	wire [16-1:0] node6446;
	wire [16-1:0] node6449;
	wire [16-1:0] node6452;
	wire [16-1:0] node6453;
	wire [16-1:0] node6454;
	wire [16-1:0] node6457;
	wire [16-1:0] node6460;
	wire [16-1:0] node6461;
	wire [16-1:0] node6464;
	wire [16-1:0] node6467;
	wire [16-1:0] node6468;
	wire [16-1:0] node6469;
	wire [16-1:0] node6470;
	wire [16-1:0] node6471;
	wire [16-1:0] node6474;
	wire [16-1:0] node6477;
	wire [16-1:0] node6478;
	wire [16-1:0] node6481;
	wire [16-1:0] node6484;
	wire [16-1:0] node6485;
	wire [16-1:0] node6486;
	wire [16-1:0] node6489;
	wire [16-1:0] node6492;
	wire [16-1:0] node6493;
	wire [16-1:0] node6496;
	wire [16-1:0] node6499;
	wire [16-1:0] node6500;
	wire [16-1:0] node6501;
	wire [16-1:0] node6502;
	wire [16-1:0] node6505;
	wire [16-1:0] node6508;
	wire [16-1:0] node6509;
	wire [16-1:0] node6512;
	wire [16-1:0] node6515;
	wire [16-1:0] node6516;
	wire [16-1:0] node6517;
	wire [16-1:0] node6520;
	wire [16-1:0] node6523;
	wire [16-1:0] node6524;
	wire [16-1:0] node6527;
	wire [16-1:0] node6530;
	wire [16-1:0] node6531;
	wire [16-1:0] node6532;
	wire [16-1:0] node6533;
	wire [16-1:0] node6534;
	wire [16-1:0] node6535;
	wire [16-1:0] node6538;
	wire [16-1:0] node6541;
	wire [16-1:0] node6542;
	wire [16-1:0] node6545;
	wire [16-1:0] node6548;
	wire [16-1:0] node6549;
	wire [16-1:0] node6550;
	wire [16-1:0] node6553;
	wire [16-1:0] node6556;
	wire [16-1:0] node6557;
	wire [16-1:0] node6560;
	wire [16-1:0] node6563;
	wire [16-1:0] node6564;
	wire [16-1:0] node6565;
	wire [16-1:0] node6566;
	wire [16-1:0] node6569;
	wire [16-1:0] node6572;
	wire [16-1:0] node6573;
	wire [16-1:0] node6576;
	wire [16-1:0] node6579;
	wire [16-1:0] node6580;
	wire [16-1:0] node6581;
	wire [16-1:0] node6584;
	wire [16-1:0] node6587;
	wire [16-1:0] node6588;
	wire [16-1:0] node6591;
	wire [16-1:0] node6594;
	wire [16-1:0] node6595;
	wire [16-1:0] node6596;
	wire [16-1:0] node6597;
	wire [16-1:0] node6598;
	wire [16-1:0] node6601;
	wire [16-1:0] node6604;
	wire [16-1:0] node6605;
	wire [16-1:0] node6608;
	wire [16-1:0] node6611;
	wire [16-1:0] node6612;
	wire [16-1:0] node6613;
	wire [16-1:0] node6616;
	wire [16-1:0] node6619;
	wire [16-1:0] node6620;
	wire [16-1:0] node6623;
	wire [16-1:0] node6626;
	wire [16-1:0] node6627;
	wire [16-1:0] node6628;
	wire [16-1:0] node6629;
	wire [16-1:0] node6632;
	wire [16-1:0] node6635;
	wire [16-1:0] node6636;
	wire [16-1:0] node6639;
	wire [16-1:0] node6642;
	wire [16-1:0] node6643;
	wire [16-1:0] node6644;
	wire [16-1:0] node6647;
	wire [16-1:0] node6650;
	wire [16-1:0] node6651;
	wire [16-1:0] node6654;
	wire [16-1:0] node6657;
	wire [16-1:0] node6658;
	wire [16-1:0] node6659;
	wire [16-1:0] node6660;
	wire [16-1:0] node6661;
	wire [16-1:0] node6662;
	wire [16-1:0] node6663;
	wire [16-1:0] node6664;
	wire [16-1:0] node6667;
	wire [16-1:0] node6670;
	wire [16-1:0] node6671;
	wire [16-1:0] node6674;
	wire [16-1:0] node6677;
	wire [16-1:0] node6678;
	wire [16-1:0] node6679;
	wire [16-1:0] node6682;
	wire [16-1:0] node6685;
	wire [16-1:0] node6686;
	wire [16-1:0] node6689;
	wire [16-1:0] node6692;
	wire [16-1:0] node6693;
	wire [16-1:0] node6694;
	wire [16-1:0] node6695;
	wire [16-1:0] node6698;
	wire [16-1:0] node6701;
	wire [16-1:0] node6702;
	wire [16-1:0] node6705;
	wire [16-1:0] node6708;
	wire [16-1:0] node6709;
	wire [16-1:0] node6710;
	wire [16-1:0] node6713;
	wire [16-1:0] node6716;
	wire [16-1:0] node6717;
	wire [16-1:0] node6720;
	wire [16-1:0] node6723;
	wire [16-1:0] node6724;
	wire [16-1:0] node6725;
	wire [16-1:0] node6726;
	wire [16-1:0] node6727;
	wire [16-1:0] node6730;
	wire [16-1:0] node6733;
	wire [16-1:0] node6734;
	wire [16-1:0] node6737;
	wire [16-1:0] node6740;
	wire [16-1:0] node6741;
	wire [16-1:0] node6742;
	wire [16-1:0] node6745;
	wire [16-1:0] node6748;
	wire [16-1:0] node6749;
	wire [16-1:0] node6752;
	wire [16-1:0] node6755;
	wire [16-1:0] node6756;
	wire [16-1:0] node6757;
	wire [16-1:0] node6758;
	wire [16-1:0] node6761;
	wire [16-1:0] node6764;
	wire [16-1:0] node6765;
	wire [16-1:0] node6768;
	wire [16-1:0] node6771;
	wire [16-1:0] node6772;
	wire [16-1:0] node6773;
	wire [16-1:0] node6776;
	wire [16-1:0] node6779;
	wire [16-1:0] node6780;
	wire [16-1:0] node6783;
	wire [16-1:0] node6786;
	wire [16-1:0] node6787;
	wire [16-1:0] node6788;
	wire [16-1:0] node6789;
	wire [16-1:0] node6790;
	wire [16-1:0] node6791;
	wire [16-1:0] node6794;
	wire [16-1:0] node6797;
	wire [16-1:0] node6798;
	wire [16-1:0] node6801;
	wire [16-1:0] node6804;
	wire [16-1:0] node6805;
	wire [16-1:0] node6806;
	wire [16-1:0] node6809;
	wire [16-1:0] node6812;
	wire [16-1:0] node6813;
	wire [16-1:0] node6816;
	wire [16-1:0] node6819;
	wire [16-1:0] node6820;
	wire [16-1:0] node6821;
	wire [16-1:0] node6822;
	wire [16-1:0] node6825;
	wire [16-1:0] node6828;
	wire [16-1:0] node6829;
	wire [16-1:0] node6832;
	wire [16-1:0] node6835;
	wire [16-1:0] node6836;
	wire [16-1:0] node6837;
	wire [16-1:0] node6840;
	wire [16-1:0] node6843;
	wire [16-1:0] node6844;
	wire [16-1:0] node6847;
	wire [16-1:0] node6850;
	wire [16-1:0] node6851;
	wire [16-1:0] node6852;
	wire [16-1:0] node6853;
	wire [16-1:0] node6854;
	wire [16-1:0] node6857;
	wire [16-1:0] node6860;
	wire [16-1:0] node6861;
	wire [16-1:0] node6864;
	wire [16-1:0] node6867;
	wire [16-1:0] node6868;
	wire [16-1:0] node6869;
	wire [16-1:0] node6872;
	wire [16-1:0] node6875;
	wire [16-1:0] node6876;
	wire [16-1:0] node6879;
	wire [16-1:0] node6882;
	wire [16-1:0] node6883;
	wire [16-1:0] node6884;
	wire [16-1:0] node6885;
	wire [16-1:0] node6888;
	wire [16-1:0] node6891;
	wire [16-1:0] node6892;
	wire [16-1:0] node6895;
	wire [16-1:0] node6898;
	wire [16-1:0] node6899;
	wire [16-1:0] node6900;
	wire [16-1:0] node6903;
	wire [16-1:0] node6906;
	wire [16-1:0] node6907;
	wire [16-1:0] node6910;
	wire [16-1:0] node6913;
	wire [16-1:0] node6914;
	wire [16-1:0] node6915;
	wire [16-1:0] node6916;
	wire [16-1:0] node6917;
	wire [16-1:0] node6918;
	wire [16-1:0] node6919;
	wire [16-1:0] node6922;
	wire [16-1:0] node6925;
	wire [16-1:0] node6926;
	wire [16-1:0] node6929;
	wire [16-1:0] node6932;
	wire [16-1:0] node6933;
	wire [16-1:0] node6934;
	wire [16-1:0] node6937;
	wire [16-1:0] node6940;
	wire [16-1:0] node6941;
	wire [16-1:0] node6944;
	wire [16-1:0] node6947;
	wire [16-1:0] node6948;
	wire [16-1:0] node6949;
	wire [16-1:0] node6950;
	wire [16-1:0] node6953;
	wire [16-1:0] node6956;
	wire [16-1:0] node6957;
	wire [16-1:0] node6960;
	wire [16-1:0] node6963;
	wire [16-1:0] node6964;
	wire [16-1:0] node6965;
	wire [16-1:0] node6968;
	wire [16-1:0] node6971;
	wire [16-1:0] node6972;
	wire [16-1:0] node6975;
	wire [16-1:0] node6978;
	wire [16-1:0] node6979;
	wire [16-1:0] node6980;
	wire [16-1:0] node6981;
	wire [16-1:0] node6982;
	wire [16-1:0] node6985;
	wire [16-1:0] node6988;
	wire [16-1:0] node6989;
	wire [16-1:0] node6992;
	wire [16-1:0] node6995;
	wire [16-1:0] node6996;
	wire [16-1:0] node6997;
	wire [16-1:0] node7000;
	wire [16-1:0] node7003;
	wire [16-1:0] node7004;
	wire [16-1:0] node7007;
	wire [16-1:0] node7010;
	wire [16-1:0] node7011;
	wire [16-1:0] node7012;
	wire [16-1:0] node7013;
	wire [16-1:0] node7016;
	wire [16-1:0] node7019;
	wire [16-1:0] node7020;
	wire [16-1:0] node7023;
	wire [16-1:0] node7026;
	wire [16-1:0] node7027;
	wire [16-1:0] node7028;
	wire [16-1:0] node7031;
	wire [16-1:0] node7034;
	wire [16-1:0] node7035;
	wire [16-1:0] node7038;
	wire [16-1:0] node7041;
	wire [16-1:0] node7042;
	wire [16-1:0] node7043;
	wire [16-1:0] node7044;
	wire [16-1:0] node7045;
	wire [16-1:0] node7046;
	wire [16-1:0] node7049;
	wire [16-1:0] node7052;
	wire [16-1:0] node7053;
	wire [16-1:0] node7056;
	wire [16-1:0] node7059;
	wire [16-1:0] node7060;
	wire [16-1:0] node7061;
	wire [16-1:0] node7064;
	wire [16-1:0] node7067;
	wire [16-1:0] node7068;
	wire [16-1:0] node7071;
	wire [16-1:0] node7074;
	wire [16-1:0] node7075;
	wire [16-1:0] node7076;
	wire [16-1:0] node7077;
	wire [16-1:0] node7080;
	wire [16-1:0] node7083;
	wire [16-1:0] node7084;
	wire [16-1:0] node7087;
	wire [16-1:0] node7090;
	wire [16-1:0] node7091;
	wire [16-1:0] node7092;
	wire [16-1:0] node7095;
	wire [16-1:0] node7098;
	wire [16-1:0] node7099;
	wire [16-1:0] node7102;
	wire [16-1:0] node7105;
	wire [16-1:0] node7106;
	wire [16-1:0] node7107;
	wire [16-1:0] node7108;
	wire [16-1:0] node7109;
	wire [16-1:0] node7112;
	wire [16-1:0] node7115;
	wire [16-1:0] node7116;
	wire [16-1:0] node7119;
	wire [16-1:0] node7122;
	wire [16-1:0] node7123;
	wire [16-1:0] node7124;
	wire [16-1:0] node7127;
	wire [16-1:0] node7130;
	wire [16-1:0] node7131;
	wire [16-1:0] node7134;
	wire [16-1:0] node7137;
	wire [16-1:0] node7138;
	wire [16-1:0] node7139;
	wire [16-1:0] node7140;
	wire [16-1:0] node7143;
	wire [16-1:0] node7146;
	wire [16-1:0] node7147;
	wire [16-1:0] node7150;
	wire [16-1:0] node7153;
	wire [16-1:0] node7154;
	wire [16-1:0] node7155;
	wire [16-1:0] node7158;
	wire [16-1:0] node7161;
	wire [16-1:0] node7162;
	wire [16-1:0] node7165;
	wire [16-1:0] node7168;
	wire [16-1:0] node7169;
	wire [16-1:0] node7170;
	wire [16-1:0] node7171;
	wire [16-1:0] node7172;
	wire [16-1:0] node7173;
	wire [16-1:0] node7174;
	wire [16-1:0] node7175;
	wire [16-1:0] node7176;
	wire [16-1:0] node7179;
	wire [16-1:0] node7182;
	wire [16-1:0] node7183;
	wire [16-1:0] node7186;
	wire [16-1:0] node7189;
	wire [16-1:0] node7190;
	wire [16-1:0] node7191;
	wire [16-1:0] node7194;
	wire [16-1:0] node7197;
	wire [16-1:0] node7198;
	wire [16-1:0] node7201;
	wire [16-1:0] node7204;
	wire [16-1:0] node7205;
	wire [16-1:0] node7206;
	wire [16-1:0] node7207;
	wire [16-1:0] node7210;
	wire [16-1:0] node7213;
	wire [16-1:0] node7214;
	wire [16-1:0] node7217;
	wire [16-1:0] node7220;
	wire [16-1:0] node7221;
	wire [16-1:0] node7222;
	wire [16-1:0] node7225;
	wire [16-1:0] node7228;
	wire [16-1:0] node7229;
	wire [16-1:0] node7232;
	wire [16-1:0] node7235;
	wire [16-1:0] node7236;
	wire [16-1:0] node7237;
	wire [16-1:0] node7238;
	wire [16-1:0] node7239;
	wire [16-1:0] node7242;
	wire [16-1:0] node7245;
	wire [16-1:0] node7246;
	wire [16-1:0] node7249;
	wire [16-1:0] node7252;
	wire [16-1:0] node7253;
	wire [16-1:0] node7254;
	wire [16-1:0] node7257;
	wire [16-1:0] node7260;
	wire [16-1:0] node7261;
	wire [16-1:0] node7264;
	wire [16-1:0] node7267;
	wire [16-1:0] node7268;
	wire [16-1:0] node7269;
	wire [16-1:0] node7270;
	wire [16-1:0] node7273;
	wire [16-1:0] node7276;
	wire [16-1:0] node7277;
	wire [16-1:0] node7280;
	wire [16-1:0] node7283;
	wire [16-1:0] node7284;
	wire [16-1:0] node7285;
	wire [16-1:0] node7288;
	wire [16-1:0] node7291;
	wire [16-1:0] node7292;
	wire [16-1:0] node7295;
	wire [16-1:0] node7298;
	wire [16-1:0] node7299;
	wire [16-1:0] node7300;
	wire [16-1:0] node7301;
	wire [16-1:0] node7302;
	wire [16-1:0] node7303;
	wire [16-1:0] node7306;
	wire [16-1:0] node7309;
	wire [16-1:0] node7310;
	wire [16-1:0] node7313;
	wire [16-1:0] node7316;
	wire [16-1:0] node7317;
	wire [16-1:0] node7318;
	wire [16-1:0] node7321;
	wire [16-1:0] node7324;
	wire [16-1:0] node7325;
	wire [16-1:0] node7328;
	wire [16-1:0] node7331;
	wire [16-1:0] node7332;
	wire [16-1:0] node7333;
	wire [16-1:0] node7334;
	wire [16-1:0] node7337;
	wire [16-1:0] node7340;
	wire [16-1:0] node7341;
	wire [16-1:0] node7344;
	wire [16-1:0] node7347;
	wire [16-1:0] node7348;
	wire [16-1:0] node7349;
	wire [16-1:0] node7352;
	wire [16-1:0] node7355;
	wire [16-1:0] node7356;
	wire [16-1:0] node7359;
	wire [16-1:0] node7362;
	wire [16-1:0] node7363;
	wire [16-1:0] node7364;
	wire [16-1:0] node7365;
	wire [16-1:0] node7366;
	wire [16-1:0] node7369;
	wire [16-1:0] node7372;
	wire [16-1:0] node7373;
	wire [16-1:0] node7376;
	wire [16-1:0] node7379;
	wire [16-1:0] node7380;
	wire [16-1:0] node7381;
	wire [16-1:0] node7384;
	wire [16-1:0] node7387;
	wire [16-1:0] node7388;
	wire [16-1:0] node7391;
	wire [16-1:0] node7394;
	wire [16-1:0] node7395;
	wire [16-1:0] node7396;
	wire [16-1:0] node7397;
	wire [16-1:0] node7400;
	wire [16-1:0] node7403;
	wire [16-1:0] node7404;
	wire [16-1:0] node7407;
	wire [16-1:0] node7410;
	wire [16-1:0] node7411;
	wire [16-1:0] node7412;
	wire [16-1:0] node7415;
	wire [16-1:0] node7418;
	wire [16-1:0] node7419;
	wire [16-1:0] node7422;
	wire [16-1:0] node7425;
	wire [16-1:0] node7426;
	wire [16-1:0] node7427;
	wire [16-1:0] node7428;
	wire [16-1:0] node7429;
	wire [16-1:0] node7430;
	wire [16-1:0] node7431;
	wire [16-1:0] node7434;
	wire [16-1:0] node7437;
	wire [16-1:0] node7438;
	wire [16-1:0] node7441;
	wire [16-1:0] node7444;
	wire [16-1:0] node7445;
	wire [16-1:0] node7446;
	wire [16-1:0] node7449;
	wire [16-1:0] node7452;
	wire [16-1:0] node7453;
	wire [16-1:0] node7456;
	wire [16-1:0] node7459;
	wire [16-1:0] node7460;
	wire [16-1:0] node7461;
	wire [16-1:0] node7462;
	wire [16-1:0] node7465;
	wire [16-1:0] node7468;
	wire [16-1:0] node7469;
	wire [16-1:0] node7472;
	wire [16-1:0] node7475;
	wire [16-1:0] node7476;
	wire [16-1:0] node7477;
	wire [16-1:0] node7480;
	wire [16-1:0] node7483;
	wire [16-1:0] node7484;
	wire [16-1:0] node7487;
	wire [16-1:0] node7490;
	wire [16-1:0] node7491;
	wire [16-1:0] node7492;
	wire [16-1:0] node7493;
	wire [16-1:0] node7494;
	wire [16-1:0] node7497;
	wire [16-1:0] node7500;
	wire [16-1:0] node7501;
	wire [16-1:0] node7504;
	wire [16-1:0] node7507;
	wire [16-1:0] node7508;
	wire [16-1:0] node7509;
	wire [16-1:0] node7512;
	wire [16-1:0] node7515;
	wire [16-1:0] node7516;
	wire [16-1:0] node7519;
	wire [16-1:0] node7522;
	wire [16-1:0] node7523;
	wire [16-1:0] node7524;
	wire [16-1:0] node7525;
	wire [16-1:0] node7528;
	wire [16-1:0] node7531;
	wire [16-1:0] node7532;
	wire [16-1:0] node7535;
	wire [16-1:0] node7538;
	wire [16-1:0] node7539;
	wire [16-1:0] node7540;
	wire [16-1:0] node7543;
	wire [16-1:0] node7546;
	wire [16-1:0] node7547;
	wire [16-1:0] node7550;
	wire [16-1:0] node7553;
	wire [16-1:0] node7554;
	wire [16-1:0] node7555;
	wire [16-1:0] node7556;
	wire [16-1:0] node7557;
	wire [16-1:0] node7558;
	wire [16-1:0] node7561;
	wire [16-1:0] node7564;
	wire [16-1:0] node7565;
	wire [16-1:0] node7568;
	wire [16-1:0] node7571;
	wire [16-1:0] node7572;
	wire [16-1:0] node7573;
	wire [16-1:0] node7576;
	wire [16-1:0] node7579;
	wire [16-1:0] node7580;
	wire [16-1:0] node7583;
	wire [16-1:0] node7586;
	wire [16-1:0] node7587;
	wire [16-1:0] node7588;
	wire [16-1:0] node7589;
	wire [16-1:0] node7592;
	wire [16-1:0] node7595;
	wire [16-1:0] node7596;
	wire [16-1:0] node7599;
	wire [16-1:0] node7602;
	wire [16-1:0] node7603;
	wire [16-1:0] node7604;
	wire [16-1:0] node7607;
	wire [16-1:0] node7610;
	wire [16-1:0] node7611;
	wire [16-1:0] node7614;
	wire [16-1:0] node7617;
	wire [16-1:0] node7618;
	wire [16-1:0] node7619;
	wire [16-1:0] node7620;
	wire [16-1:0] node7621;
	wire [16-1:0] node7624;
	wire [16-1:0] node7627;
	wire [16-1:0] node7628;
	wire [16-1:0] node7631;
	wire [16-1:0] node7634;
	wire [16-1:0] node7635;
	wire [16-1:0] node7636;
	wire [16-1:0] node7639;
	wire [16-1:0] node7642;
	wire [16-1:0] node7643;
	wire [16-1:0] node7646;
	wire [16-1:0] node7649;
	wire [16-1:0] node7650;
	wire [16-1:0] node7651;
	wire [16-1:0] node7652;
	wire [16-1:0] node7655;
	wire [16-1:0] node7658;
	wire [16-1:0] node7659;
	wire [16-1:0] node7662;
	wire [16-1:0] node7665;
	wire [16-1:0] node7666;
	wire [16-1:0] node7667;
	wire [16-1:0] node7670;
	wire [16-1:0] node7673;
	wire [16-1:0] node7674;
	wire [16-1:0] node7677;
	wire [16-1:0] node7680;
	wire [16-1:0] node7681;
	wire [16-1:0] node7682;
	wire [16-1:0] node7683;
	wire [16-1:0] node7684;
	wire [16-1:0] node7685;
	wire [16-1:0] node7686;
	wire [16-1:0] node7687;
	wire [16-1:0] node7690;
	wire [16-1:0] node7693;
	wire [16-1:0] node7694;
	wire [16-1:0] node7697;
	wire [16-1:0] node7700;
	wire [16-1:0] node7701;
	wire [16-1:0] node7702;
	wire [16-1:0] node7705;
	wire [16-1:0] node7708;
	wire [16-1:0] node7709;
	wire [16-1:0] node7712;
	wire [16-1:0] node7715;
	wire [16-1:0] node7716;
	wire [16-1:0] node7717;
	wire [16-1:0] node7718;
	wire [16-1:0] node7721;
	wire [16-1:0] node7724;
	wire [16-1:0] node7725;
	wire [16-1:0] node7728;
	wire [16-1:0] node7731;
	wire [16-1:0] node7732;
	wire [16-1:0] node7733;
	wire [16-1:0] node7736;
	wire [16-1:0] node7739;
	wire [16-1:0] node7740;
	wire [16-1:0] node7743;
	wire [16-1:0] node7746;
	wire [16-1:0] node7747;
	wire [16-1:0] node7748;
	wire [16-1:0] node7749;
	wire [16-1:0] node7750;
	wire [16-1:0] node7753;
	wire [16-1:0] node7756;
	wire [16-1:0] node7757;
	wire [16-1:0] node7760;
	wire [16-1:0] node7763;
	wire [16-1:0] node7764;
	wire [16-1:0] node7765;
	wire [16-1:0] node7768;
	wire [16-1:0] node7771;
	wire [16-1:0] node7772;
	wire [16-1:0] node7775;
	wire [16-1:0] node7778;
	wire [16-1:0] node7779;
	wire [16-1:0] node7780;
	wire [16-1:0] node7781;
	wire [16-1:0] node7784;
	wire [16-1:0] node7787;
	wire [16-1:0] node7788;
	wire [16-1:0] node7791;
	wire [16-1:0] node7794;
	wire [16-1:0] node7795;
	wire [16-1:0] node7796;
	wire [16-1:0] node7799;
	wire [16-1:0] node7802;
	wire [16-1:0] node7803;
	wire [16-1:0] node7806;
	wire [16-1:0] node7809;
	wire [16-1:0] node7810;
	wire [16-1:0] node7811;
	wire [16-1:0] node7812;
	wire [16-1:0] node7813;
	wire [16-1:0] node7814;
	wire [16-1:0] node7817;
	wire [16-1:0] node7820;
	wire [16-1:0] node7821;
	wire [16-1:0] node7824;
	wire [16-1:0] node7827;
	wire [16-1:0] node7828;
	wire [16-1:0] node7829;
	wire [16-1:0] node7832;
	wire [16-1:0] node7835;
	wire [16-1:0] node7836;
	wire [16-1:0] node7839;
	wire [16-1:0] node7842;
	wire [16-1:0] node7843;
	wire [16-1:0] node7844;
	wire [16-1:0] node7845;
	wire [16-1:0] node7848;
	wire [16-1:0] node7851;
	wire [16-1:0] node7852;
	wire [16-1:0] node7855;
	wire [16-1:0] node7858;
	wire [16-1:0] node7859;
	wire [16-1:0] node7860;
	wire [16-1:0] node7863;
	wire [16-1:0] node7866;
	wire [16-1:0] node7867;
	wire [16-1:0] node7870;
	wire [16-1:0] node7873;
	wire [16-1:0] node7874;
	wire [16-1:0] node7875;
	wire [16-1:0] node7876;
	wire [16-1:0] node7877;
	wire [16-1:0] node7880;
	wire [16-1:0] node7883;
	wire [16-1:0] node7884;
	wire [16-1:0] node7887;
	wire [16-1:0] node7890;
	wire [16-1:0] node7891;
	wire [16-1:0] node7892;
	wire [16-1:0] node7895;
	wire [16-1:0] node7898;
	wire [16-1:0] node7899;
	wire [16-1:0] node7902;
	wire [16-1:0] node7905;
	wire [16-1:0] node7906;
	wire [16-1:0] node7907;
	wire [16-1:0] node7908;
	wire [16-1:0] node7911;
	wire [16-1:0] node7914;
	wire [16-1:0] node7915;
	wire [16-1:0] node7918;
	wire [16-1:0] node7921;
	wire [16-1:0] node7922;
	wire [16-1:0] node7923;
	wire [16-1:0] node7926;
	wire [16-1:0] node7929;
	wire [16-1:0] node7930;
	wire [16-1:0] node7933;
	wire [16-1:0] node7936;
	wire [16-1:0] node7937;
	wire [16-1:0] node7938;
	wire [16-1:0] node7939;
	wire [16-1:0] node7940;
	wire [16-1:0] node7941;
	wire [16-1:0] node7942;
	wire [16-1:0] node7945;
	wire [16-1:0] node7948;
	wire [16-1:0] node7949;
	wire [16-1:0] node7952;
	wire [16-1:0] node7955;
	wire [16-1:0] node7956;
	wire [16-1:0] node7957;
	wire [16-1:0] node7960;
	wire [16-1:0] node7963;
	wire [16-1:0] node7964;
	wire [16-1:0] node7967;
	wire [16-1:0] node7970;
	wire [16-1:0] node7971;
	wire [16-1:0] node7972;
	wire [16-1:0] node7973;
	wire [16-1:0] node7976;
	wire [16-1:0] node7979;
	wire [16-1:0] node7980;
	wire [16-1:0] node7983;
	wire [16-1:0] node7986;
	wire [16-1:0] node7987;
	wire [16-1:0] node7988;
	wire [16-1:0] node7991;
	wire [16-1:0] node7994;
	wire [16-1:0] node7995;
	wire [16-1:0] node7998;
	wire [16-1:0] node8001;
	wire [16-1:0] node8002;
	wire [16-1:0] node8003;
	wire [16-1:0] node8004;
	wire [16-1:0] node8005;
	wire [16-1:0] node8008;
	wire [16-1:0] node8011;
	wire [16-1:0] node8012;
	wire [16-1:0] node8015;
	wire [16-1:0] node8018;
	wire [16-1:0] node8019;
	wire [16-1:0] node8020;
	wire [16-1:0] node8023;
	wire [16-1:0] node8026;
	wire [16-1:0] node8027;
	wire [16-1:0] node8030;
	wire [16-1:0] node8033;
	wire [16-1:0] node8034;
	wire [16-1:0] node8035;
	wire [16-1:0] node8036;
	wire [16-1:0] node8039;
	wire [16-1:0] node8042;
	wire [16-1:0] node8043;
	wire [16-1:0] node8046;
	wire [16-1:0] node8049;
	wire [16-1:0] node8050;
	wire [16-1:0] node8051;
	wire [16-1:0] node8054;
	wire [16-1:0] node8057;
	wire [16-1:0] node8058;
	wire [16-1:0] node8061;
	wire [16-1:0] node8064;
	wire [16-1:0] node8065;
	wire [16-1:0] node8066;
	wire [16-1:0] node8067;
	wire [16-1:0] node8068;
	wire [16-1:0] node8069;
	wire [16-1:0] node8072;
	wire [16-1:0] node8075;
	wire [16-1:0] node8076;
	wire [16-1:0] node8079;
	wire [16-1:0] node8082;
	wire [16-1:0] node8083;
	wire [16-1:0] node8084;
	wire [16-1:0] node8087;
	wire [16-1:0] node8090;
	wire [16-1:0] node8091;
	wire [16-1:0] node8094;
	wire [16-1:0] node8097;
	wire [16-1:0] node8098;
	wire [16-1:0] node8099;
	wire [16-1:0] node8100;
	wire [16-1:0] node8103;
	wire [16-1:0] node8106;
	wire [16-1:0] node8107;
	wire [16-1:0] node8110;
	wire [16-1:0] node8113;
	wire [16-1:0] node8114;
	wire [16-1:0] node8115;
	wire [16-1:0] node8118;
	wire [16-1:0] node8121;
	wire [16-1:0] node8122;
	wire [16-1:0] node8125;
	wire [16-1:0] node8128;
	wire [16-1:0] node8129;
	wire [16-1:0] node8130;
	wire [16-1:0] node8131;
	wire [16-1:0] node8132;
	wire [16-1:0] node8135;
	wire [16-1:0] node8138;
	wire [16-1:0] node8139;
	wire [16-1:0] node8142;
	wire [16-1:0] node8145;
	wire [16-1:0] node8146;
	wire [16-1:0] node8147;
	wire [16-1:0] node8150;
	wire [16-1:0] node8153;
	wire [16-1:0] node8154;
	wire [16-1:0] node8157;
	wire [16-1:0] node8160;
	wire [16-1:0] node8161;
	wire [16-1:0] node8162;
	wire [16-1:0] node8163;
	wire [16-1:0] node8166;
	wire [16-1:0] node8169;
	wire [16-1:0] node8170;
	wire [16-1:0] node8173;
	wire [16-1:0] node8176;
	wire [16-1:0] node8177;
	wire [16-1:0] node8178;
	wire [16-1:0] node8181;
	wire [16-1:0] node8184;
	wire [16-1:0] node8185;
	wire [16-1:0] node8188;

	assign outp = (inp[1]) ? node4096 : node1;
		assign node1 = (inp[11]) ? node2049 : node2;
			assign node2 = (inp[3]) ? node1026 : node3;
				assign node3 = (inp[9]) ? node515 : node4;
					assign node4 = (inp[14]) ? node260 : node5;
						assign node5 = (inp[10]) ? node133 : node6;
							assign node6 = (inp[12]) ? node70 : node7;
								assign node7 = (inp[6]) ? node39 : node8;
									assign node8 = (inp[8]) ? node24 : node9;
										assign node9 = (inp[0]) ? node17 : node10;
											assign node10 = (inp[13]) ? node14 : node11;
												assign node11 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node14 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node17 = (inp[5]) ? node21 : node18;
												assign node18 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node21 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node24 = (inp[7]) ? node32 : node25;
											assign node25 = (inp[0]) ? node29 : node26;
												assign node26 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node29 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node32 = (inp[4]) ? node36 : node33;
												assign node33 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node36 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
									assign node39 = (inp[7]) ? node55 : node40;
										assign node40 = (inp[13]) ? node48 : node41;
											assign node41 = (inp[8]) ? node45 : node42;
												assign node42 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node45 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node48 = (inp[15]) ? node52 : node49;
												assign node49 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node52 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node55 = (inp[2]) ? node63 : node56;
											assign node56 = (inp[13]) ? node60 : node57;
												assign node57 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node60 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node63 = (inp[4]) ? node67 : node64;
												assign node64 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node67 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node70 = (inp[13]) ? node102 : node71;
									assign node71 = (inp[2]) ? node87 : node72;
										assign node72 = (inp[4]) ? node80 : node73;
											assign node73 = (inp[0]) ? node77 : node74;
												assign node74 = (inp[6]) ? 16'b0000111111111111 : 16'b0011111111111111;
												assign node77 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node80 = (inp[7]) ? node84 : node81;
												assign node81 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node84 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node87 = (inp[8]) ? node95 : node88;
											assign node88 = (inp[15]) ? node92 : node89;
												assign node89 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node92 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node95 = (inp[7]) ? node99 : node96;
												assign node96 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node99 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node102 = (inp[2]) ? node118 : node103;
										assign node103 = (inp[0]) ? node111 : node104;
											assign node104 = (inp[7]) ? node108 : node105;
												assign node105 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node108 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node111 = (inp[8]) ? node115 : node112;
												assign node112 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node115 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node118 = (inp[6]) ? node126 : node119;
											assign node119 = (inp[4]) ? node123 : node120;
												assign node120 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node123 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node126 = (inp[0]) ? node130 : node127;
												assign node127 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node130 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
							assign node133 = (inp[0]) ? node197 : node134;
								assign node134 = (inp[13]) ? node166 : node135;
									assign node135 = (inp[5]) ? node151 : node136;
										assign node136 = (inp[4]) ? node144 : node137;
											assign node137 = (inp[8]) ? node141 : node138;
												assign node138 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node141 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node144 = (inp[2]) ? node148 : node145;
												assign node145 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node148 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node151 = (inp[8]) ? node159 : node152;
											assign node152 = (inp[12]) ? node156 : node153;
												assign node153 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node156 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node159 = (inp[2]) ? node163 : node160;
												assign node160 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node163 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node166 = (inp[2]) ? node182 : node167;
										assign node167 = (inp[7]) ? node175 : node168;
											assign node168 = (inp[12]) ? node172 : node169;
												assign node169 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node172 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node175 = (inp[4]) ? node179 : node176;
												assign node176 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node179 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node182 = (inp[5]) ? node190 : node183;
											assign node183 = (inp[8]) ? node187 : node184;
												assign node184 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node187 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node190 = (inp[6]) ? node194 : node191;
												assign node191 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node194 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node197 = (inp[7]) ? node229 : node198;
									assign node198 = (inp[15]) ? node214 : node199;
										assign node199 = (inp[13]) ? node207 : node200;
											assign node200 = (inp[6]) ? node204 : node201;
												assign node201 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node204 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node207 = (inp[6]) ? node211 : node208;
												assign node208 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node211 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node214 = (inp[12]) ? node222 : node215;
											assign node215 = (inp[6]) ? node219 : node216;
												assign node216 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node219 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node222 = (inp[8]) ? node226 : node223;
												assign node223 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node226 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node229 = (inp[4]) ? node245 : node230;
										assign node230 = (inp[2]) ? node238 : node231;
											assign node231 = (inp[6]) ? node235 : node232;
												assign node232 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node235 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node238 = (inp[5]) ? node242 : node239;
												assign node239 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node242 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node245 = (inp[13]) ? node253 : node246;
											assign node246 = (inp[6]) ? node250 : node247;
												assign node247 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node250 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node253 = (inp[5]) ? node257 : node254;
												assign node254 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node257 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node260 = (inp[6]) ? node388 : node261;
							assign node261 = (inp[5]) ? node325 : node262;
								assign node262 = (inp[7]) ? node294 : node263;
									assign node263 = (inp[4]) ? node279 : node264;
										assign node264 = (inp[12]) ? node272 : node265;
											assign node265 = (inp[13]) ? node269 : node266;
												assign node266 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node269 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node272 = (inp[8]) ? node276 : node273;
												assign node273 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node276 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node279 = (inp[10]) ? node287 : node280;
											assign node280 = (inp[2]) ? node284 : node281;
												assign node281 = (inp[8]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node284 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node287 = (inp[12]) ? node291 : node288;
												assign node288 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node291 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node294 = (inp[8]) ? node310 : node295;
										assign node295 = (inp[0]) ? node303 : node296;
											assign node296 = (inp[15]) ? node300 : node297;
												assign node297 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node300 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node303 = (inp[2]) ? node307 : node304;
												assign node304 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node307 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node310 = (inp[2]) ? node318 : node311;
											assign node311 = (inp[4]) ? node315 : node312;
												assign node312 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node315 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node318 = (inp[10]) ? node322 : node319;
												assign node319 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node322 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node325 = (inp[2]) ? node357 : node326;
									assign node326 = (inp[13]) ? node342 : node327;
										assign node327 = (inp[15]) ? node335 : node328;
											assign node328 = (inp[10]) ? node332 : node329;
												assign node329 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node332 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node335 = (inp[0]) ? node339 : node336;
												assign node336 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node339 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node342 = (inp[8]) ? node350 : node343;
											assign node343 = (inp[15]) ? node347 : node344;
												assign node344 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node347 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node350 = (inp[12]) ? node354 : node351;
												assign node351 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node354 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node357 = (inp[4]) ? node373 : node358;
										assign node358 = (inp[10]) ? node366 : node359;
											assign node359 = (inp[12]) ? node363 : node360;
												assign node360 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node363 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node366 = (inp[13]) ? node370 : node367;
												assign node367 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node370 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node373 = (inp[0]) ? node381 : node374;
											assign node374 = (inp[7]) ? node378 : node375;
												assign node375 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node378 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node381 = (inp[8]) ? node385 : node382;
												assign node382 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node385 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node388 = (inp[10]) ? node452 : node389;
								assign node389 = (inp[8]) ? node421 : node390;
									assign node390 = (inp[5]) ? node406 : node391;
										assign node391 = (inp[15]) ? node399 : node392;
											assign node392 = (inp[0]) ? node396 : node393;
												assign node393 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node396 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node399 = (inp[4]) ? node403 : node400;
												assign node400 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node403 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node406 = (inp[4]) ? node414 : node407;
											assign node407 = (inp[7]) ? node411 : node408;
												assign node408 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node411 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node414 = (inp[2]) ? node418 : node415;
												assign node415 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node418 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node421 = (inp[13]) ? node437 : node422;
										assign node422 = (inp[12]) ? node430 : node423;
											assign node423 = (inp[0]) ? node427 : node424;
												assign node424 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node427 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node430 = (inp[15]) ? node434 : node431;
												assign node431 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node434 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node437 = (inp[7]) ? node445 : node438;
											assign node438 = (inp[0]) ? node442 : node439;
												assign node439 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node442 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node445 = (inp[5]) ? node449 : node446;
												assign node446 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node449 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node452 = (inp[12]) ? node484 : node453;
									assign node453 = (inp[0]) ? node469 : node454;
										assign node454 = (inp[4]) ? node462 : node455;
											assign node455 = (inp[7]) ? node459 : node456;
												assign node456 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node459 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node462 = (inp[15]) ? node466 : node463;
												assign node463 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node466 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node469 = (inp[8]) ? node477 : node470;
											assign node470 = (inp[2]) ? node474 : node471;
												assign node471 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node474 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node477 = (inp[5]) ? node481 : node478;
												assign node478 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node481 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node484 = (inp[15]) ? node500 : node485;
										assign node485 = (inp[4]) ? node493 : node486;
											assign node486 = (inp[13]) ? node490 : node487;
												assign node487 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node490 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node493 = (inp[5]) ? node497 : node494;
												assign node494 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node497 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node500 = (inp[2]) ? node508 : node501;
											assign node501 = (inp[7]) ? node505 : node502;
												assign node502 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node505 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node508 = (inp[0]) ? node512 : node509;
												assign node509 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node512 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node515 = (inp[4]) ? node771 : node516;
						assign node516 = (inp[5]) ? node644 : node517;
							assign node517 = (inp[0]) ? node581 : node518;
								assign node518 = (inp[2]) ? node550 : node519;
									assign node519 = (inp[15]) ? node535 : node520;
										assign node520 = (inp[6]) ? node528 : node521;
											assign node521 = (inp[8]) ? node525 : node522;
												assign node522 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node525 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node528 = (inp[7]) ? node532 : node529;
												assign node529 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node532 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node535 = (inp[14]) ? node543 : node536;
											assign node536 = (inp[7]) ? node540 : node537;
												assign node537 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node540 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node543 = (inp[6]) ? node547 : node544;
												assign node544 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node547 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node550 = (inp[15]) ? node566 : node551;
										assign node551 = (inp[8]) ? node559 : node552;
											assign node552 = (inp[12]) ? node556 : node553;
												assign node553 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node556 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node559 = (inp[13]) ? node563 : node560;
												assign node560 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node563 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node566 = (inp[13]) ? node574 : node567;
											assign node567 = (inp[7]) ? node571 : node568;
												assign node568 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node571 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node574 = (inp[8]) ? node578 : node575;
												assign node575 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node578 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node581 = (inp[7]) ? node613 : node582;
									assign node582 = (inp[13]) ? node598 : node583;
										assign node583 = (inp[6]) ? node591 : node584;
											assign node584 = (inp[2]) ? node588 : node585;
												assign node585 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node588 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node591 = (inp[8]) ? node595 : node592;
												assign node592 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node595 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node598 = (inp[12]) ? node606 : node599;
											assign node599 = (inp[6]) ? node603 : node600;
												assign node600 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node603 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node606 = (inp[8]) ? node610 : node607;
												assign node607 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node610 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node613 = (inp[2]) ? node629 : node614;
										assign node614 = (inp[8]) ? node622 : node615;
											assign node615 = (inp[13]) ? node619 : node616;
												assign node616 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node619 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node622 = (inp[10]) ? node626 : node623;
												assign node623 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node626 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node629 = (inp[15]) ? node637 : node630;
											assign node630 = (inp[10]) ? node634 : node631;
												assign node631 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node634 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node637 = (inp[13]) ? node641 : node638;
												assign node638 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node641 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
							assign node644 = (inp[2]) ? node708 : node645;
								assign node645 = (inp[7]) ? node677 : node646;
									assign node646 = (inp[12]) ? node662 : node647;
										assign node647 = (inp[6]) ? node655 : node648;
											assign node648 = (inp[10]) ? node652 : node649;
												assign node649 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node652 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node655 = (inp[13]) ? node659 : node656;
												assign node656 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node659 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node662 = (inp[13]) ? node670 : node663;
											assign node663 = (inp[8]) ? node667 : node664;
												assign node664 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node667 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node670 = (inp[6]) ? node674 : node671;
												assign node671 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node674 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node677 = (inp[12]) ? node693 : node678;
										assign node678 = (inp[14]) ? node686 : node679;
											assign node679 = (inp[15]) ? node683 : node680;
												assign node680 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node683 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node686 = (inp[10]) ? node690 : node687;
												assign node687 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node690 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node693 = (inp[13]) ? node701 : node694;
											assign node694 = (inp[6]) ? node698 : node695;
												assign node695 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node698 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node701 = (inp[10]) ? node705 : node702;
												assign node702 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node705 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node708 = (inp[8]) ? node740 : node709;
									assign node709 = (inp[6]) ? node725 : node710;
										assign node710 = (inp[13]) ? node718 : node711;
											assign node711 = (inp[10]) ? node715 : node712;
												assign node712 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node715 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node718 = (inp[7]) ? node722 : node719;
												assign node719 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node722 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node725 = (inp[14]) ? node733 : node726;
											assign node726 = (inp[12]) ? node730 : node727;
												assign node727 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node730 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node733 = (inp[10]) ? node737 : node734;
												assign node734 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node737 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node740 = (inp[12]) ? node756 : node741;
										assign node741 = (inp[7]) ? node749 : node742;
											assign node742 = (inp[13]) ? node746 : node743;
												assign node743 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node746 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node749 = (inp[15]) ? node753 : node750;
												assign node750 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node753 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node756 = (inp[6]) ? node764 : node757;
											assign node757 = (inp[0]) ? node761 : node758;
												assign node758 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node761 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node764 = (inp[0]) ? node768 : node765;
												assign node765 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node768 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
						assign node771 = (inp[12]) ? node899 : node772;
							assign node772 = (inp[15]) ? node836 : node773;
								assign node773 = (inp[13]) ? node805 : node774;
									assign node774 = (inp[14]) ? node790 : node775;
										assign node775 = (inp[6]) ? node783 : node776;
											assign node776 = (inp[0]) ? node780 : node777;
												assign node777 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node780 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node783 = (inp[0]) ? node787 : node784;
												assign node784 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node787 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node790 = (inp[8]) ? node798 : node791;
											assign node791 = (inp[7]) ? node795 : node792;
												assign node792 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node795 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node798 = (inp[2]) ? node802 : node799;
												assign node799 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node802 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node805 = (inp[10]) ? node821 : node806;
										assign node806 = (inp[14]) ? node814 : node807;
											assign node807 = (inp[6]) ? node811 : node808;
												assign node808 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node811 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node814 = (inp[8]) ? node818 : node815;
												assign node815 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node818 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node821 = (inp[0]) ? node829 : node822;
											assign node822 = (inp[5]) ? node826 : node823;
												assign node823 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node826 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node829 = (inp[8]) ? node833 : node830;
												assign node830 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node833 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node836 = (inp[0]) ? node868 : node837;
									assign node837 = (inp[13]) ? node853 : node838;
										assign node838 = (inp[7]) ? node846 : node839;
											assign node839 = (inp[2]) ? node843 : node840;
												assign node840 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node843 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node846 = (inp[14]) ? node850 : node847;
												assign node847 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node850 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node853 = (inp[10]) ? node861 : node854;
											assign node854 = (inp[7]) ? node858 : node855;
												assign node855 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node858 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node861 = (inp[14]) ? node865 : node862;
												assign node862 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node865 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node868 = (inp[2]) ? node884 : node869;
										assign node869 = (inp[6]) ? node877 : node870;
											assign node870 = (inp[7]) ? node874 : node871;
												assign node871 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node874 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node877 = (inp[13]) ? node881 : node878;
												assign node878 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node881 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node884 = (inp[5]) ? node892 : node885;
											assign node885 = (inp[8]) ? node889 : node886;
												assign node886 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node889 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node892 = (inp[10]) ? node896 : node893;
												assign node893 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node896 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node899 = (inp[6]) ? node963 : node900;
								assign node900 = (inp[15]) ? node932 : node901;
									assign node901 = (inp[13]) ? node917 : node902;
										assign node902 = (inp[5]) ? node910 : node903;
											assign node903 = (inp[8]) ? node907 : node904;
												assign node904 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node907 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node910 = (inp[7]) ? node914 : node911;
												assign node911 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node914 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node917 = (inp[10]) ? node925 : node918;
											assign node918 = (inp[14]) ? node922 : node919;
												assign node919 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node922 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node925 = (inp[7]) ? node929 : node926;
												assign node926 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node929 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node932 = (inp[0]) ? node948 : node933;
										assign node933 = (inp[2]) ? node941 : node934;
											assign node934 = (inp[13]) ? node938 : node935;
												assign node935 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node938 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node941 = (inp[10]) ? node945 : node942;
												assign node942 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node945 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node948 = (inp[5]) ? node956 : node949;
											assign node949 = (inp[8]) ? node953 : node950;
												assign node950 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node953 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node956 = (inp[7]) ? node960 : node957;
												assign node957 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node960 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node963 = (inp[13]) ? node995 : node964;
									assign node964 = (inp[0]) ? node980 : node965;
										assign node965 = (inp[7]) ? node973 : node966;
											assign node966 = (inp[5]) ? node970 : node967;
												assign node967 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node970 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node973 = (inp[14]) ? node977 : node974;
												assign node974 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node977 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node980 = (inp[15]) ? node988 : node981;
											assign node981 = (inp[8]) ? node985 : node982;
												assign node982 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node985 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node988 = (inp[14]) ? node992 : node989;
												assign node989 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node992 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node995 = (inp[5]) ? node1011 : node996;
										assign node996 = (inp[7]) ? node1004 : node997;
											assign node997 = (inp[0]) ? node1001 : node998;
												assign node998 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1001 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1004 = (inp[8]) ? node1008 : node1005;
												assign node1005 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1008 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1011 = (inp[0]) ? node1019 : node1012;
											assign node1012 = (inp[15]) ? node1016 : node1013;
												assign node1013 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1016 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1019 = (inp[10]) ? node1023 : node1020;
												assign node1020 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1023 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
				assign node1026 = (inp[8]) ? node1538 : node1027;
					assign node1027 = (inp[0]) ? node1283 : node1028;
						assign node1028 = (inp[9]) ? node1156 : node1029;
							assign node1029 = (inp[13]) ? node1093 : node1030;
								assign node1030 = (inp[2]) ? node1062 : node1031;
									assign node1031 = (inp[12]) ? node1047 : node1032;
										assign node1032 = (inp[10]) ? node1040 : node1033;
											assign node1033 = (inp[14]) ? node1037 : node1034;
												assign node1034 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node1037 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1040 = (inp[5]) ? node1044 : node1041;
												assign node1041 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1044 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1047 = (inp[14]) ? node1055 : node1048;
											assign node1048 = (inp[5]) ? node1052 : node1049;
												assign node1049 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1052 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1055 = (inp[6]) ? node1059 : node1056;
												assign node1056 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1059 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1062 = (inp[12]) ? node1078 : node1063;
										assign node1063 = (inp[6]) ? node1071 : node1064;
											assign node1064 = (inp[5]) ? node1068 : node1065;
												assign node1065 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1068 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1071 = (inp[5]) ? node1075 : node1072;
												assign node1072 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1075 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1078 = (inp[14]) ? node1086 : node1079;
											assign node1079 = (inp[6]) ? node1083 : node1080;
												assign node1080 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1083 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1086 = (inp[10]) ? node1090 : node1087;
												assign node1087 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1090 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1093 = (inp[7]) ? node1125 : node1094;
									assign node1094 = (inp[4]) ? node1110 : node1095;
										assign node1095 = (inp[2]) ? node1103 : node1096;
											assign node1096 = (inp[12]) ? node1100 : node1097;
												assign node1097 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1100 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1103 = (inp[15]) ? node1107 : node1104;
												assign node1104 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1107 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1110 = (inp[6]) ? node1118 : node1111;
											assign node1111 = (inp[2]) ? node1115 : node1112;
												assign node1112 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1115 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1118 = (inp[14]) ? node1122 : node1119;
												assign node1119 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1122 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1125 = (inp[6]) ? node1141 : node1126;
										assign node1126 = (inp[14]) ? node1134 : node1127;
											assign node1127 = (inp[15]) ? node1131 : node1128;
												assign node1128 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1131 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1134 = (inp[4]) ? node1138 : node1135;
												assign node1135 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1138 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1141 = (inp[12]) ? node1149 : node1142;
											assign node1142 = (inp[5]) ? node1146 : node1143;
												assign node1143 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1146 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1149 = (inp[2]) ? node1153 : node1150;
												assign node1150 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1153 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1156 = (inp[2]) ? node1220 : node1157;
								assign node1157 = (inp[15]) ? node1189 : node1158;
									assign node1158 = (inp[13]) ? node1174 : node1159;
										assign node1159 = (inp[14]) ? node1167 : node1160;
											assign node1160 = (inp[7]) ? node1164 : node1161;
												assign node1161 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1164 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1167 = (inp[5]) ? node1171 : node1168;
												assign node1168 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1171 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1174 = (inp[14]) ? node1182 : node1175;
											assign node1175 = (inp[6]) ? node1179 : node1176;
												assign node1176 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1179 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1182 = (inp[7]) ? node1186 : node1183;
												assign node1183 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1186 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1189 = (inp[4]) ? node1205 : node1190;
										assign node1190 = (inp[13]) ? node1198 : node1191;
											assign node1191 = (inp[5]) ? node1195 : node1192;
												assign node1192 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1195 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1198 = (inp[7]) ? node1202 : node1199;
												assign node1199 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1202 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1205 = (inp[6]) ? node1213 : node1206;
											assign node1206 = (inp[10]) ? node1210 : node1207;
												assign node1207 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1210 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1213 = (inp[5]) ? node1217 : node1214;
												assign node1214 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1217 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1220 = (inp[5]) ? node1252 : node1221;
									assign node1221 = (inp[14]) ? node1237 : node1222;
										assign node1222 = (inp[12]) ? node1230 : node1223;
											assign node1223 = (inp[4]) ? node1227 : node1224;
												assign node1224 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1227 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1230 = (inp[10]) ? node1234 : node1231;
												assign node1231 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1234 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1237 = (inp[7]) ? node1245 : node1238;
											assign node1238 = (inp[10]) ? node1242 : node1239;
												assign node1239 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1242 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1245 = (inp[12]) ? node1249 : node1246;
												assign node1246 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1249 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1252 = (inp[6]) ? node1268 : node1253;
										assign node1253 = (inp[10]) ? node1261 : node1254;
											assign node1254 = (inp[13]) ? node1258 : node1255;
												assign node1255 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1258 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1261 = (inp[4]) ? node1265 : node1262;
												assign node1262 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1265 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1268 = (inp[10]) ? node1276 : node1269;
											assign node1269 = (inp[15]) ? node1273 : node1270;
												assign node1270 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1273 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1276 = (inp[13]) ? node1280 : node1277;
												assign node1277 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1280 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node1283 = (inp[4]) ? node1411 : node1284;
							assign node1284 = (inp[13]) ? node1348 : node1285;
								assign node1285 = (inp[2]) ? node1317 : node1286;
									assign node1286 = (inp[15]) ? node1302 : node1287;
										assign node1287 = (inp[12]) ? node1295 : node1288;
											assign node1288 = (inp[7]) ? node1292 : node1289;
												assign node1289 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1292 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1295 = (inp[6]) ? node1299 : node1296;
												assign node1296 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1299 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1302 = (inp[6]) ? node1310 : node1303;
											assign node1303 = (inp[12]) ? node1307 : node1304;
												assign node1304 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1307 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1310 = (inp[10]) ? node1314 : node1311;
												assign node1311 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1314 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1317 = (inp[14]) ? node1333 : node1318;
										assign node1318 = (inp[6]) ? node1326 : node1319;
											assign node1319 = (inp[10]) ? node1323 : node1320;
												assign node1320 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1323 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1326 = (inp[12]) ? node1330 : node1327;
												assign node1327 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1330 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1333 = (inp[10]) ? node1341 : node1334;
											assign node1334 = (inp[9]) ? node1338 : node1335;
												assign node1335 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1338 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1341 = (inp[15]) ? node1345 : node1342;
												assign node1342 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1345 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1348 = (inp[5]) ? node1380 : node1349;
									assign node1349 = (inp[14]) ? node1365 : node1350;
										assign node1350 = (inp[12]) ? node1358 : node1351;
											assign node1351 = (inp[10]) ? node1355 : node1352;
												assign node1352 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1355 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1358 = (inp[7]) ? node1362 : node1359;
												assign node1359 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1362 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1365 = (inp[10]) ? node1373 : node1366;
											assign node1366 = (inp[9]) ? node1370 : node1367;
												assign node1367 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1370 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1373 = (inp[15]) ? node1377 : node1374;
												assign node1374 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1377 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1380 = (inp[9]) ? node1396 : node1381;
										assign node1381 = (inp[12]) ? node1389 : node1382;
											assign node1382 = (inp[10]) ? node1386 : node1383;
												assign node1383 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1386 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1389 = (inp[7]) ? node1393 : node1390;
												assign node1390 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1393 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1396 = (inp[2]) ? node1404 : node1397;
											assign node1397 = (inp[12]) ? node1401 : node1398;
												assign node1398 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1401 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1404 = (inp[15]) ? node1408 : node1405;
												assign node1405 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node1408 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1411 = (inp[10]) ? node1475 : node1412;
								assign node1412 = (inp[12]) ? node1444 : node1413;
									assign node1413 = (inp[15]) ? node1429 : node1414;
										assign node1414 = (inp[5]) ? node1422 : node1415;
											assign node1415 = (inp[7]) ? node1419 : node1416;
												assign node1416 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1419 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1422 = (inp[6]) ? node1426 : node1423;
												assign node1423 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1426 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1429 = (inp[14]) ? node1437 : node1430;
											assign node1430 = (inp[2]) ? node1434 : node1431;
												assign node1431 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1434 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1437 = (inp[9]) ? node1441 : node1438;
												assign node1438 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1441 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1444 = (inp[13]) ? node1460 : node1445;
										assign node1445 = (inp[9]) ? node1453 : node1446;
											assign node1446 = (inp[14]) ? node1450 : node1447;
												assign node1447 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1450 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1453 = (inp[7]) ? node1457 : node1454;
												assign node1454 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1457 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1460 = (inp[2]) ? node1468 : node1461;
											assign node1461 = (inp[5]) ? node1465 : node1462;
												assign node1462 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1465 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1468 = (inp[15]) ? node1472 : node1469;
												assign node1469 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1472 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1475 = (inp[14]) ? node1507 : node1476;
									assign node1476 = (inp[7]) ? node1492 : node1477;
										assign node1477 = (inp[15]) ? node1485 : node1478;
											assign node1478 = (inp[12]) ? node1482 : node1479;
												assign node1479 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1482 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1485 = (inp[2]) ? node1489 : node1486;
												assign node1486 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1489 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1492 = (inp[13]) ? node1500 : node1493;
											assign node1493 = (inp[5]) ? node1497 : node1494;
												assign node1494 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1497 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1500 = (inp[9]) ? node1504 : node1501;
												assign node1501 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1504 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1507 = (inp[9]) ? node1523 : node1508;
										assign node1508 = (inp[12]) ? node1516 : node1509;
											assign node1509 = (inp[15]) ? node1513 : node1510;
												assign node1510 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1513 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1516 = (inp[5]) ? node1520 : node1517;
												assign node1517 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1520 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1523 = (inp[15]) ? node1531 : node1524;
											assign node1524 = (inp[7]) ? node1528 : node1525;
												assign node1525 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1528 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1531 = (inp[6]) ? node1535 : node1532;
												assign node1532 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1535 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node1538 = (inp[2]) ? node1794 : node1539;
						assign node1539 = (inp[14]) ? node1667 : node1540;
							assign node1540 = (inp[4]) ? node1604 : node1541;
								assign node1541 = (inp[6]) ? node1573 : node1542;
									assign node1542 = (inp[12]) ? node1558 : node1543;
										assign node1543 = (inp[7]) ? node1551 : node1544;
											assign node1544 = (inp[9]) ? node1548 : node1545;
												assign node1545 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1548 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1551 = (inp[13]) ? node1555 : node1552;
												assign node1552 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1555 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1558 = (inp[0]) ? node1566 : node1559;
											assign node1559 = (inp[7]) ? node1563 : node1560;
												assign node1560 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1563 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1566 = (inp[10]) ? node1570 : node1567;
												assign node1567 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1570 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1573 = (inp[9]) ? node1589 : node1574;
										assign node1574 = (inp[7]) ? node1582 : node1575;
											assign node1575 = (inp[15]) ? node1579 : node1576;
												assign node1576 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1579 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1582 = (inp[0]) ? node1586 : node1583;
												assign node1583 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1586 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1589 = (inp[13]) ? node1597 : node1590;
											assign node1590 = (inp[10]) ? node1594 : node1591;
												assign node1591 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1594 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1597 = (inp[12]) ? node1601 : node1598;
												assign node1598 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1601 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1604 = (inp[9]) ? node1636 : node1605;
									assign node1605 = (inp[10]) ? node1621 : node1606;
										assign node1606 = (inp[6]) ? node1614 : node1607;
											assign node1607 = (inp[13]) ? node1611 : node1608;
												assign node1608 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1611 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1614 = (inp[0]) ? node1618 : node1615;
												assign node1615 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1618 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1621 = (inp[15]) ? node1629 : node1622;
											assign node1622 = (inp[0]) ? node1626 : node1623;
												assign node1623 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1626 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1629 = (inp[12]) ? node1633 : node1630;
												assign node1630 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1633 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1636 = (inp[6]) ? node1652 : node1637;
										assign node1637 = (inp[12]) ? node1645 : node1638;
											assign node1638 = (inp[0]) ? node1642 : node1639;
												assign node1639 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1642 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1645 = (inp[15]) ? node1649 : node1646;
												assign node1646 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1649 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1652 = (inp[7]) ? node1660 : node1653;
											assign node1653 = (inp[10]) ? node1657 : node1654;
												assign node1654 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1657 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node1660 = (inp[0]) ? node1664 : node1661;
												assign node1661 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1664 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1667 = (inp[12]) ? node1731 : node1668;
								assign node1668 = (inp[5]) ? node1700 : node1669;
									assign node1669 = (inp[15]) ? node1685 : node1670;
										assign node1670 = (inp[9]) ? node1678 : node1671;
											assign node1671 = (inp[0]) ? node1675 : node1672;
												assign node1672 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1675 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1678 = (inp[7]) ? node1682 : node1679;
												assign node1679 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1682 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1685 = (inp[4]) ? node1693 : node1686;
											assign node1686 = (inp[0]) ? node1690 : node1687;
												assign node1687 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1690 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1693 = (inp[7]) ? node1697 : node1694;
												assign node1694 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1697 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1700 = (inp[13]) ? node1716 : node1701;
										assign node1701 = (inp[4]) ? node1709 : node1702;
											assign node1702 = (inp[0]) ? node1706 : node1703;
												assign node1703 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1706 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1709 = (inp[15]) ? node1713 : node1710;
												assign node1710 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1713 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1716 = (inp[15]) ? node1724 : node1717;
											assign node1717 = (inp[4]) ? node1721 : node1718;
												assign node1718 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1721 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1724 = (inp[9]) ? node1728 : node1725;
												assign node1725 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1728 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1731 = (inp[7]) ? node1763 : node1732;
									assign node1732 = (inp[4]) ? node1748 : node1733;
										assign node1733 = (inp[13]) ? node1741 : node1734;
											assign node1734 = (inp[0]) ? node1738 : node1735;
												assign node1735 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1738 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1741 = (inp[15]) ? node1745 : node1742;
												assign node1742 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1745 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1748 = (inp[6]) ? node1756 : node1749;
											assign node1749 = (inp[9]) ? node1753 : node1750;
												assign node1750 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1753 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1756 = (inp[15]) ? node1760 : node1757;
												assign node1757 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1760 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1763 = (inp[10]) ? node1779 : node1764;
										assign node1764 = (inp[13]) ? node1772 : node1765;
											assign node1765 = (inp[9]) ? node1769 : node1766;
												assign node1766 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1769 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1772 = (inp[15]) ? node1776 : node1773;
												assign node1773 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1776 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1779 = (inp[9]) ? node1787 : node1780;
											assign node1780 = (inp[0]) ? node1784 : node1781;
												assign node1781 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1784 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1787 = (inp[13]) ? node1791 : node1788;
												assign node1788 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1791 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1794 = (inp[9]) ? node1922 : node1795;
							assign node1795 = (inp[10]) ? node1859 : node1796;
								assign node1796 = (inp[13]) ? node1828 : node1797;
									assign node1797 = (inp[0]) ? node1813 : node1798;
										assign node1798 = (inp[7]) ? node1806 : node1799;
											assign node1799 = (inp[6]) ? node1803 : node1800;
												assign node1800 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1803 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1806 = (inp[5]) ? node1810 : node1807;
												assign node1807 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1810 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1813 = (inp[12]) ? node1821 : node1814;
											assign node1814 = (inp[5]) ? node1818 : node1815;
												assign node1815 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1818 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1821 = (inp[4]) ? node1825 : node1822;
												assign node1822 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1825 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1828 = (inp[7]) ? node1844 : node1829;
										assign node1829 = (inp[14]) ? node1837 : node1830;
											assign node1830 = (inp[4]) ? node1834 : node1831;
												assign node1831 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1834 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1837 = (inp[15]) ? node1841 : node1838;
												assign node1838 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1841 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1844 = (inp[4]) ? node1852 : node1845;
											assign node1845 = (inp[5]) ? node1849 : node1846;
												assign node1846 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1849 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1852 = (inp[0]) ? node1856 : node1853;
												assign node1853 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1856 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1859 = (inp[12]) ? node1891 : node1860;
									assign node1860 = (inp[7]) ? node1876 : node1861;
										assign node1861 = (inp[0]) ? node1869 : node1862;
											assign node1862 = (inp[14]) ? node1866 : node1863;
												assign node1863 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1866 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1869 = (inp[5]) ? node1873 : node1870;
												assign node1870 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1873 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1876 = (inp[4]) ? node1884 : node1877;
											assign node1877 = (inp[14]) ? node1881 : node1878;
												assign node1878 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1881 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1884 = (inp[5]) ? node1888 : node1885;
												assign node1885 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1888 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1891 = (inp[0]) ? node1907 : node1892;
										assign node1892 = (inp[15]) ? node1900 : node1893;
											assign node1893 = (inp[6]) ? node1897 : node1894;
												assign node1894 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node1897 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1900 = (inp[4]) ? node1904 : node1901;
												assign node1901 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1904 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1907 = (inp[6]) ? node1915 : node1908;
											assign node1908 = (inp[4]) ? node1912 : node1909;
												assign node1909 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1912 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1915 = (inp[4]) ? node1919 : node1916;
												assign node1916 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1919 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1922 = (inp[5]) ? node1986 : node1923;
								assign node1923 = (inp[15]) ? node1955 : node1924;
									assign node1924 = (inp[10]) ? node1940 : node1925;
										assign node1925 = (inp[7]) ? node1933 : node1926;
											assign node1926 = (inp[14]) ? node1930 : node1927;
												assign node1927 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1930 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1933 = (inp[13]) ? node1937 : node1934;
												assign node1934 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1937 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node1940 = (inp[6]) ? node1948 : node1941;
											assign node1941 = (inp[4]) ? node1945 : node1942;
												assign node1942 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1945 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1948 = (inp[14]) ? node1952 : node1949;
												assign node1949 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1952 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1955 = (inp[12]) ? node1971 : node1956;
										assign node1956 = (inp[6]) ? node1964 : node1957;
											assign node1957 = (inp[13]) ? node1961 : node1958;
												assign node1958 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1961 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1964 = (inp[14]) ? node1968 : node1965;
												assign node1965 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1968 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1971 = (inp[7]) ? node1979 : node1972;
											assign node1972 = (inp[0]) ? node1976 : node1973;
												assign node1973 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1976 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node1979 = (inp[14]) ? node1983 : node1980;
												assign node1980 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1983 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node1986 = (inp[6]) ? node2018 : node1987;
									assign node1987 = (inp[7]) ? node2003 : node1988;
										assign node1988 = (inp[13]) ? node1996 : node1989;
											assign node1989 = (inp[12]) ? node1993 : node1990;
												assign node1990 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1993 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1996 = (inp[4]) ? node2000 : node1997;
												assign node1997 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2000 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2003 = (inp[10]) ? node2011 : node2004;
											assign node2004 = (inp[15]) ? node2008 : node2005;
												assign node2005 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2008 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2011 = (inp[15]) ? node2015 : node2012;
												assign node2012 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2015 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2018 = (inp[14]) ? node2034 : node2019;
										assign node2019 = (inp[13]) ? node2027 : node2020;
											assign node2020 = (inp[10]) ? node2024 : node2021;
												assign node2021 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2024 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2027 = (inp[12]) ? node2031 : node2028;
												assign node2028 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2031 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node2034 = (inp[13]) ? node2042 : node2035;
											assign node2035 = (inp[4]) ? node2039 : node2036;
												assign node2036 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2039 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node2042 = (inp[15]) ? node2046 : node2043;
												assign node2043 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node2046 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
			assign node2049 = (inp[3]) ? node3073 : node2050;
				assign node2050 = (inp[13]) ? node2562 : node2051;
					assign node2051 = (inp[2]) ? node2307 : node2052;
						assign node2052 = (inp[6]) ? node2180 : node2053;
							assign node2053 = (inp[15]) ? node2117 : node2054;
								assign node2054 = (inp[7]) ? node2086 : node2055;
									assign node2055 = (inp[9]) ? node2071 : node2056;
										assign node2056 = (inp[5]) ? node2064 : node2057;
											assign node2057 = (inp[10]) ? node2061 : node2058;
												assign node2058 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node2061 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node2064 = (inp[14]) ? node2068 : node2065;
												assign node2065 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2068 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2071 = (inp[14]) ? node2079 : node2072;
											assign node2072 = (inp[8]) ? node2076 : node2073;
												assign node2073 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2076 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2079 = (inp[10]) ? node2083 : node2080;
												assign node2080 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node2083 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node2086 = (inp[14]) ? node2102 : node2087;
										assign node2087 = (inp[0]) ? node2095 : node2088;
											assign node2088 = (inp[10]) ? node2092 : node2089;
												assign node2089 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2092 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2095 = (inp[8]) ? node2099 : node2096;
												assign node2096 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2099 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2102 = (inp[9]) ? node2110 : node2103;
											assign node2103 = (inp[10]) ? node2107 : node2104;
												assign node2104 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2107 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2110 = (inp[4]) ? node2114 : node2111;
												assign node2111 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2114 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node2117 = (inp[12]) ? node2149 : node2118;
									assign node2118 = (inp[10]) ? node2134 : node2119;
										assign node2119 = (inp[8]) ? node2127 : node2120;
											assign node2120 = (inp[4]) ? node2124 : node2121;
												assign node2121 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2124 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2127 = (inp[9]) ? node2131 : node2128;
												assign node2128 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2131 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2134 = (inp[0]) ? node2142 : node2135;
											assign node2135 = (inp[7]) ? node2139 : node2136;
												assign node2136 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2139 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2142 = (inp[14]) ? node2146 : node2143;
												assign node2143 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2146 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2149 = (inp[0]) ? node2165 : node2150;
										assign node2150 = (inp[9]) ? node2158 : node2151;
											assign node2151 = (inp[5]) ? node2155 : node2152;
												assign node2152 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2155 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2158 = (inp[4]) ? node2162 : node2159;
												assign node2159 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2162 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2165 = (inp[5]) ? node2173 : node2166;
											assign node2166 = (inp[10]) ? node2170 : node2167;
												assign node2167 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2170 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2173 = (inp[10]) ? node2177 : node2174;
												assign node2174 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2177 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node2180 = (inp[8]) ? node2244 : node2181;
								assign node2181 = (inp[5]) ? node2213 : node2182;
									assign node2182 = (inp[10]) ? node2198 : node2183;
										assign node2183 = (inp[12]) ? node2191 : node2184;
											assign node2184 = (inp[15]) ? node2188 : node2185;
												assign node2185 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2188 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2191 = (inp[7]) ? node2195 : node2192;
												assign node2192 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2195 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2198 = (inp[7]) ? node2206 : node2199;
											assign node2199 = (inp[0]) ? node2203 : node2200;
												assign node2200 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2203 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2206 = (inp[12]) ? node2210 : node2207;
												assign node2207 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2210 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2213 = (inp[10]) ? node2229 : node2214;
										assign node2214 = (inp[4]) ? node2222 : node2215;
											assign node2215 = (inp[12]) ? node2219 : node2216;
												assign node2216 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2219 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2222 = (inp[9]) ? node2226 : node2223;
												assign node2223 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2226 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node2229 = (inp[4]) ? node2237 : node2230;
											assign node2230 = (inp[14]) ? node2234 : node2231;
												assign node2231 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2234 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2237 = (inp[7]) ? node2241 : node2238;
												assign node2238 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2241 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2244 = (inp[7]) ? node2276 : node2245;
									assign node2245 = (inp[15]) ? node2261 : node2246;
										assign node2246 = (inp[4]) ? node2254 : node2247;
											assign node2247 = (inp[10]) ? node2251 : node2248;
												assign node2248 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2251 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2254 = (inp[12]) ? node2258 : node2255;
												assign node2255 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2258 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2261 = (inp[12]) ? node2269 : node2262;
											assign node2262 = (inp[10]) ? node2266 : node2263;
												assign node2263 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2266 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2269 = (inp[14]) ? node2273 : node2270;
												assign node2270 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2273 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2276 = (inp[0]) ? node2292 : node2277;
										assign node2277 = (inp[5]) ? node2285 : node2278;
											assign node2278 = (inp[4]) ? node2282 : node2279;
												assign node2279 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2282 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2285 = (inp[15]) ? node2289 : node2286;
												assign node2286 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2289 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2292 = (inp[12]) ? node2300 : node2293;
											assign node2293 = (inp[5]) ? node2297 : node2294;
												assign node2294 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2297 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2300 = (inp[14]) ? node2304 : node2301;
												assign node2301 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2304 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node2307 = (inp[0]) ? node2435 : node2308;
							assign node2308 = (inp[9]) ? node2372 : node2309;
								assign node2309 = (inp[7]) ? node2341 : node2310;
									assign node2310 = (inp[14]) ? node2326 : node2311;
										assign node2311 = (inp[12]) ? node2319 : node2312;
											assign node2312 = (inp[15]) ? node2316 : node2313;
												assign node2313 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2316 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2319 = (inp[8]) ? node2323 : node2320;
												assign node2320 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2323 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2326 = (inp[6]) ? node2334 : node2327;
											assign node2327 = (inp[12]) ? node2331 : node2328;
												assign node2328 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2331 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2334 = (inp[12]) ? node2338 : node2335;
												assign node2335 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2338 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2341 = (inp[4]) ? node2357 : node2342;
										assign node2342 = (inp[12]) ? node2350 : node2343;
											assign node2343 = (inp[6]) ? node2347 : node2344;
												assign node2344 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2347 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2350 = (inp[8]) ? node2354 : node2351;
												assign node2351 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2354 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2357 = (inp[5]) ? node2365 : node2358;
											assign node2358 = (inp[8]) ? node2362 : node2359;
												assign node2359 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2362 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2365 = (inp[12]) ? node2369 : node2366;
												assign node2366 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2369 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node2372 = (inp[4]) ? node2404 : node2373;
									assign node2373 = (inp[10]) ? node2389 : node2374;
										assign node2374 = (inp[5]) ? node2382 : node2375;
											assign node2375 = (inp[15]) ? node2379 : node2376;
												assign node2376 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2379 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2382 = (inp[7]) ? node2386 : node2383;
												assign node2383 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2386 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2389 = (inp[8]) ? node2397 : node2390;
											assign node2390 = (inp[7]) ? node2394 : node2391;
												assign node2391 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2394 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2397 = (inp[12]) ? node2401 : node2398;
												assign node2398 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2401 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2404 = (inp[8]) ? node2420 : node2405;
										assign node2405 = (inp[7]) ? node2413 : node2406;
											assign node2406 = (inp[14]) ? node2410 : node2407;
												assign node2407 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2410 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2413 = (inp[6]) ? node2417 : node2414;
												assign node2414 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2417 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2420 = (inp[5]) ? node2428 : node2421;
											assign node2421 = (inp[12]) ? node2425 : node2422;
												assign node2422 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2425 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2428 = (inp[14]) ? node2432 : node2429;
												assign node2429 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2432 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node2435 = (inp[10]) ? node2499 : node2436;
								assign node2436 = (inp[7]) ? node2468 : node2437;
									assign node2437 = (inp[6]) ? node2453 : node2438;
										assign node2438 = (inp[8]) ? node2446 : node2439;
											assign node2439 = (inp[5]) ? node2443 : node2440;
												assign node2440 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2443 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2446 = (inp[9]) ? node2450 : node2447;
												assign node2447 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2450 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2453 = (inp[12]) ? node2461 : node2454;
											assign node2454 = (inp[9]) ? node2458 : node2455;
												assign node2455 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2458 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2461 = (inp[15]) ? node2465 : node2462;
												assign node2462 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2465 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2468 = (inp[9]) ? node2484 : node2469;
										assign node2469 = (inp[4]) ? node2477 : node2470;
											assign node2470 = (inp[5]) ? node2474 : node2471;
												assign node2471 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2474 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2477 = (inp[12]) ? node2481 : node2478;
												assign node2478 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2481 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2484 = (inp[14]) ? node2492 : node2485;
											assign node2485 = (inp[8]) ? node2489 : node2486;
												assign node2486 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2489 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2492 = (inp[6]) ? node2496 : node2493;
												assign node2493 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2496 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
								assign node2499 = (inp[9]) ? node2531 : node2500;
									assign node2500 = (inp[5]) ? node2516 : node2501;
										assign node2501 = (inp[15]) ? node2509 : node2502;
											assign node2502 = (inp[7]) ? node2506 : node2503;
												assign node2503 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2506 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2509 = (inp[8]) ? node2513 : node2510;
												assign node2510 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2513 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2516 = (inp[12]) ? node2524 : node2517;
											assign node2517 = (inp[7]) ? node2521 : node2518;
												assign node2518 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2521 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2524 = (inp[8]) ? node2528 : node2525;
												assign node2525 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2528 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2531 = (inp[14]) ? node2547 : node2532;
										assign node2532 = (inp[5]) ? node2540 : node2533;
											assign node2533 = (inp[6]) ? node2537 : node2534;
												assign node2534 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2537 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2540 = (inp[12]) ? node2544 : node2541;
												assign node2541 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2544 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node2547 = (inp[6]) ? node2555 : node2548;
											assign node2548 = (inp[15]) ? node2552 : node2549;
												assign node2549 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2552 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2555 = (inp[8]) ? node2559 : node2556;
												assign node2556 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2559 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node2562 = (inp[14]) ? node2818 : node2563;
						assign node2563 = (inp[9]) ? node2691 : node2564;
							assign node2564 = (inp[0]) ? node2628 : node2565;
								assign node2565 = (inp[4]) ? node2597 : node2566;
									assign node2566 = (inp[15]) ? node2582 : node2567;
										assign node2567 = (inp[8]) ? node2575 : node2568;
											assign node2568 = (inp[10]) ? node2572 : node2569;
												assign node2569 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2572 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2575 = (inp[2]) ? node2579 : node2576;
												assign node2576 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2579 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2582 = (inp[2]) ? node2590 : node2583;
											assign node2583 = (inp[10]) ? node2587 : node2584;
												assign node2584 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2587 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2590 = (inp[10]) ? node2594 : node2591;
												assign node2591 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2594 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2597 = (inp[7]) ? node2613 : node2598;
										assign node2598 = (inp[6]) ? node2606 : node2599;
											assign node2599 = (inp[5]) ? node2603 : node2600;
												assign node2600 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2603 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2606 = (inp[12]) ? node2610 : node2607;
												assign node2607 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2610 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2613 = (inp[12]) ? node2621 : node2614;
											assign node2614 = (inp[8]) ? node2618 : node2615;
												assign node2615 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2618 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2621 = (inp[15]) ? node2625 : node2622;
												assign node2622 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2625 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2628 = (inp[6]) ? node2660 : node2629;
									assign node2629 = (inp[10]) ? node2645 : node2630;
										assign node2630 = (inp[15]) ? node2638 : node2631;
											assign node2631 = (inp[4]) ? node2635 : node2632;
												assign node2632 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2635 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2638 = (inp[5]) ? node2642 : node2639;
												assign node2639 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2642 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2645 = (inp[12]) ? node2653 : node2646;
											assign node2646 = (inp[8]) ? node2650 : node2647;
												assign node2647 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2650 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2653 = (inp[15]) ? node2657 : node2654;
												assign node2654 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2657 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2660 = (inp[10]) ? node2676 : node2661;
										assign node2661 = (inp[8]) ? node2669 : node2662;
											assign node2662 = (inp[2]) ? node2666 : node2663;
												assign node2663 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2666 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2669 = (inp[5]) ? node2673 : node2670;
												assign node2670 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2673 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2676 = (inp[7]) ? node2684 : node2677;
											assign node2677 = (inp[15]) ? node2681 : node2678;
												assign node2678 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2681 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2684 = (inp[8]) ? node2688 : node2685;
												assign node2685 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2688 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node2691 = (inp[0]) ? node2755 : node2692;
								assign node2692 = (inp[12]) ? node2724 : node2693;
									assign node2693 = (inp[2]) ? node2709 : node2694;
										assign node2694 = (inp[7]) ? node2702 : node2695;
											assign node2695 = (inp[10]) ? node2699 : node2696;
												assign node2696 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2699 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2702 = (inp[8]) ? node2706 : node2703;
												assign node2703 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2706 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2709 = (inp[8]) ? node2717 : node2710;
											assign node2710 = (inp[10]) ? node2714 : node2711;
												assign node2711 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2714 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2717 = (inp[4]) ? node2721 : node2718;
												assign node2718 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2721 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2724 = (inp[6]) ? node2740 : node2725;
										assign node2725 = (inp[4]) ? node2733 : node2726;
											assign node2726 = (inp[5]) ? node2730 : node2727;
												assign node2727 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2730 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2733 = (inp[15]) ? node2737 : node2734;
												assign node2734 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2737 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2740 = (inp[10]) ? node2748 : node2741;
											assign node2741 = (inp[15]) ? node2745 : node2742;
												assign node2742 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2745 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2748 = (inp[5]) ? node2752 : node2749;
												assign node2749 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2752 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2755 = (inp[15]) ? node2787 : node2756;
									assign node2756 = (inp[4]) ? node2772 : node2757;
										assign node2757 = (inp[10]) ? node2765 : node2758;
											assign node2758 = (inp[8]) ? node2762 : node2759;
												assign node2759 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2762 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2765 = (inp[5]) ? node2769 : node2766;
												assign node2766 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2769 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2772 = (inp[7]) ? node2780 : node2773;
											assign node2773 = (inp[6]) ? node2777 : node2774;
												assign node2774 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2777 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node2780 = (inp[12]) ? node2784 : node2781;
												assign node2781 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2784 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2787 = (inp[10]) ? node2803 : node2788;
										assign node2788 = (inp[8]) ? node2796 : node2789;
											assign node2789 = (inp[2]) ? node2793 : node2790;
												assign node2790 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2793 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2796 = (inp[5]) ? node2800 : node2797;
												assign node2797 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2800 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2803 = (inp[12]) ? node2811 : node2804;
											assign node2804 = (inp[4]) ? node2808 : node2805;
												assign node2805 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2808 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2811 = (inp[7]) ? node2815 : node2812;
												assign node2812 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2815 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node2818 = (inp[10]) ? node2946 : node2819;
							assign node2819 = (inp[12]) ? node2883 : node2820;
								assign node2820 = (inp[4]) ? node2852 : node2821;
									assign node2821 = (inp[6]) ? node2837 : node2822;
										assign node2822 = (inp[0]) ? node2830 : node2823;
											assign node2823 = (inp[2]) ? node2827 : node2824;
												assign node2824 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2827 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2830 = (inp[9]) ? node2834 : node2831;
												assign node2831 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2834 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2837 = (inp[0]) ? node2845 : node2838;
											assign node2838 = (inp[9]) ? node2842 : node2839;
												assign node2839 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2842 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2845 = (inp[7]) ? node2849 : node2846;
												assign node2846 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2849 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2852 = (inp[8]) ? node2868 : node2853;
										assign node2853 = (inp[15]) ? node2861 : node2854;
											assign node2854 = (inp[0]) ? node2858 : node2855;
												assign node2855 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2858 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2861 = (inp[9]) ? node2865 : node2862;
												assign node2862 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2865 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2868 = (inp[5]) ? node2876 : node2869;
											assign node2869 = (inp[0]) ? node2873 : node2870;
												assign node2870 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2873 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2876 = (inp[7]) ? node2880 : node2877;
												assign node2877 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2880 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2883 = (inp[7]) ? node2915 : node2884;
									assign node2884 = (inp[5]) ? node2900 : node2885;
										assign node2885 = (inp[8]) ? node2893 : node2886;
											assign node2886 = (inp[6]) ? node2890 : node2887;
												assign node2887 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2890 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2893 = (inp[0]) ? node2897 : node2894;
												assign node2894 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2897 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2900 = (inp[4]) ? node2908 : node2901;
											assign node2901 = (inp[9]) ? node2905 : node2902;
												assign node2902 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2905 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2908 = (inp[2]) ? node2912 : node2909;
												assign node2909 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2912 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2915 = (inp[15]) ? node2931 : node2916;
										assign node2916 = (inp[5]) ? node2924 : node2917;
											assign node2917 = (inp[8]) ? node2921 : node2918;
												assign node2918 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2921 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2924 = (inp[0]) ? node2928 : node2925;
												assign node2925 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2928 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2931 = (inp[9]) ? node2939 : node2932;
											assign node2932 = (inp[0]) ? node2936 : node2933;
												assign node2933 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2936 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2939 = (inp[5]) ? node2943 : node2940;
												assign node2940 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2943 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node2946 = (inp[2]) ? node3010 : node2947;
								assign node2947 = (inp[8]) ? node2979 : node2948;
									assign node2948 = (inp[15]) ? node2964 : node2949;
										assign node2949 = (inp[9]) ? node2957 : node2950;
											assign node2950 = (inp[6]) ? node2954 : node2951;
												assign node2951 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2954 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2957 = (inp[7]) ? node2961 : node2958;
												assign node2958 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2961 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2964 = (inp[7]) ? node2972 : node2965;
											assign node2965 = (inp[12]) ? node2969 : node2966;
												assign node2966 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2969 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2972 = (inp[0]) ? node2976 : node2973;
												assign node2973 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2976 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2979 = (inp[4]) ? node2995 : node2980;
										assign node2980 = (inp[6]) ? node2988 : node2981;
											assign node2981 = (inp[15]) ? node2985 : node2982;
												assign node2982 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2985 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2988 = (inp[15]) ? node2992 : node2989;
												assign node2989 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2992 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2995 = (inp[6]) ? node3003 : node2996;
											assign node2996 = (inp[12]) ? node3000 : node2997;
												assign node2997 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3000 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3003 = (inp[5]) ? node3007 : node3004;
												assign node3004 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3007 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3010 = (inp[4]) ? node3042 : node3011;
									assign node3011 = (inp[7]) ? node3027 : node3012;
										assign node3012 = (inp[15]) ? node3020 : node3013;
											assign node3013 = (inp[6]) ? node3017 : node3014;
												assign node3014 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3017 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3020 = (inp[5]) ? node3024 : node3021;
												assign node3021 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3024 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3027 = (inp[5]) ? node3035 : node3028;
											assign node3028 = (inp[0]) ? node3032 : node3029;
												assign node3029 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3032 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3035 = (inp[9]) ? node3039 : node3036;
												assign node3036 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3039 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3042 = (inp[12]) ? node3058 : node3043;
										assign node3043 = (inp[6]) ? node3051 : node3044;
											assign node3044 = (inp[7]) ? node3048 : node3045;
												assign node3045 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3048 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3051 = (inp[15]) ? node3055 : node3052;
												assign node3052 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3055 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3058 = (inp[9]) ? node3066 : node3059;
											assign node3059 = (inp[7]) ? node3063 : node3060;
												assign node3060 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3063 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3066 = (inp[15]) ? node3070 : node3067;
												assign node3067 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3070 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
				assign node3073 = (inp[12]) ? node3585 : node3074;
					assign node3074 = (inp[5]) ? node3330 : node3075;
						assign node3075 = (inp[10]) ? node3203 : node3076;
							assign node3076 = (inp[9]) ? node3140 : node3077;
								assign node3077 = (inp[7]) ? node3109 : node3078;
									assign node3078 = (inp[15]) ? node3094 : node3079;
										assign node3079 = (inp[0]) ? node3087 : node3080;
											assign node3080 = (inp[6]) ? node3084 : node3081;
												assign node3081 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3084 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3087 = (inp[8]) ? node3091 : node3088;
												assign node3088 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3091 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3094 = (inp[13]) ? node3102 : node3095;
											assign node3095 = (inp[8]) ? node3099 : node3096;
												assign node3096 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3099 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3102 = (inp[2]) ? node3106 : node3103;
												assign node3103 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3106 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3109 = (inp[8]) ? node3125 : node3110;
										assign node3110 = (inp[2]) ? node3118 : node3111;
											assign node3111 = (inp[6]) ? node3115 : node3112;
												assign node3112 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3115 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3118 = (inp[4]) ? node3122 : node3119;
												assign node3119 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3122 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3125 = (inp[6]) ? node3133 : node3126;
											assign node3126 = (inp[0]) ? node3130 : node3127;
												assign node3127 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3130 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3133 = (inp[2]) ? node3137 : node3134;
												assign node3134 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3137 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node3140 = (inp[14]) ? node3172 : node3141;
									assign node3141 = (inp[6]) ? node3157 : node3142;
										assign node3142 = (inp[0]) ? node3150 : node3143;
											assign node3143 = (inp[13]) ? node3147 : node3144;
												assign node3144 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3147 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3150 = (inp[4]) ? node3154 : node3151;
												assign node3151 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3154 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3157 = (inp[8]) ? node3165 : node3158;
											assign node3158 = (inp[7]) ? node3162 : node3159;
												assign node3159 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3162 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3165 = (inp[15]) ? node3169 : node3166;
												assign node3166 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3169 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3172 = (inp[2]) ? node3188 : node3173;
										assign node3173 = (inp[4]) ? node3181 : node3174;
											assign node3174 = (inp[6]) ? node3178 : node3175;
												assign node3175 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3178 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3181 = (inp[15]) ? node3185 : node3182;
												assign node3182 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3185 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3188 = (inp[0]) ? node3196 : node3189;
											assign node3189 = (inp[8]) ? node3193 : node3190;
												assign node3190 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3193 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3196 = (inp[7]) ? node3200 : node3197;
												assign node3197 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3200 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node3203 = (inp[4]) ? node3267 : node3204;
								assign node3204 = (inp[6]) ? node3236 : node3205;
									assign node3205 = (inp[8]) ? node3221 : node3206;
										assign node3206 = (inp[15]) ? node3214 : node3207;
											assign node3207 = (inp[13]) ? node3211 : node3208;
												assign node3208 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3211 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3214 = (inp[0]) ? node3218 : node3215;
												assign node3215 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3218 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3221 = (inp[14]) ? node3229 : node3222;
											assign node3222 = (inp[0]) ? node3226 : node3223;
												assign node3223 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3226 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3229 = (inp[9]) ? node3233 : node3230;
												assign node3230 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3233 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3236 = (inp[2]) ? node3252 : node3237;
										assign node3237 = (inp[13]) ? node3245 : node3238;
											assign node3238 = (inp[15]) ? node3242 : node3239;
												assign node3239 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3242 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3245 = (inp[7]) ? node3249 : node3246;
												assign node3246 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3249 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3252 = (inp[8]) ? node3260 : node3253;
											assign node3253 = (inp[7]) ? node3257 : node3254;
												assign node3254 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3257 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3260 = (inp[9]) ? node3264 : node3261;
												assign node3261 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3264 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3267 = (inp[13]) ? node3299 : node3268;
									assign node3268 = (inp[7]) ? node3284 : node3269;
										assign node3269 = (inp[14]) ? node3277 : node3270;
											assign node3270 = (inp[2]) ? node3274 : node3271;
												assign node3271 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3274 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3277 = (inp[9]) ? node3281 : node3278;
												assign node3278 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3281 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3284 = (inp[0]) ? node3292 : node3285;
											assign node3285 = (inp[8]) ? node3289 : node3286;
												assign node3286 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3289 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3292 = (inp[8]) ? node3296 : node3293;
												assign node3293 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3296 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3299 = (inp[14]) ? node3315 : node3300;
										assign node3300 = (inp[15]) ? node3308 : node3301;
											assign node3301 = (inp[7]) ? node3305 : node3302;
												assign node3302 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3305 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3308 = (inp[2]) ? node3312 : node3309;
												assign node3309 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3312 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3315 = (inp[2]) ? node3323 : node3316;
											assign node3316 = (inp[0]) ? node3320 : node3317;
												assign node3317 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3320 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3323 = (inp[8]) ? node3327 : node3324;
												assign node3324 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3327 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node3330 = (inp[10]) ? node3458 : node3331;
							assign node3331 = (inp[8]) ? node3395 : node3332;
								assign node3332 = (inp[13]) ? node3364 : node3333;
									assign node3333 = (inp[9]) ? node3349 : node3334;
										assign node3334 = (inp[6]) ? node3342 : node3335;
											assign node3335 = (inp[2]) ? node3339 : node3336;
												assign node3336 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3339 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3342 = (inp[0]) ? node3346 : node3343;
												assign node3343 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3346 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3349 = (inp[15]) ? node3357 : node3350;
											assign node3350 = (inp[4]) ? node3354 : node3351;
												assign node3351 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3354 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3357 = (inp[6]) ? node3361 : node3358;
												assign node3358 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3361 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3364 = (inp[7]) ? node3380 : node3365;
										assign node3365 = (inp[9]) ? node3373 : node3366;
											assign node3366 = (inp[4]) ? node3370 : node3367;
												assign node3367 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3370 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3373 = (inp[14]) ? node3377 : node3374;
												assign node3374 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3377 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3380 = (inp[15]) ? node3388 : node3381;
											assign node3381 = (inp[4]) ? node3385 : node3382;
												assign node3382 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3385 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3388 = (inp[2]) ? node3392 : node3389;
												assign node3389 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3392 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3395 = (inp[9]) ? node3427 : node3396;
									assign node3396 = (inp[14]) ? node3412 : node3397;
										assign node3397 = (inp[15]) ? node3405 : node3398;
											assign node3398 = (inp[7]) ? node3402 : node3399;
												assign node3399 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3402 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3405 = (inp[2]) ? node3409 : node3406;
												assign node3406 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3409 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3412 = (inp[0]) ? node3420 : node3413;
											assign node3413 = (inp[6]) ? node3417 : node3414;
												assign node3414 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3417 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3420 = (inp[13]) ? node3424 : node3421;
												assign node3421 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3424 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3427 = (inp[2]) ? node3443 : node3428;
										assign node3428 = (inp[14]) ? node3436 : node3429;
											assign node3429 = (inp[13]) ? node3433 : node3430;
												assign node3430 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3433 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3436 = (inp[7]) ? node3440 : node3437;
												assign node3437 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3440 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3443 = (inp[4]) ? node3451 : node3444;
											assign node3444 = (inp[0]) ? node3448 : node3445;
												assign node3445 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3448 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3451 = (inp[14]) ? node3455 : node3452;
												assign node3452 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3455 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node3458 = (inp[4]) ? node3522 : node3459;
								assign node3459 = (inp[7]) ? node3491 : node3460;
									assign node3460 = (inp[2]) ? node3476 : node3461;
										assign node3461 = (inp[9]) ? node3469 : node3462;
											assign node3462 = (inp[14]) ? node3466 : node3463;
												assign node3463 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3466 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3469 = (inp[15]) ? node3473 : node3470;
												assign node3470 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3473 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3476 = (inp[15]) ? node3484 : node3477;
											assign node3477 = (inp[0]) ? node3481 : node3478;
												assign node3478 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3481 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3484 = (inp[14]) ? node3488 : node3485;
												assign node3485 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3488 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3491 = (inp[14]) ? node3507 : node3492;
										assign node3492 = (inp[6]) ? node3500 : node3493;
											assign node3493 = (inp[2]) ? node3497 : node3494;
												assign node3494 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3497 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3500 = (inp[13]) ? node3504 : node3501;
												assign node3501 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3504 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3507 = (inp[8]) ? node3515 : node3508;
											assign node3508 = (inp[15]) ? node3512 : node3509;
												assign node3509 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3512 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3515 = (inp[0]) ? node3519 : node3516;
												assign node3516 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3519 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3522 = (inp[2]) ? node3554 : node3523;
									assign node3523 = (inp[13]) ? node3539 : node3524;
										assign node3524 = (inp[9]) ? node3532 : node3525;
											assign node3525 = (inp[15]) ? node3529 : node3526;
												assign node3526 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3529 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3532 = (inp[14]) ? node3536 : node3533;
												assign node3533 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3536 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3539 = (inp[14]) ? node3547 : node3540;
											assign node3540 = (inp[15]) ? node3544 : node3541;
												assign node3541 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3544 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3547 = (inp[9]) ? node3551 : node3548;
												assign node3548 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3551 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3554 = (inp[14]) ? node3570 : node3555;
										assign node3555 = (inp[6]) ? node3563 : node3556;
											assign node3556 = (inp[0]) ? node3560 : node3557;
												assign node3557 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3560 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3563 = (inp[9]) ? node3567 : node3564;
												assign node3564 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3567 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3570 = (inp[7]) ? node3578 : node3571;
											assign node3571 = (inp[15]) ? node3575 : node3572;
												assign node3572 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3575 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3578 = (inp[0]) ? node3582 : node3579;
												assign node3579 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3582 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node3585 = (inp[14]) ? node3841 : node3586;
						assign node3586 = (inp[7]) ? node3714 : node3587;
							assign node3587 = (inp[9]) ? node3651 : node3588;
								assign node3588 = (inp[6]) ? node3620 : node3589;
									assign node3589 = (inp[10]) ? node3605 : node3590;
										assign node3590 = (inp[2]) ? node3598 : node3591;
											assign node3591 = (inp[0]) ? node3595 : node3592;
												assign node3592 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3595 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3598 = (inp[13]) ? node3602 : node3599;
												assign node3599 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3602 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3605 = (inp[4]) ? node3613 : node3606;
											assign node3606 = (inp[0]) ? node3610 : node3607;
												assign node3607 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3610 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3613 = (inp[13]) ? node3617 : node3614;
												assign node3614 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3617 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3620 = (inp[5]) ? node3636 : node3621;
										assign node3621 = (inp[15]) ? node3629 : node3622;
											assign node3622 = (inp[4]) ? node3626 : node3623;
												assign node3623 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3626 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3629 = (inp[4]) ? node3633 : node3630;
												assign node3630 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3633 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3636 = (inp[0]) ? node3644 : node3637;
											assign node3637 = (inp[4]) ? node3641 : node3638;
												assign node3638 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3641 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3644 = (inp[8]) ? node3648 : node3645;
												assign node3645 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3648 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3651 = (inp[0]) ? node3683 : node3652;
									assign node3652 = (inp[13]) ? node3668 : node3653;
										assign node3653 = (inp[2]) ? node3661 : node3654;
											assign node3654 = (inp[4]) ? node3658 : node3655;
												assign node3655 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3658 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3661 = (inp[8]) ? node3665 : node3662;
												assign node3662 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3665 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3668 = (inp[15]) ? node3676 : node3669;
											assign node3669 = (inp[8]) ? node3673 : node3670;
												assign node3670 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3673 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node3676 = (inp[5]) ? node3680 : node3677;
												assign node3677 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3680 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3683 = (inp[15]) ? node3699 : node3684;
										assign node3684 = (inp[13]) ? node3692 : node3685;
											assign node3685 = (inp[2]) ? node3689 : node3686;
												assign node3686 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3689 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3692 = (inp[8]) ? node3696 : node3693;
												assign node3693 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3696 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3699 = (inp[10]) ? node3707 : node3700;
											assign node3700 = (inp[13]) ? node3704 : node3701;
												assign node3701 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3704 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3707 = (inp[5]) ? node3711 : node3708;
												assign node3708 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3711 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node3714 = (inp[0]) ? node3778 : node3715;
								assign node3715 = (inp[6]) ? node3747 : node3716;
									assign node3716 = (inp[10]) ? node3732 : node3717;
										assign node3717 = (inp[2]) ? node3725 : node3718;
											assign node3718 = (inp[4]) ? node3722 : node3719;
												assign node3719 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3722 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3725 = (inp[8]) ? node3729 : node3726;
												assign node3726 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3729 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node3732 = (inp[8]) ? node3740 : node3733;
											assign node3733 = (inp[2]) ? node3737 : node3734;
												assign node3734 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3737 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3740 = (inp[5]) ? node3744 : node3741;
												assign node3741 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3744 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3747 = (inp[4]) ? node3763 : node3748;
										assign node3748 = (inp[13]) ? node3756 : node3749;
											assign node3749 = (inp[15]) ? node3753 : node3750;
												assign node3750 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3753 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3756 = (inp[8]) ? node3760 : node3757;
												assign node3757 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node3760 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3763 = (inp[5]) ? node3771 : node3764;
											assign node3764 = (inp[8]) ? node3768 : node3765;
												assign node3765 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3768 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3771 = (inp[8]) ? node3775 : node3772;
												assign node3772 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3775 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3778 = (inp[10]) ? node3810 : node3779;
									assign node3779 = (inp[2]) ? node3795 : node3780;
										assign node3780 = (inp[8]) ? node3788 : node3781;
											assign node3781 = (inp[5]) ? node3785 : node3782;
												assign node3782 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3785 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3788 = (inp[15]) ? node3792 : node3789;
												assign node3789 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3792 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3795 = (inp[9]) ? node3803 : node3796;
											assign node3796 = (inp[5]) ? node3800 : node3797;
												assign node3797 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3800 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3803 = (inp[13]) ? node3807 : node3804;
												assign node3804 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3807 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3810 = (inp[4]) ? node3826 : node3811;
										assign node3811 = (inp[15]) ? node3819 : node3812;
											assign node3812 = (inp[6]) ? node3816 : node3813;
												assign node3813 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3816 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3819 = (inp[13]) ? node3823 : node3820;
												assign node3820 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3823 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3826 = (inp[2]) ? node3834 : node3827;
											assign node3827 = (inp[6]) ? node3831 : node3828;
												assign node3828 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3831 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3834 = (inp[8]) ? node3838 : node3835;
												assign node3835 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3838 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node3841 = (inp[2]) ? node3969 : node3842;
							assign node3842 = (inp[6]) ? node3906 : node3843;
								assign node3843 = (inp[15]) ? node3875 : node3844;
									assign node3844 = (inp[5]) ? node3860 : node3845;
										assign node3845 = (inp[8]) ? node3853 : node3846;
											assign node3846 = (inp[7]) ? node3850 : node3847;
												assign node3847 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3850 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3853 = (inp[0]) ? node3857 : node3854;
												assign node3854 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3857 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3860 = (inp[7]) ? node3868 : node3861;
											assign node3861 = (inp[4]) ? node3865 : node3862;
												assign node3862 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3865 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3868 = (inp[13]) ? node3872 : node3869;
												assign node3869 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3872 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3875 = (inp[9]) ? node3891 : node3876;
										assign node3876 = (inp[10]) ? node3884 : node3877;
											assign node3877 = (inp[8]) ? node3881 : node3878;
												assign node3878 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3881 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3884 = (inp[5]) ? node3888 : node3885;
												assign node3885 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3888 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3891 = (inp[0]) ? node3899 : node3892;
											assign node3892 = (inp[10]) ? node3896 : node3893;
												assign node3893 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3896 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3899 = (inp[13]) ? node3903 : node3900;
												assign node3900 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3903 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3906 = (inp[10]) ? node3938 : node3907;
									assign node3907 = (inp[8]) ? node3923 : node3908;
										assign node3908 = (inp[15]) ? node3916 : node3909;
											assign node3909 = (inp[13]) ? node3913 : node3910;
												assign node3910 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3913 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3916 = (inp[9]) ? node3920 : node3917;
												assign node3917 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3920 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3923 = (inp[7]) ? node3931 : node3924;
											assign node3924 = (inp[4]) ? node3928 : node3925;
												assign node3925 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3928 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3931 = (inp[9]) ? node3935 : node3932;
												assign node3932 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3935 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3938 = (inp[4]) ? node3954 : node3939;
										assign node3939 = (inp[5]) ? node3947 : node3940;
											assign node3940 = (inp[13]) ? node3944 : node3941;
												assign node3941 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3944 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3947 = (inp[7]) ? node3951 : node3948;
												assign node3948 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3951 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3954 = (inp[15]) ? node3962 : node3955;
											assign node3955 = (inp[9]) ? node3959 : node3956;
												assign node3956 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3959 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3962 = (inp[0]) ? node3966 : node3963;
												assign node3963 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3966 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node3969 = (inp[13]) ? node4033 : node3970;
								assign node3970 = (inp[4]) ? node4002 : node3971;
									assign node3971 = (inp[8]) ? node3987 : node3972;
										assign node3972 = (inp[7]) ? node3980 : node3973;
											assign node3973 = (inp[15]) ? node3977 : node3974;
												assign node3974 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3977 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3980 = (inp[10]) ? node3984 : node3981;
												assign node3981 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3984 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3987 = (inp[6]) ? node3995 : node3988;
											assign node3988 = (inp[7]) ? node3992 : node3989;
												assign node3989 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3992 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3995 = (inp[9]) ? node3999 : node3996;
												assign node3996 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3999 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4002 = (inp[9]) ? node4018 : node4003;
										assign node4003 = (inp[10]) ? node4011 : node4004;
											assign node4004 = (inp[6]) ? node4008 : node4005;
												assign node4005 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4008 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4011 = (inp[8]) ? node4015 : node4012;
												assign node4012 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4015 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4018 = (inp[8]) ? node4026 : node4019;
											assign node4019 = (inp[10]) ? node4023 : node4020;
												assign node4020 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4023 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4026 = (inp[6]) ? node4030 : node4027;
												assign node4027 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4030 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node4033 = (inp[5]) ? node4065 : node4034;
									assign node4034 = (inp[9]) ? node4050 : node4035;
										assign node4035 = (inp[4]) ? node4043 : node4036;
											assign node4036 = (inp[10]) ? node4040 : node4037;
												assign node4037 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4040 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4043 = (inp[15]) ? node4047 : node4044;
												assign node4044 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4047 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4050 = (inp[6]) ? node4058 : node4051;
											assign node4051 = (inp[8]) ? node4055 : node4052;
												assign node4052 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4055 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4058 = (inp[10]) ? node4062 : node4059;
												assign node4059 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4062 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node4065 = (inp[0]) ? node4081 : node4066;
										assign node4066 = (inp[15]) ? node4074 : node4067;
											assign node4067 = (inp[6]) ? node4071 : node4068;
												assign node4068 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4071 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4074 = (inp[9]) ? node4078 : node4075;
												assign node4075 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4078 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node4081 = (inp[4]) ? node4089 : node4082;
											assign node4082 = (inp[6]) ? node4086 : node4083;
												assign node4083 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4086 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4089 = (inp[8]) ? node4093 : node4090;
												assign node4090 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node4093 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
		assign node4096 = (inp[6]) ? node6144 : node4097;
			assign node4097 = (inp[0]) ? node5121 : node4098;
				assign node4098 = (inp[11]) ? node4610 : node4099;
					assign node4099 = (inp[4]) ? node4355 : node4100;
						assign node4100 = (inp[9]) ? node4228 : node4101;
							assign node4101 = (inp[14]) ? node4165 : node4102;
								assign node4102 = (inp[15]) ? node4134 : node4103;
									assign node4103 = (inp[2]) ? node4119 : node4104;
										assign node4104 = (inp[5]) ? node4112 : node4105;
											assign node4105 = (inp[8]) ? node4109 : node4106;
												assign node4106 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node4109 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node4112 = (inp[13]) ? node4116 : node4113;
												assign node4113 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4116 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node4119 = (inp[5]) ? node4127 : node4120;
											assign node4120 = (inp[12]) ? node4124 : node4121;
												assign node4121 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4124 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4127 = (inp[13]) ? node4131 : node4128;
												assign node4128 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4131 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node4134 = (inp[10]) ? node4150 : node4135;
										assign node4135 = (inp[3]) ? node4143 : node4136;
											assign node4136 = (inp[2]) ? node4140 : node4137;
												assign node4137 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4140 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4143 = (inp[5]) ? node4147 : node4144;
												assign node4144 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4147 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4150 = (inp[13]) ? node4158 : node4151;
											assign node4151 = (inp[5]) ? node4155 : node4152;
												assign node4152 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4155 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4158 = (inp[3]) ? node4162 : node4159;
												assign node4159 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4162 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node4165 = (inp[8]) ? node4197 : node4166;
									assign node4166 = (inp[5]) ? node4182 : node4167;
										assign node4167 = (inp[3]) ? node4175 : node4168;
											assign node4168 = (inp[15]) ? node4172 : node4169;
												assign node4169 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4172 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4175 = (inp[15]) ? node4179 : node4176;
												assign node4176 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4179 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4182 = (inp[3]) ? node4190 : node4183;
											assign node4183 = (inp[2]) ? node4187 : node4184;
												assign node4184 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4187 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4190 = (inp[7]) ? node4194 : node4191;
												assign node4191 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4194 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4197 = (inp[10]) ? node4213 : node4198;
										assign node4198 = (inp[7]) ? node4206 : node4199;
											assign node4199 = (inp[15]) ? node4203 : node4200;
												assign node4200 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4203 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4206 = (inp[2]) ? node4210 : node4207;
												assign node4207 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4210 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4213 = (inp[15]) ? node4221 : node4214;
											assign node4214 = (inp[7]) ? node4218 : node4215;
												assign node4215 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4218 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4221 = (inp[12]) ? node4225 : node4222;
												assign node4222 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4225 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
							assign node4228 = (inp[7]) ? node4292 : node4229;
								assign node4229 = (inp[5]) ? node4261 : node4230;
									assign node4230 = (inp[12]) ? node4246 : node4231;
										assign node4231 = (inp[8]) ? node4239 : node4232;
											assign node4232 = (inp[10]) ? node4236 : node4233;
												assign node4233 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4236 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4239 = (inp[14]) ? node4243 : node4240;
												assign node4240 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4243 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4246 = (inp[13]) ? node4254 : node4247;
											assign node4247 = (inp[14]) ? node4251 : node4248;
												assign node4248 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4251 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4254 = (inp[10]) ? node4258 : node4255;
												assign node4255 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4258 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4261 = (inp[15]) ? node4277 : node4262;
										assign node4262 = (inp[2]) ? node4270 : node4263;
											assign node4263 = (inp[3]) ? node4267 : node4264;
												assign node4264 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4267 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4270 = (inp[8]) ? node4274 : node4271;
												assign node4271 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4274 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4277 = (inp[2]) ? node4285 : node4278;
											assign node4278 = (inp[12]) ? node4282 : node4279;
												assign node4279 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4282 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4285 = (inp[10]) ? node4289 : node4286;
												assign node4286 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4289 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node4292 = (inp[13]) ? node4324 : node4293;
									assign node4293 = (inp[2]) ? node4309 : node4294;
										assign node4294 = (inp[14]) ? node4302 : node4295;
											assign node4295 = (inp[10]) ? node4299 : node4296;
												assign node4296 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4299 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4302 = (inp[3]) ? node4306 : node4303;
												assign node4303 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4306 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4309 = (inp[8]) ? node4317 : node4310;
											assign node4310 = (inp[3]) ? node4314 : node4311;
												assign node4311 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4314 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4317 = (inp[10]) ? node4321 : node4318;
												assign node4318 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4321 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4324 = (inp[10]) ? node4340 : node4325;
										assign node4325 = (inp[15]) ? node4333 : node4326;
											assign node4326 = (inp[8]) ? node4330 : node4327;
												assign node4327 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4330 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4333 = (inp[2]) ? node4337 : node4334;
												assign node4334 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4337 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4340 = (inp[5]) ? node4348 : node4341;
											assign node4341 = (inp[14]) ? node4345 : node4342;
												assign node4342 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4345 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4348 = (inp[2]) ? node4352 : node4349;
												assign node4349 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4352 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
						assign node4355 = (inp[8]) ? node4483 : node4356;
							assign node4356 = (inp[2]) ? node4420 : node4357;
								assign node4357 = (inp[12]) ? node4389 : node4358;
									assign node4358 = (inp[7]) ? node4374 : node4359;
										assign node4359 = (inp[10]) ? node4367 : node4360;
											assign node4360 = (inp[13]) ? node4364 : node4361;
												assign node4361 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4364 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4367 = (inp[5]) ? node4371 : node4368;
												assign node4368 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4371 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4374 = (inp[15]) ? node4382 : node4375;
											assign node4375 = (inp[13]) ? node4379 : node4376;
												assign node4376 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4379 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4382 = (inp[14]) ? node4386 : node4383;
												assign node4383 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4386 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4389 = (inp[13]) ? node4405 : node4390;
										assign node4390 = (inp[10]) ? node4398 : node4391;
											assign node4391 = (inp[9]) ? node4395 : node4392;
												assign node4392 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4395 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4398 = (inp[15]) ? node4402 : node4399;
												assign node4399 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4402 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4405 = (inp[3]) ? node4413 : node4406;
											assign node4406 = (inp[9]) ? node4410 : node4407;
												assign node4407 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4410 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4413 = (inp[10]) ? node4417 : node4414;
												assign node4414 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4417 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node4420 = (inp[15]) ? node4452 : node4421;
									assign node4421 = (inp[13]) ? node4437 : node4422;
										assign node4422 = (inp[12]) ? node4430 : node4423;
											assign node4423 = (inp[7]) ? node4427 : node4424;
												assign node4424 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4427 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4430 = (inp[3]) ? node4434 : node4431;
												assign node4431 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4434 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4437 = (inp[9]) ? node4445 : node4438;
											assign node4438 = (inp[10]) ? node4442 : node4439;
												assign node4439 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4442 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4445 = (inp[7]) ? node4449 : node4446;
												assign node4446 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4449 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4452 = (inp[3]) ? node4468 : node4453;
										assign node4453 = (inp[7]) ? node4461 : node4454;
											assign node4454 = (inp[13]) ? node4458 : node4455;
												assign node4455 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4458 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4461 = (inp[5]) ? node4465 : node4462;
												assign node4462 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4465 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4468 = (inp[13]) ? node4476 : node4469;
											assign node4469 = (inp[10]) ? node4473 : node4470;
												assign node4470 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4473 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4476 = (inp[10]) ? node4480 : node4477;
												assign node4477 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4480 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4483 = (inp[14]) ? node4547 : node4484;
								assign node4484 = (inp[5]) ? node4516 : node4485;
									assign node4485 = (inp[10]) ? node4501 : node4486;
										assign node4486 = (inp[3]) ? node4494 : node4487;
											assign node4487 = (inp[15]) ? node4491 : node4488;
												assign node4488 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4491 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4494 = (inp[9]) ? node4498 : node4495;
												assign node4495 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4498 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4501 = (inp[15]) ? node4509 : node4502;
											assign node4502 = (inp[12]) ? node4506 : node4503;
												assign node4503 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4506 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4509 = (inp[7]) ? node4513 : node4510;
												assign node4510 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4513 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4516 = (inp[7]) ? node4532 : node4517;
										assign node4517 = (inp[9]) ? node4525 : node4518;
											assign node4518 = (inp[12]) ? node4522 : node4519;
												assign node4519 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4522 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4525 = (inp[2]) ? node4529 : node4526;
												assign node4526 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4529 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4532 = (inp[13]) ? node4540 : node4533;
											assign node4533 = (inp[3]) ? node4537 : node4534;
												assign node4534 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4537 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node4540 = (inp[2]) ? node4544 : node4541;
												assign node4541 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4544 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4547 = (inp[3]) ? node4579 : node4548;
									assign node4548 = (inp[7]) ? node4564 : node4549;
										assign node4549 = (inp[2]) ? node4557 : node4550;
											assign node4550 = (inp[15]) ? node4554 : node4551;
												assign node4551 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4554 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4557 = (inp[10]) ? node4561 : node4558;
												assign node4558 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4561 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4564 = (inp[9]) ? node4572 : node4565;
											assign node4565 = (inp[5]) ? node4569 : node4566;
												assign node4566 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4569 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4572 = (inp[12]) ? node4576 : node4573;
												assign node4573 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4576 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4579 = (inp[5]) ? node4595 : node4580;
										assign node4580 = (inp[7]) ? node4588 : node4581;
											assign node4581 = (inp[13]) ? node4585 : node4582;
												assign node4582 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4585 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4588 = (inp[12]) ? node4592 : node4589;
												assign node4589 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4592 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4595 = (inp[10]) ? node4603 : node4596;
											assign node4596 = (inp[9]) ? node4600 : node4597;
												assign node4597 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4600 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4603 = (inp[13]) ? node4607 : node4604;
												assign node4604 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4607 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node4610 = (inp[14]) ? node4866 : node4611;
						assign node4611 = (inp[9]) ? node4739 : node4612;
							assign node4612 = (inp[7]) ? node4676 : node4613;
								assign node4613 = (inp[4]) ? node4645 : node4614;
									assign node4614 = (inp[2]) ? node4630 : node4615;
										assign node4615 = (inp[12]) ? node4623 : node4616;
											assign node4616 = (inp[8]) ? node4620 : node4617;
												assign node4617 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4620 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4623 = (inp[5]) ? node4627 : node4624;
												assign node4624 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4627 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4630 = (inp[8]) ? node4638 : node4631;
											assign node4631 = (inp[13]) ? node4635 : node4632;
												assign node4632 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4635 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4638 = (inp[3]) ? node4642 : node4639;
												assign node4639 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4642 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4645 = (inp[10]) ? node4661 : node4646;
										assign node4646 = (inp[3]) ? node4654 : node4647;
											assign node4647 = (inp[15]) ? node4651 : node4648;
												assign node4648 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4651 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4654 = (inp[12]) ? node4658 : node4655;
												assign node4655 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4658 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4661 = (inp[5]) ? node4669 : node4662;
											assign node4662 = (inp[2]) ? node4666 : node4663;
												assign node4663 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4666 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4669 = (inp[3]) ? node4673 : node4670;
												assign node4670 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4673 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node4676 = (inp[5]) ? node4708 : node4677;
									assign node4677 = (inp[12]) ? node4693 : node4678;
										assign node4678 = (inp[2]) ? node4686 : node4679;
											assign node4679 = (inp[13]) ? node4683 : node4680;
												assign node4680 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4683 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4686 = (inp[15]) ? node4690 : node4687;
												assign node4687 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4690 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4693 = (inp[8]) ? node4701 : node4694;
											assign node4694 = (inp[15]) ? node4698 : node4695;
												assign node4695 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4698 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4701 = (inp[4]) ? node4705 : node4702;
												assign node4702 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4705 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4708 = (inp[3]) ? node4724 : node4709;
										assign node4709 = (inp[15]) ? node4717 : node4710;
											assign node4710 = (inp[4]) ? node4714 : node4711;
												assign node4711 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4714 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4717 = (inp[10]) ? node4721 : node4718;
												assign node4718 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4721 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4724 = (inp[12]) ? node4732 : node4725;
											assign node4725 = (inp[15]) ? node4729 : node4726;
												assign node4726 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4729 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4732 = (inp[15]) ? node4736 : node4733;
												assign node4733 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4736 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4739 = (inp[12]) ? node4803 : node4740;
								assign node4740 = (inp[3]) ? node4772 : node4741;
									assign node4741 = (inp[13]) ? node4757 : node4742;
										assign node4742 = (inp[7]) ? node4750 : node4743;
											assign node4743 = (inp[8]) ? node4747 : node4744;
												assign node4744 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4747 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4750 = (inp[8]) ? node4754 : node4751;
												assign node4751 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4754 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4757 = (inp[4]) ? node4765 : node4758;
											assign node4758 = (inp[15]) ? node4762 : node4759;
												assign node4759 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4762 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4765 = (inp[5]) ? node4769 : node4766;
												assign node4766 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4769 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4772 = (inp[8]) ? node4788 : node4773;
										assign node4773 = (inp[7]) ? node4781 : node4774;
											assign node4774 = (inp[10]) ? node4778 : node4775;
												assign node4775 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4778 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4781 = (inp[2]) ? node4785 : node4782;
												assign node4782 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4785 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node4788 = (inp[13]) ? node4796 : node4789;
											assign node4789 = (inp[10]) ? node4793 : node4790;
												assign node4790 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4793 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4796 = (inp[2]) ? node4800 : node4797;
												assign node4797 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4800 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4803 = (inp[15]) ? node4835 : node4804;
									assign node4804 = (inp[4]) ? node4820 : node4805;
										assign node4805 = (inp[10]) ? node4813 : node4806;
											assign node4806 = (inp[2]) ? node4810 : node4807;
												assign node4807 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4810 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4813 = (inp[2]) ? node4817 : node4814;
												assign node4814 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4817 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4820 = (inp[8]) ? node4828 : node4821;
											assign node4821 = (inp[10]) ? node4825 : node4822;
												assign node4822 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4825 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4828 = (inp[5]) ? node4832 : node4829;
												assign node4829 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4832 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4835 = (inp[2]) ? node4851 : node4836;
										assign node4836 = (inp[13]) ? node4844 : node4837;
											assign node4837 = (inp[7]) ? node4841 : node4838;
												assign node4838 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4841 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4844 = (inp[4]) ? node4848 : node4845;
												assign node4845 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4848 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4851 = (inp[7]) ? node4859 : node4852;
											assign node4852 = (inp[10]) ? node4856 : node4853;
												assign node4853 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4856 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4859 = (inp[13]) ? node4863 : node4860;
												assign node4860 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4863 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node4866 = (inp[7]) ? node4994 : node4867;
							assign node4867 = (inp[15]) ? node4931 : node4868;
								assign node4868 = (inp[8]) ? node4900 : node4869;
									assign node4869 = (inp[10]) ? node4885 : node4870;
										assign node4870 = (inp[4]) ? node4878 : node4871;
											assign node4871 = (inp[5]) ? node4875 : node4872;
												assign node4872 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4875 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4878 = (inp[3]) ? node4882 : node4879;
												assign node4879 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4882 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4885 = (inp[12]) ? node4893 : node4886;
											assign node4886 = (inp[2]) ? node4890 : node4887;
												assign node4887 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4890 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4893 = (inp[4]) ? node4897 : node4894;
												assign node4894 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4897 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4900 = (inp[3]) ? node4916 : node4901;
										assign node4901 = (inp[5]) ? node4909 : node4902;
											assign node4902 = (inp[9]) ? node4906 : node4903;
												assign node4903 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4906 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4909 = (inp[2]) ? node4913 : node4910;
												assign node4910 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4913 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4916 = (inp[5]) ? node4924 : node4917;
											assign node4917 = (inp[9]) ? node4921 : node4918;
												assign node4918 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4921 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4924 = (inp[9]) ? node4928 : node4925;
												assign node4925 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4928 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4931 = (inp[12]) ? node4963 : node4932;
									assign node4932 = (inp[5]) ? node4948 : node4933;
										assign node4933 = (inp[10]) ? node4941 : node4934;
											assign node4934 = (inp[8]) ? node4938 : node4935;
												assign node4935 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4938 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4941 = (inp[4]) ? node4945 : node4942;
												assign node4942 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4945 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4948 = (inp[2]) ? node4956 : node4949;
											assign node4949 = (inp[13]) ? node4953 : node4950;
												assign node4950 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4953 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4956 = (inp[4]) ? node4960 : node4957;
												assign node4957 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4960 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4963 = (inp[2]) ? node4979 : node4964;
										assign node4964 = (inp[5]) ? node4972 : node4965;
											assign node4965 = (inp[8]) ? node4969 : node4966;
												assign node4966 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4969 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4972 = (inp[3]) ? node4976 : node4973;
												assign node4973 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4976 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4979 = (inp[9]) ? node4987 : node4980;
											assign node4980 = (inp[10]) ? node4984 : node4981;
												assign node4981 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4984 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4987 = (inp[3]) ? node4991 : node4988;
												assign node4988 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4991 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node4994 = (inp[15]) ? node5058 : node4995;
								assign node4995 = (inp[2]) ? node5027 : node4996;
									assign node4996 = (inp[5]) ? node5012 : node4997;
										assign node4997 = (inp[13]) ? node5005 : node4998;
											assign node4998 = (inp[4]) ? node5002 : node4999;
												assign node4999 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5002 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5005 = (inp[12]) ? node5009 : node5006;
												assign node5006 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5009 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5012 = (inp[9]) ? node5020 : node5013;
											assign node5013 = (inp[4]) ? node5017 : node5014;
												assign node5014 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5017 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5020 = (inp[3]) ? node5024 : node5021;
												assign node5021 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5024 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5027 = (inp[5]) ? node5043 : node5028;
										assign node5028 = (inp[9]) ? node5036 : node5029;
											assign node5029 = (inp[10]) ? node5033 : node5030;
												assign node5030 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5033 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5036 = (inp[8]) ? node5040 : node5037;
												assign node5037 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5040 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5043 = (inp[3]) ? node5051 : node5044;
											assign node5044 = (inp[12]) ? node5048 : node5045;
												assign node5045 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5048 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5051 = (inp[13]) ? node5055 : node5052;
												assign node5052 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5055 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5058 = (inp[3]) ? node5090 : node5059;
									assign node5059 = (inp[10]) ? node5075 : node5060;
										assign node5060 = (inp[12]) ? node5068 : node5061;
											assign node5061 = (inp[13]) ? node5065 : node5062;
												assign node5062 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5065 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5068 = (inp[4]) ? node5072 : node5069;
												assign node5069 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5072 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5075 = (inp[13]) ? node5083 : node5076;
											assign node5076 = (inp[8]) ? node5080 : node5077;
												assign node5077 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5080 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5083 = (inp[5]) ? node5087 : node5084;
												assign node5084 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5087 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5090 = (inp[2]) ? node5106 : node5091;
										assign node5091 = (inp[13]) ? node5099 : node5092;
											assign node5092 = (inp[4]) ? node5096 : node5093;
												assign node5093 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5096 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5099 = (inp[9]) ? node5103 : node5100;
												assign node5100 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5103 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5106 = (inp[13]) ? node5114 : node5107;
											assign node5107 = (inp[5]) ? node5111 : node5108;
												assign node5108 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5111 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5114 = (inp[5]) ? node5118 : node5115;
												assign node5115 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5118 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
				assign node5121 = (inp[13]) ? node5633 : node5122;
					assign node5122 = (inp[3]) ? node5378 : node5123;
						assign node5123 = (inp[5]) ? node5251 : node5124;
							assign node5124 = (inp[10]) ? node5188 : node5125;
								assign node5125 = (inp[4]) ? node5157 : node5126;
									assign node5126 = (inp[15]) ? node5142 : node5127;
										assign node5127 = (inp[7]) ? node5135 : node5128;
											assign node5128 = (inp[8]) ? node5132 : node5129;
												assign node5129 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node5132 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node5135 = (inp[2]) ? node5139 : node5136;
												assign node5136 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5139 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node5142 = (inp[14]) ? node5150 : node5143;
											assign node5143 = (inp[11]) ? node5147 : node5144;
												assign node5144 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5147 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5150 = (inp[2]) ? node5154 : node5151;
												assign node5151 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5154 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node5157 = (inp[9]) ? node5173 : node5158;
										assign node5158 = (inp[7]) ? node5166 : node5159;
											assign node5159 = (inp[15]) ? node5163 : node5160;
												assign node5160 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5163 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5166 = (inp[8]) ? node5170 : node5167;
												assign node5167 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5170 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5173 = (inp[14]) ? node5181 : node5174;
											assign node5174 = (inp[8]) ? node5178 : node5175;
												assign node5175 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5178 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5181 = (inp[7]) ? node5185 : node5182;
												assign node5182 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5185 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node5188 = (inp[12]) ? node5220 : node5189;
									assign node5189 = (inp[8]) ? node5205 : node5190;
										assign node5190 = (inp[4]) ? node5198 : node5191;
											assign node5191 = (inp[15]) ? node5195 : node5192;
												assign node5192 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5195 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5198 = (inp[2]) ? node5202 : node5199;
												assign node5199 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5202 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5205 = (inp[9]) ? node5213 : node5206;
											assign node5206 = (inp[11]) ? node5210 : node5207;
												assign node5207 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5210 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5213 = (inp[11]) ? node5217 : node5214;
												assign node5214 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5217 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5220 = (inp[4]) ? node5236 : node5221;
										assign node5221 = (inp[11]) ? node5229 : node5222;
											assign node5222 = (inp[8]) ? node5226 : node5223;
												assign node5223 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5226 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5229 = (inp[15]) ? node5233 : node5230;
												assign node5230 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5233 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5236 = (inp[15]) ? node5244 : node5237;
											assign node5237 = (inp[9]) ? node5241 : node5238;
												assign node5238 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5241 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5244 = (inp[8]) ? node5248 : node5245;
												assign node5245 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5248 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node5251 = (inp[7]) ? node5315 : node5252;
								assign node5252 = (inp[11]) ? node5284 : node5253;
									assign node5253 = (inp[2]) ? node5269 : node5254;
										assign node5254 = (inp[4]) ? node5262 : node5255;
											assign node5255 = (inp[12]) ? node5259 : node5256;
												assign node5256 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5259 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5262 = (inp[10]) ? node5266 : node5263;
												assign node5263 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5266 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5269 = (inp[10]) ? node5277 : node5270;
											assign node5270 = (inp[4]) ? node5274 : node5271;
												assign node5271 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5274 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5277 = (inp[15]) ? node5281 : node5278;
												assign node5278 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5281 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5284 = (inp[4]) ? node5300 : node5285;
										assign node5285 = (inp[10]) ? node5293 : node5286;
											assign node5286 = (inp[2]) ? node5290 : node5287;
												assign node5287 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5290 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5293 = (inp[9]) ? node5297 : node5294;
												assign node5294 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5297 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5300 = (inp[2]) ? node5308 : node5301;
											assign node5301 = (inp[10]) ? node5305 : node5302;
												assign node5302 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5305 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5308 = (inp[8]) ? node5312 : node5309;
												assign node5309 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5312 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5315 = (inp[9]) ? node5347 : node5316;
									assign node5316 = (inp[10]) ? node5332 : node5317;
										assign node5317 = (inp[14]) ? node5325 : node5318;
											assign node5318 = (inp[8]) ? node5322 : node5319;
												assign node5319 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5322 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5325 = (inp[4]) ? node5329 : node5326;
												assign node5326 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5329 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5332 = (inp[8]) ? node5340 : node5333;
											assign node5333 = (inp[4]) ? node5337 : node5334;
												assign node5334 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5337 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5340 = (inp[4]) ? node5344 : node5341;
												assign node5341 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5344 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5347 = (inp[10]) ? node5363 : node5348;
										assign node5348 = (inp[2]) ? node5356 : node5349;
											assign node5349 = (inp[4]) ? node5353 : node5350;
												assign node5350 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5353 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5356 = (inp[11]) ? node5360 : node5357;
												assign node5357 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5360 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5363 = (inp[15]) ? node5371 : node5364;
											assign node5364 = (inp[12]) ? node5368 : node5365;
												assign node5365 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5368 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5371 = (inp[14]) ? node5375 : node5372;
												assign node5372 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5375 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node5378 = (inp[12]) ? node5506 : node5379;
							assign node5379 = (inp[11]) ? node5443 : node5380;
								assign node5380 = (inp[8]) ? node5412 : node5381;
									assign node5381 = (inp[5]) ? node5397 : node5382;
										assign node5382 = (inp[7]) ? node5390 : node5383;
											assign node5383 = (inp[9]) ? node5387 : node5384;
												assign node5384 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5387 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5390 = (inp[10]) ? node5394 : node5391;
												assign node5391 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5394 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5397 = (inp[2]) ? node5405 : node5398;
											assign node5398 = (inp[7]) ? node5402 : node5399;
												assign node5399 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5402 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5405 = (inp[15]) ? node5409 : node5406;
												assign node5406 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5409 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5412 = (inp[7]) ? node5428 : node5413;
										assign node5413 = (inp[9]) ? node5421 : node5414;
											assign node5414 = (inp[15]) ? node5418 : node5415;
												assign node5415 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5418 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5421 = (inp[4]) ? node5425 : node5422;
												assign node5422 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5425 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5428 = (inp[14]) ? node5436 : node5429;
											assign node5429 = (inp[2]) ? node5433 : node5430;
												assign node5430 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5433 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5436 = (inp[5]) ? node5440 : node5437;
												assign node5437 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5440 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5443 = (inp[14]) ? node5475 : node5444;
									assign node5444 = (inp[4]) ? node5460 : node5445;
										assign node5445 = (inp[7]) ? node5453 : node5446;
											assign node5446 = (inp[9]) ? node5450 : node5447;
												assign node5447 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5450 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5453 = (inp[5]) ? node5457 : node5454;
												assign node5454 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5457 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5460 = (inp[8]) ? node5468 : node5461;
											assign node5461 = (inp[15]) ? node5465 : node5462;
												assign node5462 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5465 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5468 = (inp[2]) ? node5472 : node5469;
												assign node5469 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5472 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node5475 = (inp[4]) ? node5491 : node5476;
										assign node5476 = (inp[8]) ? node5484 : node5477;
											assign node5477 = (inp[10]) ? node5481 : node5478;
												assign node5478 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5481 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5484 = (inp[9]) ? node5488 : node5485;
												assign node5485 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5488 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5491 = (inp[15]) ? node5499 : node5492;
											assign node5492 = (inp[9]) ? node5496 : node5493;
												assign node5493 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5496 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5499 = (inp[7]) ? node5503 : node5500;
												assign node5500 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5503 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node5506 = (inp[15]) ? node5570 : node5507;
								assign node5507 = (inp[5]) ? node5539 : node5508;
									assign node5508 = (inp[8]) ? node5524 : node5509;
										assign node5509 = (inp[4]) ? node5517 : node5510;
											assign node5510 = (inp[10]) ? node5514 : node5511;
												assign node5511 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5514 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5517 = (inp[7]) ? node5521 : node5518;
												assign node5518 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5521 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5524 = (inp[14]) ? node5532 : node5525;
											assign node5525 = (inp[10]) ? node5529 : node5526;
												assign node5526 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5529 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5532 = (inp[9]) ? node5536 : node5533;
												assign node5533 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5536 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5539 = (inp[7]) ? node5555 : node5540;
										assign node5540 = (inp[9]) ? node5548 : node5541;
											assign node5541 = (inp[10]) ? node5545 : node5542;
												assign node5542 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5545 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5548 = (inp[4]) ? node5552 : node5549;
												assign node5549 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5552 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5555 = (inp[9]) ? node5563 : node5556;
											assign node5556 = (inp[8]) ? node5560 : node5557;
												assign node5557 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5560 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5563 = (inp[11]) ? node5567 : node5564;
												assign node5564 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5567 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5570 = (inp[7]) ? node5602 : node5571;
									assign node5571 = (inp[14]) ? node5587 : node5572;
										assign node5572 = (inp[11]) ? node5580 : node5573;
											assign node5573 = (inp[2]) ? node5577 : node5574;
												assign node5574 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5577 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5580 = (inp[10]) ? node5584 : node5581;
												assign node5581 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5584 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5587 = (inp[2]) ? node5595 : node5588;
											assign node5588 = (inp[8]) ? node5592 : node5589;
												assign node5589 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5592 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5595 = (inp[9]) ? node5599 : node5596;
												assign node5596 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5599 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5602 = (inp[8]) ? node5618 : node5603;
										assign node5603 = (inp[4]) ? node5611 : node5604;
											assign node5604 = (inp[11]) ? node5608 : node5605;
												assign node5605 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5608 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5611 = (inp[14]) ? node5615 : node5612;
												assign node5612 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5615 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5618 = (inp[9]) ? node5626 : node5619;
											assign node5619 = (inp[10]) ? node5623 : node5620;
												assign node5620 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5623 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5626 = (inp[10]) ? node5630 : node5627;
												assign node5627 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5630 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node5633 = (inp[9]) ? node5889 : node5634;
						assign node5634 = (inp[2]) ? node5762 : node5635;
							assign node5635 = (inp[4]) ? node5699 : node5636;
								assign node5636 = (inp[5]) ? node5668 : node5637;
									assign node5637 = (inp[3]) ? node5653 : node5638;
										assign node5638 = (inp[8]) ? node5646 : node5639;
											assign node5639 = (inp[14]) ? node5643 : node5640;
												assign node5640 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5643 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5646 = (inp[11]) ? node5650 : node5647;
												assign node5647 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5650 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5653 = (inp[12]) ? node5661 : node5654;
											assign node5654 = (inp[11]) ? node5658 : node5655;
												assign node5655 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5658 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5661 = (inp[11]) ? node5665 : node5662;
												assign node5662 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5665 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5668 = (inp[8]) ? node5684 : node5669;
										assign node5669 = (inp[11]) ? node5677 : node5670;
											assign node5670 = (inp[15]) ? node5674 : node5671;
												assign node5671 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5674 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5677 = (inp[10]) ? node5681 : node5678;
												assign node5678 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5681 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5684 = (inp[12]) ? node5692 : node5685;
											assign node5685 = (inp[10]) ? node5689 : node5686;
												assign node5686 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5689 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5692 = (inp[10]) ? node5696 : node5693;
												assign node5693 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5696 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5699 = (inp[14]) ? node5731 : node5700;
									assign node5700 = (inp[5]) ? node5716 : node5701;
										assign node5701 = (inp[7]) ? node5709 : node5702;
											assign node5702 = (inp[10]) ? node5706 : node5703;
												assign node5703 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5706 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5709 = (inp[11]) ? node5713 : node5710;
												assign node5710 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5713 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5716 = (inp[8]) ? node5724 : node5717;
											assign node5717 = (inp[12]) ? node5721 : node5718;
												assign node5718 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5721 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5724 = (inp[15]) ? node5728 : node5725;
												assign node5725 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5728 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5731 = (inp[10]) ? node5747 : node5732;
										assign node5732 = (inp[5]) ? node5740 : node5733;
											assign node5733 = (inp[8]) ? node5737 : node5734;
												assign node5734 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5737 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5740 = (inp[8]) ? node5744 : node5741;
												assign node5741 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5744 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5747 = (inp[15]) ? node5755 : node5748;
											assign node5748 = (inp[5]) ? node5752 : node5749;
												assign node5749 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5752 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5755 = (inp[7]) ? node5759 : node5756;
												assign node5756 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5759 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node5762 = (inp[8]) ? node5826 : node5763;
								assign node5763 = (inp[10]) ? node5795 : node5764;
									assign node5764 = (inp[15]) ? node5780 : node5765;
										assign node5765 = (inp[3]) ? node5773 : node5766;
											assign node5766 = (inp[5]) ? node5770 : node5767;
												assign node5767 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5770 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5773 = (inp[14]) ? node5777 : node5774;
												assign node5774 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5777 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5780 = (inp[3]) ? node5788 : node5781;
											assign node5781 = (inp[14]) ? node5785 : node5782;
												assign node5782 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5785 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5788 = (inp[5]) ? node5792 : node5789;
												assign node5789 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5792 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5795 = (inp[4]) ? node5811 : node5796;
										assign node5796 = (inp[11]) ? node5804 : node5797;
											assign node5797 = (inp[12]) ? node5801 : node5798;
												assign node5798 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5801 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5804 = (inp[3]) ? node5808 : node5805;
												assign node5805 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5808 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5811 = (inp[14]) ? node5819 : node5812;
											assign node5812 = (inp[7]) ? node5816 : node5813;
												assign node5813 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5816 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5819 = (inp[5]) ? node5823 : node5820;
												assign node5820 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5823 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5826 = (inp[3]) ? node5858 : node5827;
									assign node5827 = (inp[10]) ? node5843 : node5828;
										assign node5828 = (inp[15]) ? node5836 : node5829;
											assign node5829 = (inp[14]) ? node5833 : node5830;
												assign node5830 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5833 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5836 = (inp[7]) ? node5840 : node5837;
												assign node5837 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5840 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5843 = (inp[15]) ? node5851 : node5844;
											assign node5844 = (inp[4]) ? node5848 : node5845;
												assign node5845 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5848 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5851 = (inp[11]) ? node5855 : node5852;
												assign node5852 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5855 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5858 = (inp[12]) ? node5874 : node5859;
										assign node5859 = (inp[14]) ? node5867 : node5860;
											assign node5860 = (inp[4]) ? node5864 : node5861;
												assign node5861 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5864 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5867 = (inp[5]) ? node5871 : node5868;
												assign node5868 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5871 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5874 = (inp[4]) ? node5882 : node5875;
											assign node5875 = (inp[14]) ? node5879 : node5876;
												assign node5876 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5879 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5882 = (inp[14]) ? node5886 : node5883;
												assign node5883 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5886 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node5889 = (inp[12]) ? node6017 : node5890;
							assign node5890 = (inp[7]) ? node5954 : node5891;
								assign node5891 = (inp[4]) ? node5923 : node5892;
									assign node5892 = (inp[8]) ? node5908 : node5893;
										assign node5893 = (inp[15]) ? node5901 : node5894;
											assign node5894 = (inp[11]) ? node5898 : node5895;
												assign node5895 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5898 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5901 = (inp[14]) ? node5905 : node5902;
												assign node5902 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5905 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5908 = (inp[14]) ? node5916 : node5909;
											assign node5909 = (inp[10]) ? node5913 : node5910;
												assign node5910 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5913 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5916 = (inp[2]) ? node5920 : node5917;
												assign node5917 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5920 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node5923 = (inp[3]) ? node5939 : node5924;
										assign node5924 = (inp[2]) ? node5932 : node5925;
											assign node5925 = (inp[14]) ? node5929 : node5926;
												assign node5926 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5929 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5932 = (inp[8]) ? node5936 : node5933;
												assign node5933 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5936 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5939 = (inp[5]) ? node5947 : node5940;
											assign node5940 = (inp[14]) ? node5944 : node5941;
												assign node5941 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5944 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5947 = (inp[15]) ? node5951 : node5948;
												assign node5948 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5951 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5954 = (inp[11]) ? node5986 : node5955;
									assign node5955 = (inp[4]) ? node5971 : node5956;
										assign node5956 = (inp[10]) ? node5964 : node5957;
											assign node5957 = (inp[15]) ? node5961 : node5958;
												assign node5958 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5961 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5964 = (inp[15]) ? node5968 : node5965;
												assign node5965 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5968 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5971 = (inp[14]) ? node5979 : node5972;
											assign node5972 = (inp[8]) ? node5976 : node5973;
												assign node5973 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5976 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5979 = (inp[8]) ? node5983 : node5980;
												assign node5980 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5983 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5986 = (inp[10]) ? node6002 : node5987;
										assign node5987 = (inp[14]) ? node5995 : node5988;
											assign node5988 = (inp[15]) ? node5992 : node5989;
												assign node5989 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5992 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5995 = (inp[2]) ? node5999 : node5996;
												assign node5996 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5999 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6002 = (inp[5]) ? node6010 : node6003;
											assign node6003 = (inp[15]) ? node6007 : node6004;
												assign node6004 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6007 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6010 = (inp[4]) ? node6014 : node6011;
												assign node6011 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6014 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node6017 = (inp[11]) ? node6081 : node6018;
								assign node6018 = (inp[8]) ? node6050 : node6019;
									assign node6019 = (inp[7]) ? node6035 : node6020;
										assign node6020 = (inp[15]) ? node6028 : node6021;
											assign node6021 = (inp[14]) ? node6025 : node6022;
												assign node6022 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6025 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6028 = (inp[3]) ? node6032 : node6029;
												assign node6029 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6032 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6035 = (inp[2]) ? node6043 : node6036;
											assign node6036 = (inp[3]) ? node6040 : node6037;
												assign node6037 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6040 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6043 = (inp[10]) ? node6047 : node6044;
												assign node6044 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6047 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node6050 = (inp[7]) ? node6066 : node6051;
										assign node6051 = (inp[15]) ? node6059 : node6052;
											assign node6052 = (inp[10]) ? node6056 : node6053;
												assign node6053 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6056 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6059 = (inp[10]) ? node6063 : node6060;
												assign node6060 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6063 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6066 = (inp[4]) ? node6074 : node6067;
											assign node6067 = (inp[15]) ? node6071 : node6068;
												assign node6068 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6071 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6074 = (inp[3]) ? node6078 : node6075;
												assign node6075 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6078 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node6081 = (inp[15]) ? node6113 : node6082;
									assign node6082 = (inp[10]) ? node6098 : node6083;
										assign node6083 = (inp[14]) ? node6091 : node6084;
											assign node6084 = (inp[7]) ? node6088 : node6085;
												assign node6085 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6088 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6091 = (inp[3]) ? node6095 : node6092;
												assign node6092 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6095 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6098 = (inp[4]) ? node6106 : node6099;
											assign node6099 = (inp[7]) ? node6103 : node6100;
												assign node6100 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6103 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6106 = (inp[14]) ? node6110 : node6107;
												assign node6107 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6110 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000011111;
									assign node6113 = (inp[2]) ? node6129 : node6114;
										assign node6114 = (inp[3]) ? node6122 : node6115;
											assign node6115 = (inp[4]) ? node6119 : node6116;
												assign node6116 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6119 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6122 = (inp[7]) ? node6126 : node6123;
												assign node6123 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6126 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node6129 = (inp[5]) ? node6137 : node6130;
											assign node6130 = (inp[4]) ? node6134 : node6131;
												assign node6131 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6134 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node6137 = (inp[7]) ? node6141 : node6138;
												assign node6138 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node6141 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
			assign node6144 = (inp[2]) ? node7168 : node6145;
				assign node6145 = (inp[13]) ? node6657 : node6146;
					assign node6146 = (inp[12]) ? node6402 : node6147;
						assign node6147 = (inp[3]) ? node6275 : node6148;
							assign node6148 = (inp[15]) ? node6212 : node6149;
								assign node6149 = (inp[11]) ? node6181 : node6150;
									assign node6150 = (inp[14]) ? node6166 : node6151;
										assign node6151 = (inp[5]) ? node6159 : node6152;
											assign node6152 = (inp[4]) ? node6156 : node6153;
												assign node6153 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node6156 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6159 = (inp[10]) ? node6163 : node6160;
												assign node6160 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6163 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node6166 = (inp[7]) ? node6174 : node6167;
											assign node6167 = (inp[5]) ? node6171 : node6168;
												assign node6168 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6171 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6174 = (inp[9]) ? node6178 : node6175;
												assign node6175 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6178 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6181 = (inp[9]) ? node6197 : node6182;
										assign node6182 = (inp[8]) ? node6190 : node6183;
											assign node6183 = (inp[5]) ? node6187 : node6184;
												assign node6184 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6187 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6190 = (inp[0]) ? node6194 : node6191;
												assign node6191 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6194 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6197 = (inp[7]) ? node6205 : node6198;
											assign node6198 = (inp[8]) ? node6202 : node6199;
												assign node6199 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6202 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6205 = (inp[10]) ? node6209 : node6206;
												assign node6206 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6209 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node6212 = (inp[0]) ? node6244 : node6213;
									assign node6213 = (inp[10]) ? node6229 : node6214;
										assign node6214 = (inp[5]) ? node6222 : node6215;
											assign node6215 = (inp[14]) ? node6219 : node6216;
												assign node6216 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6219 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6222 = (inp[4]) ? node6226 : node6223;
												assign node6223 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6226 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6229 = (inp[11]) ? node6237 : node6230;
											assign node6230 = (inp[9]) ? node6234 : node6231;
												assign node6231 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6234 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6237 = (inp[14]) ? node6241 : node6238;
												assign node6238 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6241 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6244 = (inp[10]) ? node6260 : node6245;
										assign node6245 = (inp[14]) ? node6253 : node6246;
											assign node6246 = (inp[11]) ? node6250 : node6247;
												assign node6247 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6250 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6253 = (inp[4]) ? node6257 : node6254;
												assign node6254 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6257 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6260 = (inp[7]) ? node6268 : node6261;
											assign node6261 = (inp[9]) ? node6265 : node6262;
												assign node6262 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6265 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6268 = (inp[5]) ? node6272 : node6269;
												assign node6269 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6272 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
							assign node6275 = (inp[11]) ? node6339 : node6276;
								assign node6276 = (inp[5]) ? node6308 : node6277;
									assign node6277 = (inp[10]) ? node6293 : node6278;
										assign node6278 = (inp[7]) ? node6286 : node6279;
											assign node6279 = (inp[15]) ? node6283 : node6280;
												assign node6280 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6283 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6286 = (inp[0]) ? node6290 : node6287;
												assign node6287 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6290 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6293 = (inp[8]) ? node6301 : node6294;
											assign node6294 = (inp[14]) ? node6298 : node6295;
												assign node6295 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6298 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6301 = (inp[15]) ? node6305 : node6302;
												assign node6302 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node6305 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6308 = (inp[15]) ? node6324 : node6309;
										assign node6309 = (inp[8]) ? node6317 : node6310;
											assign node6310 = (inp[0]) ? node6314 : node6311;
												assign node6311 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6314 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6317 = (inp[9]) ? node6321 : node6318;
												assign node6318 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6321 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6324 = (inp[8]) ? node6332 : node6325;
											assign node6325 = (inp[0]) ? node6329 : node6326;
												assign node6326 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6329 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6332 = (inp[7]) ? node6336 : node6333;
												assign node6333 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6336 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node6339 = (inp[15]) ? node6371 : node6340;
									assign node6340 = (inp[14]) ? node6356 : node6341;
										assign node6341 = (inp[4]) ? node6349 : node6342;
											assign node6342 = (inp[7]) ? node6346 : node6343;
												assign node6343 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6346 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6349 = (inp[10]) ? node6353 : node6350;
												assign node6350 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6353 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6356 = (inp[7]) ? node6364 : node6357;
											assign node6357 = (inp[8]) ? node6361 : node6358;
												assign node6358 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6361 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6364 = (inp[0]) ? node6368 : node6365;
												assign node6365 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6368 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6371 = (inp[10]) ? node6387 : node6372;
										assign node6372 = (inp[4]) ? node6380 : node6373;
											assign node6373 = (inp[9]) ? node6377 : node6374;
												assign node6374 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6377 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6380 = (inp[14]) ? node6384 : node6381;
												assign node6381 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6384 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6387 = (inp[5]) ? node6395 : node6388;
											assign node6388 = (inp[0]) ? node6392 : node6389;
												assign node6389 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6392 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6395 = (inp[4]) ? node6399 : node6396;
												assign node6396 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6399 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node6402 = (inp[15]) ? node6530 : node6403;
							assign node6403 = (inp[8]) ? node6467 : node6404;
								assign node6404 = (inp[9]) ? node6436 : node6405;
									assign node6405 = (inp[0]) ? node6421 : node6406;
										assign node6406 = (inp[10]) ? node6414 : node6407;
											assign node6407 = (inp[14]) ? node6411 : node6408;
												assign node6408 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6411 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6414 = (inp[4]) ? node6418 : node6415;
												assign node6415 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6418 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6421 = (inp[5]) ? node6429 : node6422;
											assign node6422 = (inp[4]) ? node6426 : node6423;
												assign node6423 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6426 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6429 = (inp[10]) ? node6433 : node6430;
												assign node6430 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6433 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6436 = (inp[4]) ? node6452 : node6437;
										assign node6437 = (inp[14]) ? node6445 : node6438;
											assign node6438 = (inp[11]) ? node6442 : node6439;
												assign node6439 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6442 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6445 = (inp[7]) ? node6449 : node6446;
												assign node6446 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6449 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6452 = (inp[3]) ? node6460 : node6453;
											assign node6453 = (inp[11]) ? node6457 : node6454;
												assign node6454 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6457 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6460 = (inp[5]) ? node6464 : node6461;
												assign node6461 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6464 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node6467 = (inp[11]) ? node6499 : node6468;
									assign node6468 = (inp[4]) ? node6484 : node6469;
										assign node6469 = (inp[5]) ? node6477 : node6470;
											assign node6470 = (inp[3]) ? node6474 : node6471;
												assign node6471 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6474 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6477 = (inp[10]) ? node6481 : node6478;
												assign node6478 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6481 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6484 = (inp[7]) ? node6492 : node6485;
											assign node6485 = (inp[3]) ? node6489 : node6486;
												assign node6486 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6489 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6492 = (inp[9]) ? node6496 : node6493;
												assign node6493 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6496 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6499 = (inp[0]) ? node6515 : node6500;
										assign node6500 = (inp[9]) ? node6508 : node6501;
											assign node6501 = (inp[14]) ? node6505 : node6502;
												assign node6502 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6505 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6508 = (inp[14]) ? node6512 : node6509;
												assign node6509 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6512 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6515 = (inp[9]) ? node6523 : node6516;
											assign node6516 = (inp[4]) ? node6520 : node6517;
												assign node6517 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6520 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6523 = (inp[14]) ? node6527 : node6524;
												assign node6524 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6527 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node6530 = (inp[7]) ? node6594 : node6531;
								assign node6531 = (inp[4]) ? node6563 : node6532;
									assign node6532 = (inp[8]) ? node6548 : node6533;
										assign node6533 = (inp[14]) ? node6541 : node6534;
											assign node6534 = (inp[11]) ? node6538 : node6535;
												assign node6535 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6538 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6541 = (inp[3]) ? node6545 : node6542;
												assign node6542 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6545 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6548 = (inp[5]) ? node6556 : node6549;
											assign node6549 = (inp[14]) ? node6553 : node6550;
												assign node6550 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6553 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node6556 = (inp[0]) ? node6560 : node6557;
												assign node6557 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6560 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6563 = (inp[11]) ? node6579 : node6564;
										assign node6564 = (inp[14]) ? node6572 : node6565;
											assign node6565 = (inp[3]) ? node6569 : node6566;
												assign node6566 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6569 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6572 = (inp[5]) ? node6576 : node6573;
												assign node6573 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6576 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6579 = (inp[9]) ? node6587 : node6580;
											assign node6580 = (inp[5]) ? node6584 : node6581;
												assign node6581 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6584 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6587 = (inp[0]) ? node6591 : node6588;
												assign node6588 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6591 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node6594 = (inp[14]) ? node6626 : node6595;
									assign node6595 = (inp[3]) ? node6611 : node6596;
										assign node6596 = (inp[8]) ? node6604 : node6597;
											assign node6597 = (inp[4]) ? node6601 : node6598;
												assign node6598 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6601 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6604 = (inp[9]) ? node6608 : node6605;
												assign node6605 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6608 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6611 = (inp[0]) ? node6619 : node6612;
											assign node6612 = (inp[11]) ? node6616 : node6613;
												assign node6613 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6616 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6619 = (inp[10]) ? node6623 : node6620;
												assign node6620 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6623 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node6626 = (inp[5]) ? node6642 : node6627;
										assign node6627 = (inp[0]) ? node6635 : node6628;
											assign node6628 = (inp[9]) ? node6632 : node6629;
												assign node6629 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6632 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6635 = (inp[4]) ? node6639 : node6636;
												assign node6636 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6639 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6642 = (inp[8]) ? node6650 : node6643;
											assign node6643 = (inp[0]) ? node6647 : node6644;
												assign node6644 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6647 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6650 = (inp[11]) ? node6654 : node6651;
												assign node6651 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6654 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node6657 = (inp[10]) ? node6913 : node6658;
						assign node6658 = (inp[0]) ? node6786 : node6659;
							assign node6659 = (inp[12]) ? node6723 : node6660;
								assign node6660 = (inp[9]) ? node6692 : node6661;
									assign node6661 = (inp[5]) ? node6677 : node6662;
										assign node6662 = (inp[15]) ? node6670 : node6663;
											assign node6663 = (inp[11]) ? node6667 : node6664;
												assign node6664 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6667 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6670 = (inp[11]) ? node6674 : node6671;
												assign node6671 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6674 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6677 = (inp[7]) ? node6685 : node6678;
											assign node6678 = (inp[8]) ? node6682 : node6679;
												assign node6679 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6682 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6685 = (inp[14]) ? node6689 : node6686;
												assign node6686 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6689 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6692 = (inp[8]) ? node6708 : node6693;
										assign node6693 = (inp[14]) ? node6701 : node6694;
											assign node6694 = (inp[4]) ? node6698 : node6695;
												assign node6695 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6698 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6701 = (inp[5]) ? node6705 : node6702;
												assign node6702 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6705 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6708 = (inp[14]) ? node6716 : node6709;
											assign node6709 = (inp[3]) ? node6713 : node6710;
												assign node6710 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6713 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6716 = (inp[3]) ? node6720 : node6717;
												assign node6717 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6720 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node6723 = (inp[15]) ? node6755 : node6724;
									assign node6724 = (inp[9]) ? node6740 : node6725;
										assign node6725 = (inp[8]) ? node6733 : node6726;
											assign node6726 = (inp[3]) ? node6730 : node6727;
												assign node6727 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6730 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6733 = (inp[5]) ? node6737 : node6734;
												assign node6734 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6737 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6740 = (inp[7]) ? node6748 : node6741;
											assign node6741 = (inp[8]) ? node6745 : node6742;
												assign node6742 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6745 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6748 = (inp[11]) ? node6752 : node6749;
												assign node6749 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6752 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6755 = (inp[5]) ? node6771 : node6756;
										assign node6756 = (inp[7]) ? node6764 : node6757;
											assign node6757 = (inp[14]) ? node6761 : node6758;
												assign node6758 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6761 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6764 = (inp[3]) ? node6768 : node6765;
												assign node6765 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6768 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6771 = (inp[4]) ? node6779 : node6772;
											assign node6772 = (inp[9]) ? node6776 : node6773;
												assign node6773 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6776 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6779 = (inp[7]) ? node6783 : node6780;
												assign node6780 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6783 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node6786 = (inp[4]) ? node6850 : node6787;
								assign node6787 = (inp[12]) ? node6819 : node6788;
									assign node6788 = (inp[15]) ? node6804 : node6789;
										assign node6789 = (inp[7]) ? node6797 : node6790;
											assign node6790 = (inp[11]) ? node6794 : node6791;
												assign node6791 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6794 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6797 = (inp[9]) ? node6801 : node6798;
												assign node6798 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6801 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6804 = (inp[3]) ? node6812 : node6805;
											assign node6805 = (inp[8]) ? node6809 : node6806;
												assign node6806 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6809 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6812 = (inp[8]) ? node6816 : node6813;
												assign node6813 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6816 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6819 = (inp[14]) ? node6835 : node6820;
										assign node6820 = (inp[5]) ? node6828 : node6821;
											assign node6821 = (inp[8]) ? node6825 : node6822;
												assign node6822 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6825 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6828 = (inp[11]) ? node6832 : node6829;
												assign node6829 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6832 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6835 = (inp[9]) ? node6843 : node6836;
											assign node6836 = (inp[7]) ? node6840 : node6837;
												assign node6837 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6840 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6843 = (inp[15]) ? node6847 : node6844;
												assign node6844 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6847 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node6850 = (inp[5]) ? node6882 : node6851;
									assign node6851 = (inp[9]) ? node6867 : node6852;
										assign node6852 = (inp[12]) ? node6860 : node6853;
											assign node6853 = (inp[8]) ? node6857 : node6854;
												assign node6854 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6857 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6860 = (inp[8]) ? node6864 : node6861;
												assign node6861 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6864 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6867 = (inp[15]) ? node6875 : node6868;
											assign node6868 = (inp[11]) ? node6872 : node6869;
												assign node6869 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6872 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6875 = (inp[7]) ? node6879 : node6876;
												assign node6876 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6879 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node6882 = (inp[14]) ? node6898 : node6883;
										assign node6883 = (inp[3]) ? node6891 : node6884;
											assign node6884 = (inp[11]) ? node6888 : node6885;
												assign node6885 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6888 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6891 = (inp[15]) ? node6895 : node6892;
												assign node6892 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6895 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6898 = (inp[8]) ? node6906 : node6899;
											assign node6899 = (inp[11]) ? node6903 : node6900;
												assign node6900 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6903 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6906 = (inp[9]) ? node6910 : node6907;
												assign node6907 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node6910 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node6913 = (inp[14]) ? node7041 : node6914;
							assign node6914 = (inp[5]) ? node6978 : node6915;
								assign node6915 = (inp[9]) ? node6947 : node6916;
									assign node6916 = (inp[8]) ? node6932 : node6917;
										assign node6917 = (inp[4]) ? node6925 : node6918;
											assign node6918 = (inp[7]) ? node6922 : node6919;
												assign node6919 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6922 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6925 = (inp[7]) ? node6929 : node6926;
												assign node6926 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6929 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6932 = (inp[15]) ? node6940 : node6933;
											assign node6933 = (inp[7]) ? node6937 : node6934;
												assign node6934 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6937 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6940 = (inp[0]) ? node6944 : node6941;
												assign node6941 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6944 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6947 = (inp[8]) ? node6963 : node6948;
										assign node6948 = (inp[3]) ? node6956 : node6949;
											assign node6949 = (inp[15]) ? node6953 : node6950;
												assign node6950 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6953 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6956 = (inp[12]) ? node6960 : node6957;
												assign node6957 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6960 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6963 = (inp[12]) ? node6971 : node6964;
											assign node6964 = (inp[11]) ? node6968 : node6965;
												assign node6965 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6968 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6971 = (inp[0]) ? node6975 : node6972;
												assign node6972 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6975 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
								assign node6978 = (inp[7]) ? node7010 : node6979;
									assign node6979 = (inp[12]) ? node6995 : node6980;
										assign node6980 = (inp[8]) ? node6988 : node6981;
											assign node6981 = (inp[3]) ? node6985 : node6982;
												assign node6982 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6985 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6988 = (inp[4]) ? node6992 : node6989;
												assign node6989 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6992 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6995 = (inp[4]) ? node7003 : node6996;
											assign node6996 = (inp[15]) ? node7000 : node6997;
												assign node6997 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7000 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7003 = (inp[0]) ? node7007 : node7004;
												assign node7004 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7007 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7010 = (inp[11]) ? node7026 : node7011;
										assign node7011 = (inp[12]) ? node7019 : node7012;
											assign node7012 = (inp[0]) ? node7016 : node7013;
												assign node7013 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7016 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7019 = (inp[8]) ? node7023 : node7020;
												assign node7020 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node7023 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7026 = (inp[3]) ? node7034 : node7027;
											assign node7027 = (inp[0]) ? node7031 : node7028;
												assign node7028 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7031 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7034 = (inp[9]) ? node7038 : node7035;
												assign node7035 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7038 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7041 = (inp[8]) ? node7105 : node7042;
								assign node7042 = (inp[3]) ? node7074 : node7043;
									assign node7043 = (inp[9]) ? node7059 : node7044;
										assign node7044 = (inp[15]) ? node7052 : node7045;
											assign node7045 = (inp[4]) ? node7049 : node7046;
												assign node7046 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7049 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7052 = (inp[11]) ? node7056 : node7053;
												assign node7053 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7056 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7059 = (inp[0]) ? node7067 : node7060;
											assign node7060 = (inp[7]) ? node7064 : node7061;
												assign node7061 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7064 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7067 = (inp[11]) ? node7071 : node7068;
												assign node7068 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7071 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7074 = (inp[12]) ? node7090 : node7075;
										assign node7075 = (inp[4]) ? node7083 : node7076;
											assign node7076 = (inp[9]) ? node7080 : node7077;
												assign node7077 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7080 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7083 = (inp[11]) ? node7087 : node7084;
												assign node7084 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7087 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7090 = (inp[0]) ? node7098 : node7091;
											assign node7091 = (inp[5]) ? node7095 : node7092;
												assign node7092 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7095 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7098 = (inp[11]) ? node7102 : node7099;
												assign node7099 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7102 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7105 = (inp[0]) ? node7137 : node7106;
									assign node7106 = (inp[9]) ? node7122 : node7107;
										assign node7107 = (inp[15]) ? node7115 : node7108;
											assign node7108 = (inp[12]) ? node7112 : node7109;
												assign node7109 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7112 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7115 = (inp[12]) ? node7119 : node7116;
												assign node7116 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7119 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7122 = (inp[12]) ? node7130 : node7123;
											assign node7123 = (inp[11]) ? node7127 : node7124;
												assign node7124 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7127 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7130 = (inp[7]) ? node7134 : node7131;
												assign node7131 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7134 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7137 = (inp[9]) ? node7153 : node7138;
										assign node7138 = (inp[3]) ? node7146 : node7139;
											assign node7139 = (inp[15]) ? node7143 : node7140;
												assign node7140 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7143 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7146 = (inp[4]) ? node7150 : node7147;
												assign node7147 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7150 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7153 = (inp[12]) ? node7161 : node7154;
											assign node7154 = (inp[15]) ? node7158 : node7155;
												assign node7155 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7158 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7161 = (inp[3]) ? node7165 : node7162;
												assign node7162 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node7165 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node7168 = (inp[15]) ? node7680 : node7169;
					assign node7169 = (inp[11]) ? node7425 : node7170;
						assign node7170 = (inp[5]) ? node7298 : node7171;
							assign node7171 = (inp[7]) ? node7235 : node7172;
								assign node7172 = (inp[0]) ? node7204 : node7173;
									assign node7173 = (inp[10]) ? node7189 : node7174;
										assign node7174 = (inp[8]) ? node7182 : node7175;
											assign node7175 = (inp[4]) ? node7179 : node7176;
												assign node7176 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7179 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7182 = (inp[12]) ? node7186 : node7183;
												assign node7183 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7186 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7189 = (inp[3]) ? node7197 : node7190;
											assign node7190 = (inp[12]) ? node7194 : node7191;
												assign node7191 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7194 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7197 = (inp[8]) ? node7201 : node7198;
												assign node7198 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7201 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7204 = (inp[4]) ? node7220 : node7205;
										assign node7205 = (inp[10]) ? node7213 : node7206;
											assign node7206 = (inp[12]) ? node7210 : node7207;
												assign node7207 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7210 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7213 = (inp[9]) ? node7217 : node7214;
												assign node7214 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7217 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7220 = (inp[3]) ? node7228 : node7221;
											assign node7221 = (inp[10]) ? node7225 : node7222;
												assign node7222 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7225 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7228 = (inp[9]) ? node7232 : node7229;
												assign node7229 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7232 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node7235 = (inp[13]) ? node7267 : node7236;
									assign node7236 = (inp[10]) ? node7252 : node7237;
										assign node7237 = (inp[4]) ? node7245 : node7238;
											assign node7238 = (inp[12]) ? node7242 : node7239;
												assign node7239 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7242 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7245 = (inp[3]) ? node7249 : node7246;
												assign node7246 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7249 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7252 = (inp[9]) ? node7260 : node7253;
											assign node7253 = (inp[3]) ? node7257 : node7254;
												assign node7254 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7257 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7260 = (inp[4]) ? node7264 : node7261;
												assign node7261 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7264 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7267 = (inp[3]) ? node7283 : node7268;
										assign node7268 = (inp[10]) ? node7276 : node7269;
											assign node7269 = (inp[8]) ? node7273 : node7270;
												assign node7270 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7273 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7276 = (inp[4]) ? node7280 : node7277;
												assign node7277 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7280 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7283 = (inp[12]) ? node7291 : node7284;
											assign node7284 = (inp[8]) ? node7288 : node7285;
												assign node7285 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7288 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7291 = (inp[4]) ? node7295 : node7292;
												assign node7292 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7295 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node7298 = (inp[14]) ? node7362 : node7299;
								assign node7299 = (inp[7]) ? node7331 : node7300;
									assign node7300 = (inp[3]) ? node7316 : node7301;
										assign node7301 = (inp[13]) ? node7309 : node7302;
											assign node7302 = (inp[10]) ? node7306 : node7303;
												assign node7303 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7306 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7309 = (inp[4]) ? node7313 : node7310;
												assign node7310 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7313 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7316 = (inp[12]) ? node7324 : node7317;
											assign node7317 = (inp[0]) ? node7321 : node7318;
												assign node7318 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7321 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7324 = (inp[0]) ? node7328 : node7325;
												assign node7325 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7328 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7331 = (inp[0]) ? node7347 : node7332;
										assign node7332 = (inp[8]) ? node7340 : node7333;
											assign node7333 = (inp[4]) ? node7337 : node7334;
												assign node7334 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7337 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7340 = (inp[13]) ? node7344 : node7341;
												assign node7341 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7344 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7347 = (inp[13]) ? node7355 : node7348;
											assign node7348 = (inp[3]) ? node7352 : node7349;
												assign node7349 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7352 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7355 = (inp[4]) ? node7359 : node7356;
												assign node7356 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7359 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7362 = (inp[10]) ? node7394 : node7363;
									assign node7363 = (inp[0]) ? node7379 : node7364;
										assign node7364 = (inp[3]) ? node7372 : node7365;
											assign node7365 = (inp[7]) ? node7369 : node7366;
												assign node7366 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7369 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7372 = (inp[13]) ? node7376 : node7373;
												assign node7373 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7376 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7379 = (inp[8]) ? node7387 : node7380;
											assign node7380 = (inp[9]) ? node7384 : node7381;
												assign node7381 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7384 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7387 = (inp[9]) ? node7391 : node7388;
												assign node7388 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7391 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7394 = (inp[7]) ? node7410 : node7395;
										assign node7395 = (inp[13]) ? node7403 : node7396;
											assign node7396 = (inp[12]) ? node7400 : node7397;
												assign node7397 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7400 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7403 = (inp[8]) ? node7407 : node7404;
												assign node7404 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7407 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7410 = (inp[4]) ? node7418 : node7411;
											assign node7411 = (inp[13]) ? node7415 : node7412;
												assign node7412 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7415 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7418 = (inp[3]) ? node7422 : node7419;
												assign node7419 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7422 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node7425 = (inp[0]) ? node7553 : node7426;
							assign node7426 = (inp[7]) ? node7490 : node7427;
								assign node7427 = (inp[14]) ? node7459 : node7428;
									assign node7428 = (inp[12]) ? node7444 : node7429;
										assign node7429 = (inp[4]) ? node7437 : node7430;
											assign node7430 = (inp[5]) ? node7434 : node7431;
												assign node7431 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7434 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7437 = (inp[3]) ? node7441 : node7438;
												assign node7438 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7441 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7444 = (inp[9]) ? node7452 : node7445;
											assign node7445 = (inp[3]) ? node7449 : node7446;
												assign node7446 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7449 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7452 = (inp[5]) ? node7456 : node7453;
												assign node7453 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7456 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7459 = (inp[8]) ? node7475 : node7460;
										assign node7460 = (inp[3]) ? node7468 : node7461;
											assign node7461 = (inp[13]) ? node7465 : node7462;
												assign node7462 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node7465 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7468 = (inp[5]) ? node7472 : node7469;
												assign node7469 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7472 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7475 = (inp[10]) ? node7483 : node7476;
											assign node7476 = (inp[4]) ? node7480 : node7477;
												assign node7477 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7480 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7483 = (inp[4]) ? node7487 : node7484;
												assign node7484 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7487 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7490 = (inp[4]) ? node7522 : node7491;
									assign node7491 = (inp[9]) ? node7507 : node7492;
										assign node7492 = (inp[5]) ? node7500 : node7493;
											assign node7493 = (inp[12]) ? node7497 : node7494;
												assign node7494 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7497 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7500 = (inp[3]) ? node7504 : node7501;
												assign node7501 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7504 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7507 = (inp[13]) ? node7515 : node7508;
											assign node7508 = (inp[3]) ? node7512 : node7509;
												assign node7509 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7512 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7515 = (inp[3]) ? node7519 : node7516;
												assign node7516 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7519 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7522 = (inp[14]) ? node7538 : node7523;
										assign node7523 = (inp[12]) ? node7531 : node7524;
											assign node7524 = (inp[13]) ? node7528 : node7525;
												assign node7525 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7528 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7531 = (inp[5]) ? node7535 : node7532;
												assign node7532 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7535 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7538 = (inp[5]) ? node7546 : node7539;
											assign node7539 = (inp[13]) ? node7543 : node7540;
												assign node7540 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7543 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7546 = (inp[12]) ? node7550 : node7547;
												assign node7547 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7550 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7553 = (inp[8]) ? node7617 : node7554;
								assign node7554 = (inp[9]) ? node7586 : node7555;
									assign node7555 = (inp[13]) ? node7571 : node7556;
										assign node7556 = (inp[12]) ? node7564 : node7557;
											assign node7557 = (inp[14]) ? node7561 : node7558;
												assign node7558 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7561 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7564 = (inp[3]) ? node7568 : node7565;
												assign node7565 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7568 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7571 = (inp[4]) ? node7579 : node7572;
											assign node7572 = (inp[3]) ? node7576 : node7573;
												assign node7573 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7576 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7579 = (inp[5]) ? node7583 : node7580;
												assign node7580 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7583 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7586 = (inp[10]) ? node7602 : node7587;
										assign node7587 = (inp[3]) ? node7595 : node7588;
											assign node7588 = (inp[5]) ? node7592 : node7589;
												assign node7589 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7592 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7595 = (inp[14]) ? node7599 : node7596;
												assign node7596 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7599 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7602 = (inp[7]) ? node7610 : node7603;
											assign node7603 = (inp[4]) ? node7607 : node7604;
												assign node7604 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7607 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7610 = (inp[12]) ? node7614 : node7611;
												assign node7611 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7614 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7617 = (inp[5]) ? node7649 : node7618;
									assign node7618 = (inp[13]) ? node7634 : node7619;
										assign node7619 = (inp[12]) ? node7627 : node7620;
											assign node7620 = (inp[14]) ? node7624 : node7621;
												assign node7621 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7624 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7627 = (inp[14]) ? node7631 : node7628;
												assign node7628 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7631 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7634 = (inp[4]) ? node7642 : node7635;
											assign node7635 = (inp[7]) ? node7639 : node7636;
												assign node7636 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7639 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7642 = (inp[9]) ? node7646 : node7643;
												assign node7643 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7646 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7649 = (inp[3]) ? node7665 : node7650;
										assign node7650 = (inp[7]) ? node7658 : node7651;
											assign node7651 = (inp[4]) ? node7655 : node7652;
												assign node7652 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7655 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7658 = (inp[4]) ? node7662 : node7659;
												assign node7659 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7662 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7665 = (inp[13]) ? node7673 : node7666;
											assign node7666 = (inp[4]) ? node7670 : node7667;
												assign node7667 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7670 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7673 = (inp[10]) ? node7677 : node7674;
												assign node7674 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node7677 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node7680 = (inp[8]) ? node7936 : node7681;
						assign node7681 = (inp[10]) ? node7809 : node7682;
							assign node7682 = (inp[5]) ? node7746 : node7683;
								assign node7683 = (inp[12]) ? node7715 : node7684;
									assign node7684 = (inp[0]) ? node7700 : node7685;
										assign node7685 = (inp[9]) ? node7693 : node7686;
											assign node7686 = (inp[3]) ? node7690 : node7687;
												assign node7687 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7690 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7693 = (inp[11]) ? node7697 : node7694;
												assign node7694 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7697 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7700 = (inp[3]) ? node7708 : node7701;
											assign node7701 = (inp[14]) ? node7705 : node7702;
												assign node7702 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7705 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7708 = (inp[9]) ? node7712 : node7709;
												assign node7709 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7712 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7715 = (inp[3]) ? node7731 : node7716;
										assign node7716 = (inp[4]) ? node7724 : node7717;
											assign node7717 = (inp[7]) ? node7721 : node7718;
												assign node7718 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7721 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7724 = (inp[0]) ? node7728 : node7725;
												assign node7725 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7728 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7731 = (inp[11]) ? node7739 : node7732;
											assign node7732 = (inp[14]) ? node7736 : node7733;
												assign node7733 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7736 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7739 = (inp[0]) ? node7743 : node7740;
												assign node7740 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7743 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7746 = (inp[11]) ? node7778 : node7747;
									assign node7747 = (inp[3]) ? node7763 : node7748;
										assign node7748 = (inp[9]) ? node7756 : node7749;
											assign node7749 = (inp[14]) ? node7753 : node7750;
												assign node7750 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7753 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7756 = (inp[12]) ? node7760 : node7757;
												assign node7757 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7760 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7763 = (inp[7]) ? node7771 : node7764;
											assign node7764 = (inp[13]) ? node7768 : node7765;
												assign node7765 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7768 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7771 = (inp[14]) ? node7775 : node7772;
												assign node7772 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7775 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7778 = (inp[9]) ? node7794 : node7779;
										assign node7779 = (inp[14]) ? node7787 : node7780;
											assign node7780 = (inp[3]) ? node7784 : node7781;
												assign node7781 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7784 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7787 = (inp[7]) ? node7791 : node7788;
												assign node7788 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7791 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7794 = (inp[4]) ? node7802 : node7795;
											assign node7795 = (inp[7]) ? node7799 : node7796;
												assign node7796 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7799 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7802 = (inp[12]) ? node7806 : node7803;
												assign node7803 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7806 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7809 = (inp[12]) ? node7873 : node7810;
								assign node7810 = (inp[11]) ? node7842 : node7811;
									assign node7811 = (inp[14]) ? node7827 : node7812;
										assign node7812 = (inp[0]) ? node7820 : node7813;
											assign node7813 = (inp[7]) ? node7817 : node7814;
												assign node7814 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7817 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7820 = (inp[3]) ? node7824 : node7821;
												assign node7821 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7824 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7827 = (inp[0]) ? node7835 : node7828;
											assign node7828 = (inp[3]) ? node7832 : node7829;
												assign node7829 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7832 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7835 = (inp[4]) ? node7839 : node7836;
												assign node7836 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7839 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7842 = (inp[5]) ? node7858 : node7843;
										assign node7843 = (inp[9]) ? node7851 : node7844;
											assign node7844 = (inp[0]) ? node7848 : node7845;
												assign node7845 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7848 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7851 = (inp[4]) ? node7855 : node7852;
												assign node7852 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7855 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7858 = (inp[9]) ? node7866 : node7859;
											assign node7859 = (inp[13]) ? node7863 : node7860;
												assign node7860 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7863 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7866 = (inp[4]) ? node7870 : node7867;
												assign node7867 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7870 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7873 = (inp[5]) ? node7905 : node7874;
									assign node7874 = (inp[7]) ? node7890 : node7875;
										assign node7875 = (inp[0]) ? node7883 : node7876;
											assign node7876 = (inp[13]) ? node7880 : node7877;
												assign node7877 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7880 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7883 = (inp[9]) ? node7887 : node7884;
												assign node7884 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7887 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7890 = (inp[11]) ? node7898 : node7891;
											assign node7891 = (inp[13]) ? node7895 : node7892;
												assign node7892 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node7895 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7898 = (inp[9]) ? node7902 : node7899;
												assign node7899 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7902 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7905 = (inp[4]) ? node7921 : node7906;
										assign node7906 = (inp[3]) ? node7914 : node7907;
											assign node7907 = (inp[14]) ? node7911 : node7908;
												assign node7908 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7911 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7914 = (inp[9]) ? node7918 : node7915;
												assign node7915 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7918 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7921 = (inp[11]) ? node7929 : node7922;
											assign node7922 = (inp[3]) ? node7926 : node7923;
												assign node7923 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7926 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7929 = (inp[13]) ? node7933 : node7930;
												assign node7930 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node7933 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node7936 = (inp[14]) ? node8064 : node7937;
							assign node7937 = (inp[13]) ? node8001 : node7938;
								assign node7938 = (inp[4]) ? node7970 : node7939;
									assign node7939 = (inp[0]) ? node7955 : node7940;
										assign node7940 = (inp[9]) ? node7948 : node7941;
											assign node7941 = (inp[7]) ? node7945 : node7942;
												assign node7942 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7945 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7948 = (inp[5]) ? node7952 : node7949;
												assign node7949 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7952 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7955 = (inp[7]) ? node7963 : node7956;
											assign node7956 = (inp[3]) ? node7960 : node7957;
												assign node7957 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7960 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7963 = (inp[9]) ? node7967 : node7964;
												assign node7964 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7967 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7970 = (inp[11]) ? node7986 : node7971;
										assign node7971 = (inp[3]) ? node7979 : node7972;
											assign node7972 = (inp[0]) ? node7976 : node7973;
												assign node7973 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7976 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7979 = (inp[0]) ? node7983 : node7980;
												assign node7980 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7983 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7986 = (inp[5]) ? node7994 : node7987;
											assign node7987 = (inp[9]) ? node7991 : node7988;
												assign node7988 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7991 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7994 = (inp[3]) ? node7998 : node7995;
												assign node7995 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7998 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node8001 = (inp[9]) ? node8033 : node8002;
									assign node8002 = (inp[0]) ? node8018 : node8003;
										assign node8003 = (inp[12]) ? node8011 : node8004;
											assign node8004 = (inp[11]) ? node8008 : node8005;
												assign node8005 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8008 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8011 = (inp[3]) ? node8015 : node8012;
												assign node8012 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8015 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8018 = (inp[5]) ? node8026 : node8019;
											assign node8019 = (inp[11]) ? node8023 : node8020;
												assign node8020 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8023 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8026 = (inp[7]) ? node8030 : node8027;
												assign node8027 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8030 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node8033 = (inp[4]) ? node8049 : node8034;
										assign node8034 = (inp[11]) ? node8042 : node8035;
											assign node8035 = (inp[12]) ? node8039 : node8036;
												assign node8036 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8039 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8042 = (inp[5]) ? node8046 : node8043;
												assign node8043 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8046 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node8049 = (inp[3]) ? node8057 : node8050;
											assign node8050 = (inp[0]) ? node8054 : node8051;
												assign node8051 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8054 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8057 = (inp[11]) ? node8061 : node8058;
												assign node8058 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8061 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node8064 = (inp[7]) ? node8128 : node8065;
								assign node8065 = (inp[13]) ? node8097 : node8066;
									assign node8066 = (inp[12]) ? node8082 : node8067;
										assign node8067 = (inp[4]) ? node8075 : node8068;
											assign node8068 = (inp[9]) ? node8072 : node8069;
												assign node8069 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8072 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8075 = (inp[5]) ? node8079 : node8076;
												assign node8076 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8079 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8082 = (inp[9]) ? node8090 : node8083;
											assign node8083 = (inp[4]) ? node8087 : node8084;
												assign node8084 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8087 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8090 = (inp[11]) ? node8094 : node8091;
												assign node8091 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8094 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node8097 = (inp[11]) ? node8113 : node8098;
										assign node8098 = (inp[3]) ? node8106 : node8099;
											assign node8099 = (inp[12]) ? node8103 : node8100;
												assign node8100 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8103 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8106 = (inp[4]) ? node8110 : node8107;
												assign node8107 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8110 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node8113 = (inp[0]) ? node8121 : node8114;
											assign node8114 = (inp[5]) ? node8118 : node8115;
												assign node8115 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8118 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8121 = (inp[12]) ? node8125 : node8122;
												assign node8122 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8125 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node8128 = (inp[3]) ? node8160 : node8129;
									assign node8129 = (inp[0]) ? node8145 : node8130;
										assign node8130 = (inp[5]) ? node8138 : node8131;
											assign node8131 = (inp[12]) ? node8135 : node8132;
												assign node8132 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8135 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8138 = (inp[11]) ? node8142 : node8139;
												assign node8139 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8142 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node8145 = (inp[9]) ? node8153 : node8146;
											assign node8146 = (inp[11]) ? node8150 : node8147;
												assign node8147 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8150 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8153 = (inp[4]) ? node8157 : node8154;
												assign node8154 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8157 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node8160 = (inp[11]) ? node8176 : node8161;
										assign node8161 = (inp[5]) ? node8169 : node8162;
											assign node8162 = (inp[13]) ? node8166 : node8163;
												assign node8163 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8166 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8169 = (inp[9]) ? node8173 : node8170;
												assign node8170 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8173 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node8176 = (inp[12]) ? node8184 : node8177;
											assign node8177 = (inp[10]) ? node8181 : node8178;
												assign node8178 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8181 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node8184 = (inp[0]) ? node8188 : node8185;
												assign node8185 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node8188 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;

endmodule