module dtc_split125_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node3;
	wire [40-1:0] node5;
	wire [40-1:0] node7;
	wire [40-1:0] node8;
	wire [40-1:0] node10;
	wire [40-1:0] node15;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node41;
	wire [40-1:0] node44;
	wire [40-1:0] node46;
	wire [40-1:0] node48;
	wire [40-1:0] node50;
	wire [40-1:0] node51;
	wire [40-1:0] node53;
	wire [40-1:0] node56;
	wire [40-1:0] node57;
	wire [40-1:0] node60;
	wire [40-1:0] node63;
	wire [40-1:0] node64;
	wire [40-1:0] node66;
	wire [40-1:0] node67;
	wire [40-1:0] node68;
	wire [40-1:0] node70;
	wire [40-1:0] node72;
	wire [40-1:0] node76;
	wire [40-1:0] node77;
	wire [40-1:0] node78;
	wire [40-1:0] node80;
	wire [40-1:0] node83;
	wire [40-1:0] node85;
	wire [40-1:0] node89;
	wire [40-1:0] node90;
	wire [40-1:0] node91;
	wire [40-1:0] node94;
	wire [40-1:0] node97;
	wire [40-1:0] node99;
	wire [40-1:0] node100;
	wire [40-1:0] node102;
	wire [40-1:0] node104;
	wire [40-1:0] node107;
	wire [40-1:0] node108;
	wire [40-1:0] node109;
	wire [40-1:0] node110;
	wire [40-1:0] node113;
	wire [40-1:0] node116;
	wire [40-1:0] node118;
	wire [40-1:0] node121;
	wire [40-1:0] node122;
	wire [40-1:0] node123;
	wire [40-1:0] node127;
	wire [40-1:0] node130;
	wire [40-1:0] node131;
	wire [40-1:0] node132;
	wire [40-1:0] node135;
	wire [40-1:0] node136;
	wire [40-1:0] node137;
	wire [40-1:0] node138;
	wire [40-1:0] node139;
	wire [40-1:0] node142;
	wire [40-1:0] node145;
	wire [40-1:0] node146;
	wire [40-1:0] node149;
	wire [40-1:0] node152;
	wire [40-1:0] node153;
	wire [40-1:0] node154;
	wire [40-1:0] node157;
	wire [40-1:0] node160;
	wire [40-1:0] node161;
	wire [40-1:0] node164;
	wire [40-1:0] node167;
	wire [40-1:0] node168;
	wire [40-1:0] node169;
	wire [40-1:0] node170;
	wire [40-1:0] node173;
	wire [40-1:0] node176;
	wire [40-1:0] node177;
	wire [40-1:0] node180;
	wire [40-1:0] node183;
	wire [40-1:0] node184;
	wire [40-1:0] node185;
	wire [40-1:0] node188;
	wire [40-1:0] node191;
	wire [40-1:0] node192;
	wire [40-1:0] node195;
	wire [40-1:0] node198;
	wire [40-1:0] node199;
	wire [40-1:0] node202;
	wire [40-1:0] node204;
	wire [40-1:0] node205;
	wire [40-1:0] node206;
	wire [40-1:0] node207;
	wire [40-1:0] node208;
	wire [40-1:0] node209;
	wire [40-1:0] node210;
	wire [40-1:0] node212;
	wire [40-1:0] node215;
	wire [40-1:0] node216;
	wire [40-1:0] node219;
	wire [40-1:0] node222;
	wire [40-1:0] node223;
	wire [40-1:0] node224;
	wire [40-1:0] node227;
	wire [40-1:0] node230;
	wire [40-1:0] node231;
	wire [40-1:0] node234;
	wire [40-1:0] node237;
	wire [40-1:0] node238;
	wire [40-1:0] node239;
	wire [40-1:0] node240;
	wire [40-1:0] node243;
	wire [40-1:0] node246;
	wire [40-1:0] node247;
	wire [40-1:0] node250;
	wire [40-1:0] node253;
	wire [40-1:0] node254;
	wire [40-1:0] node255;
	wire [40-1:0] node258;
	wire [40-1:0] node261;
	wire [40-1:0] node262;
	wire [40-1:0] node265;
	wire [40-1:0] node268;
	wire [40-1:0] node269;
	wire [40-1:0] node271;
	wire [40-1:0] node273;
	wire [40-1:0] node275;
	wire [40-1:0] node278;
	wire [40-1:0] node279;
	wire [40-1:0] node280;
	wire [40-1:0] node282;
	wire [40-1:0] node285;
	wire [40-1:0] node286;
	wire [40-1:0] node289;
	wire [40-1:0] node292;
	wire [40-1:0] node293;
	wire [40-1:0] node294;
	wire [40-1:0] node297;
	wire [40-1:0] node300;
	wire [40-1:0] node301;
	wire [40-1:0] node304;
	wire [40-1:0] node307;
	wire [40-1:0] node308;
	wire [40-1:0] node309;
	wire [40-1:0] node310;
	wire [40-1:0] node311;
	wire [40-1:0] node312;
	wire [40-1:0] node315;
	wire [40-1:0] node318;
	wire [40-1:0] node320;
	wire [40-1:0] node323;
	wire [40-1:0] node324;
	wire [40-1:0] node325;
	wire [40-1:0] node331;
	wire [40-1:0] node333;
	wire [40-1:0] node334;
	wire [40-1:0] node335;
	wire [40-1:0] node336;
	wire [40-1:0] node339;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node346;
	wire [40-1:0] node349;
	wire [40-1:0] node350;
	wire [40-1:0] node351;
	wire [40-1:0] node354;
	wire [40-1:0] node357;
	wire [40-1:0] node358;
	wire [40-1:0] node361;
	wire [40-1:0] node364;
	wire [40-1:0] node365;
	wire [40-1:0] node366;
	wire [40-1:0] node368;
	wire [40-1:0] node370;
	wire [40-1:0] node371;
	wire [40-1:0] node373;
	wire [40-1:0] node376;
	wire [40-1:0] node377;
	wire [40-1:0] node380;
	wire [40-1:0] node383;
	wire [40-1:0] node384;
	wire [40-1:0] node385;
	wire [40-1:0] node386;
	wire [40-1:0] node388;
	wire [40-1:0] node391;
	wire [40-1:0] node392;
	wire [40-1:0] node396;
	wire [40-1:0] node397;
	wire [40-1:0] node399;
	wire [40-1:0] node402;
	wire [40-1:0] node403;
	wire [40-1:0] node408;
	wire [40-1:0] node409;
	wire [40-1:0] node411;
	wire [40-1:0] node412;
	wire [40-1:0] node413;
	wire [40-1:0] node415;
	wire [40-1:0] node418;
	wire [40-1:0] node419;
	wire [40-1:0] node422;
	wire [40-1:0] node425;
	wire [40-1:0] node426;
	wire [40-1:0] node427;
	wire [40-1:0] node430;
	wire [40-1:0] node433;
	wire [40-1:0] node434;
	wire [40-1:0] node437;
	wire [40-1:0] node440;
	wire [40-1:0] node441;
	wire [40-1:0] node442;
	wire [40-1:0] node443;
	wire [40-1:0] node444;
	wire [40-1:0] node447;
	wire [40-1:0] node450;
	wire [40-1:0] node451;
	wire [40-1:0] node454;
	wire [40-1:0] node457;
	wire [40-1:0] node458;
	wire [40-1:0] node459;
	wire [40-1:0] node462;
	wire [40-1:0] node465;
	wire [40-1:0] node467;

	assign outp = (inp[9]) ? node130 : node1;
		assign node1 = (inp[1]) ? node15 : node2;
			assign node2 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node3;
				assign node3 = (inp[4]) ? node5 : 40'b0000000000000000000000000000000000000000;
					assign node5 = (inp[8]) ? node7 : 40'b0000000000000000000000000000000000000000;
						assign node7 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node8;
							assign node8 = (inp[7]) ? node10 : 40'b0000000000000000000000000000000000000000;
								assign node10 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
			assign node15 = (inp[4]) ? node17 : 40'b0000000001000000000000000000000000000000;
				assign node17 = (inp[8]) ? node63 : node18;
					assign node18 = (inp[7]) ? node44 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[11]) ? node24 : node21;
								assign node21 = (inp[3]) ? 40'b0000000000100010000000000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[3]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000000010000001000000000000000000;
							assign node27 = (inp[11]) ? node31 : node28;
								assign node28 = (inp[3]) ? 40'b0000000000100000000000000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[3]) ? node33 : 40'b0000000000000000000001000000000010000000;
									assign node33 = (inp[10]) ? node39 : node34;
										assign node34 = (inp[0]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[13]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[0]) ? node41 : 40'b0000000000000010010000010000000010000000;
											assign node41 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000010000010000000010000000;
						assign node44 = (inp[3]) ? node46 : 40'b0000000000000000000000000000000000000000;
							assign node46 = (inp[11]) ? node48 : 40'b0000000000000000000000000000000000000000;
								assign node48 = (inp[14]) ? node50 : 40'b0000000000000000000000000000000000000000;
									assign node50 = (inp[10]) ? node56 : node51;
										assign node51 = (inp[13]) ? node53 : 40'b0000000000000000000000000000000000000000;
											assign node53 = (inp[0]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node56 = (inp[13]) ? node60 : node57;
											assign node57 = (inp[0]) ? 40'b0000000000000000000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node60 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000110000000;
					assign node63 = (inp[14]) ? node89 : node64;
						assign node64 = (inp[0]) ? node66 : 40'b0000000000000000000000000000000000000000;
							assign node66 = (inp[13]) ? node76 : node67;
								assign node67 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node68;
									assign node68 = (inp[12]) ? node70 : 40'b0000000000000000000000000000000000000000;
										assign node70 = (inp[3]) ? node72 : 40'b0000000000000000000000000000000000000000;
											assign node72 = (inp[11]) ? 40'b0000000010000001010000000000010000000000 : 40'b0000000010000001010000000000000000000000;
								assign node76 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node77;
									assign node77 = (inp[7]) ? node83 : node78;
										assign node78 = (inp[10]) ? node80 : 40'b0000000000000000000000000000000000000000;
											assign node80 = (inp[3]) ? 40'b0000000000000000000000000000001000000000 : 40'b0000000000000000000000000000000000000000;
										assign node83 = (inp[3]) ? node85 : 40'b0000000000000000000000000000000000000000;
											assign node85 = (inp[10]) ? 40'b0000000000000000000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
						assign node89 = (inp[3]) ? node97 : node90;
							assign node90 = (inp[7]) ? node94 : node91;
								assign node91 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node94 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
							assign node97 = (inp[0]) ? node99 : 40'b0000000000000000000000000000000000000000;
								assign node99 = (inp[15]) ? node107 : node100;
									assign node100 = (inp[13]) ? node102 : 40'b0000000000000000000000000000000000000000;
										assign node102 = (inp[10]) ? node104 : 40'b0000000000000000000000000000000000000000;
											assign node104 = (inp[6]) ? 40'b0000000010001000000000000000000001000010 : 40'b0100000000000000000000011000000100000000;
									assign node107 = (inp[7]) ? node121 : node108;
										assign node108 = (inp[11]) ? node116 : node109;
											assign node109 = (inp[6]) ? node113 : node110;
												assign node110 = (inp[5]) ? 40'b0000000000000000000100000000001001000010 : 40'b0000000000000000000000000000000000000000;
												assign node113 = (inp[5]) ? 40'b0000000010000000010100100000000001000000 : 40'b0000000000000000000100000000000001000010;
											assign node116 = (inp[13]) ? node118 : 40'b0000000000000000000000000000000000000000;
												assign node118 = (inp[10]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000010001010010000100000000001000000;
										assign node121 = (inp[13]) ? node127 : node122;
											assign node122 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node123;
												assign node123 = (inp[2]) ? 40'b0100000000000001000000001000001100000000 : 40'b0000000000000000000000000000000000000000;
											assign node127 = (inp[11]) ? 40'b0100000000000010000000100000000100000011 : 40'b0100000000000000000000011000000100000000;
		assign node130 = (inp[1]) ? node198 : node131;
			assign node131 = (inp[8]) ? node135 : node132;
				assign node132 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node135 = (inp[7]) ? node167 : node136;
					assign node136 = (inp[3]) ? node152 : node137;
						assign node137 = (inp[11]) ? node145 : node138;
							assign node138 = (inp[14]) ? node142 : node139;
								assign node139 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node142 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
							assign node145 = (inp[14]) ? node149 : node146;
								assign node146 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node149 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
						assign node152 = (inp[14]) ? node160 : node153;
							assign node153 = (inp[11]) ? node157 : node154;
								assign node154 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node157 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
							assign node160 = (inp[11]) ? node164 : node161;
								assign node161 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
								assign node164 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node167 = (inp[11]) ? node183 : node168;
						assign node168 = (inp[14]) ? node176 : node169;
							assign node169 = (inp[3]) ? node173 : node170;
								assign node170 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node173 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
							assign node176 = (inp[3]) ? node180 : node177;
								assign node177 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node180 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
						assign node183 = (inp[3]) ? node191 : node184;
							assign node184 = (inp[14]) ? node188 : node185;
								assign node185 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
								assign node188 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
							assign node191 = (inp[14]) ? node195 : node192;
								assign node192 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
								assign node195 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node198 = (inp[4]) ? node202 : node199;
				assign node199 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node202 = (inp[8]) ? node204 : 40'b0000100000000000000000000000000000000000;
					assign node204 = (inp[7]) ? node364 : node205;
						assign node205 = (inp[3]) ? node307 : node206;
							assign node206 = (inp[14]) ? node268 : node207;
								assign node207 = (inp[11]) ? node237 : node208;
									assign node208 = (inp[10]) ? node222 : node209;
										assign node209 = (inp[13]) ? node215 : node210;
											assign node210 = (inp[0]) ? node212 : 40'b1001000000010101010110000010101000010000;
												assign node212 = (inp[12]) ? 40'b0000000000011101010110000010101000010000 : 40'b0000000000001101010110000010101000010000;
											assign node215 = (inp[15]) ? node219 : node216;
												assign node216 = (inp[5]) ? 40'b0001000000011101010010000011001000010000 : 40'b1000000000011101010010000010001000010000;
												assign node219 = (inp[6]) ? 40'b0000000000001101010010000011001000010000 : 40'b1001000000000101010010000001001000010000;
										assign node222 = (inp[6]) ? node230 : node223;
											assign node223 = (inp[15]) ? node227 : node224;
												assign node224 = (inp[12]) ? 40'b1000000000010001010010000001001000010000 : 40'b1000000000010001010110000010001000010000;
												assign node227 = (inp[0]) ? 40'b1000000000000001010010000010101000010000 : 40'b0001000000000001010110000010101000010000;
											assign node230 = (inp[12]) ? node234 : node231;
												assign node231 = (inp[5]) ? 40'b1001000000010001010010000001001000010000 : 40'b0000000000001001010110000010001000010000;
												assign node234 = (inp[13]) ? 40'b0001000000011001010010000011001000010000 : 40'b0001000000011001010010000011101000010000;
									assign node237 = (inp[15]) ? node253 : node238;
										assign node238 = (inp[13]) ? node246 : node239;
											assign node239 = (inp[12]) ? node243 : node240;
												assign node240 = (inp[6]) ? 40'b1000000000011001010010000010101000000000 : 40'b0000000000010001010110000010101000000000;
												assign node243 = (inp[2]) ? 40'b0000000000010001010010000001101000000000 : 40'b0000000000011001010010000011101000000000;
											assign node246 = (inp[10]) ? node250 : node247;
												assign node247 = (inp[2]) ? 40'b0000000000010101010110000010001000000000 : 40'b1000000000010101010010000000001000000000;
												assign node250 = (inp[12]) ? 40'b0001000000011001010010000010001000000000 : 40'b0000000000010001010110000010001000000000;
										assign node253 = (inp[13]) ? node261 : node254;
											assign node254 = (inp[0]) ? node258 : node255;
												assign node255 = (inp[6]) ? 40'b1001000000001001010010000010101000000000 : 40'b1001000000000001010110000010101000000000;
												assign node258 = (inp[10]) ? 40'b0000000000001001010010000010101000000000 : 40'b0000000000000101010110000010101000000000;
											assign node261 = (inp[5]) ? node265 : node262;
												assign node262 = (inp[10]) ? 40'b1001000000000001010010000000001000000000 : 40'b1001000000001101010010000010001000000000;
												assign node265 = (inp[2]) ? 40'b0001000000000001010110000011001000000000 : 40'b1001000000000101010110000010001000000000;
								assign node268 = (inp[11]) ? node278 : node269;
									assign node269 = (inp[15]) ? node271 : 40'b0000000000000000000000000000000000000000;
										assign node271 = (inp[0]) ? node273 : 40'b0000000000000000000000000000000000000000;
											assign node273 = (inp[2]) ? node275 : 40'b0000000000000000000000000000000000000000;
												assign node275 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000100001100000010000000000000;
									assign node278 = (inp[13]) ? node292 : node279;
										assign node279 = (inp[2]) ? node285 : node280;
											assign node280 = (inp[0]) ? node282 : 40'b1001010000000100000000000001100000000000;
												assign node282 = (inp[15]) ? 40'b1000010000000000000000000001100000000000 : 40'b1000010000010000000000000001100000000000;
											assign node285 = (inp[5]) ? node289 : node286;
												assign node286 = (inp[15]) ? 40'b0000010000001000000000000011100000000000 : 40'b1001010000010000000000000001100000000000;
												assign node289 = (inp[10]) ? 40'b0000010000000000000100000010100000000000 : 40'b0000010000000100000100000011100000000000;
										assign node292 = (inp[0]) ? node300 : node293;
											assign node293 = (inp[10]) ? node297 : node294;
												assign node294 = (inp[5]) ? 40'b1001010000000100000100000010000000000000 : 40'b1001010000000100000000000001000000000000;
												assign node297 = (inp[2]) ? 40'b0001010000000000000000000001000000000000 : 40'b0001010000001000000000000010000000000000;
											assign node300 = (inp[10]) ? node304 : node301;
												assign node301 = (inp[15]) ? 40'b0000010000001100000100000010000000000000 : 40'b1000010000011100000000000010000000000000;
												assign node304 = (inp[5]) ? 40'b0000010000011000000000000011000000000000 : 40'b0000010000001000000000000010000000000000;
							assign node307 = (inp[14]) ? node331 : node308;
								assign node308 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node309;
									assign node309 = (inp[6]) ? node323 : node310;
										assign node310 = (inp[15]) ? node318 : node311;
											assign node311 = (inp[2]) ? node315 : node312;
												assign node312 = (inp[0]) ? 40'b1000000000010000000000000000000000100000 : 40'b1001000000010000000000000000000000100000;
												assign node315 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node318 = (inp[0]) ? node320 : 40'b0000000000000000000000000000000000000000;
												assign node320 = (inp[2]) ? 40'b0000000000000100000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
										assign node323 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node324;
											assign node324 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node325;
												assign node325 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
								assign node331 = (inp[11]) ? node333 : 40'b0000000000000000000000000000000000000000;
									assign node333 = (inp[10]) ? node349 : node334;
										assign node334 = (inp[13]) ? node342 : node335;
											assign node335 = (inp[0]) ? node339 : node336;
												assign node336 = (inp[5]) ? 40'b0011000000010100000100000010100000000000 : 40'b1011000000000100000000000001100000000000;
												assign node339 = (inp[15]) ? 40'b0010000000001100000000000010100000000000 : 40'b0010000000011100000000000010100000000000;
											assign node342 = (inp[15]) ? node346 : node343;
												assign node343 = (inp[2]) ? 40'b0011000000010100000000000001000000000000 : 40'b1010000000010100000000000000000000000000;
												assign node346 = (inp[0]) ? 40'b1010000000000100000100000011000000000000 : 40'b1011000000000100000000000001000000000000;
										assign node349 = (inp[0]) ? node357 : node350;
											assign node350 = (inp[5]) ? node354 : node351;
												assign node351 = (inp[2]) ? 40'b0011000000001000000100000010000000000000 : 40'b1011000000001000000000000010100000000000;
												assign node354 = (inp[12]) ? 40'b0011000000010000000100000011100000000000 : 40'b1011000000010000000100000010000000000000;
											assign node357 = (inp[13]) ? node361 : node358;
												assign node358 = (inp[2]) ? 40'b0010000000010000000000000001100000000000 : 40'b0010000000001000000000000010100000000000;
												assign node361 = (inp[15]) ? 40'b1010000000000000000000000001000000000000 : 40'b0010000000011000000100000011000000000000;
						assign node364 = (inp[3]) ? node408 : node365;
							assign node365 = (inp[11]) ? node383 : node366;
								assign node366 = (inp[14]) ? node368 : 40'b0000000000000000000000000000000000000000;
									assign node368 = (inp[0]) ? node370 : 40'b0000000000000000000000000000000000000000;
										assign node370 = (inp[15]) ? node376 : node371;
											assign node371 = (inp[13]) ? node373 : 40'b0000000000000000000000000000000000000000;
												assign node373 = (inp[10]) ? 40'b0000001100010000000100000011000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node376 = (inp[2]) ? node380 : node377;
												assign node377 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000001100001000000000000010000000000000;
												assign node380 = (inp[5]) ? 40'b0000001100000000000100000011100000000000 : 40'b0000001100001000000000000011100000000000;
								assign node383 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node384;
									assign node384 = (inp[15]) ? node396 : node385;
										assign node385 = (inp[0]) ? node391 : node386;
											assign node386 = (inp[10]) ? node388 : 40'b0000000000000000000000000000000000000000;
												assign node388 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
											assign node391 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node392;
												assign node392 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
										assign node396 = (inp[10]) ? node402 : node397;
											assign node397 = (inp[0]) ? node399 : 40'b0000000000000000000000000000000000000000;
												assign node399 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
											assign node402 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node403;
												assign node403 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
							assign node408 = (inp[14]) ? node440 : node409;
								assign node409 = (inp[11]) ? node411 : 40'b0000000000000000000000000000000000000000;
									assign node411 = (inp[10]) ? node425 : node412;
										assign node412 = (inp[5]) ? node418 : node413;
											assign node413 = (inp[0]) ? node415 : 40'b0001001000001100000100000010000000001000;
												assign node415 = (inp[12]) ? 40'b1000001000011100000000000010000000001000 : 40'b1000001000001100000000000010100000001000;
											assign node418 = (inp[12]) ? node422 : node419;
												assign node419 = (inp[2]) ? 40'b0001001000000100000100000011000000001000 : 40'b1001001000010100000000000001000000001000;
												assign node422 = (inp[13]) ? 40'b0000001000010100000000000001000000001000 : 40'b0000001000010100000000000001100000001000;
										assign node425 = (inp[15]) ? node433 : node426;
											assign node426 = (inp[12]) ? node430 : node427;
												assign node427 = (inp[5]) ? 40'b0000001000010000000100000010100000001000 : 40'b0000001000011000000100000010100000001000;
												assign node430 = (inp[6]) ? 40'b0000001000011000000000000011000000001000 : 40'b0000001000011000000100000010000000001000;
											assign node433 = (inp[0]) ? node437 : node434;
												assign node434 = (inp[6]) ? 40'b0001001000001000000000000010000000001000 : 40'b1001001000000000000100000010000000001000;
												assign node437 = (inp[13]) ? 40'b0000001000000000000100000010000000001000 : 40'b1000001000001000000000000010100000001000;
								assign node440 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node441;
									assign node441 = (inp[10]) ? node457 : node442;
										assign node442 = (inp[12]) ? node450 : node443;
											assign node443 = (inp[6]) ? node447 : node444;
												assign node444 = (inp[15]) ? 40'b1001001000000100000100000010100000000000 : 40'b1001001000010100000100000010100000000000;
												assign node447 = (inp[13]) ? 40'b1000001000011100000000000010000000000000 : 40'b1001001000001100000000000010100000000000;
											assign node450 = (inp[0]) ? node454 : node451;
												assign node451 = (inp[6]) ? 40'b0001001000001100000000000011100000000000 : 40'b0001001000001100000100000010100000000000;
												assign node454 = (inp[15]) ? 40'b0000001000001100000000000010100000000000 : 40'b0000001000011100000000000011100000000000;
										assign node457 = (inp[15]) ? node465 : node458;
											assign node458 = (inp[0]) ? node462 : node459;
												assign node459 = (inp[5]) ? 40'b1001001000010000000100000010000000000000 : 40'b1001001000011000000000000010000000000000;
												assign node462 = (inp[2]) ? 40'b0000001000011000000000000011000000000000 : 40'b1000001000010000000000000001000000000000;
											assign node465 = (inp[12]) ? node467 : 40'b1001001000000000000100000010000000000000;
												assign node467 = (inp[2]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000001000000000000011100000000000;

endmodule