module dtc_split5_bm81 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node361;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node814;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node830;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node974;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node989;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1139;
	wire [3-1:0] node1143;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1151;
	wire [3-1:0] node1154;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1163;
	wire [3-1:0] node1167;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1176;

	assign outp = (inp[9]) ? node366 : node1;
		assign node1 = (inp[6]) ? node261 : node2;
			assign node2 = (inp[3]) ? node186 : node3;
				assign node3 = (inp[4]) ? node85 : node4;
					assign node4 = (inp[7]) ? node18 : node5;
						assign node5 = (inp[11]) ? 3'b001 : node6;
							assign node6 = (inp[8]) ? node8 : 3'b001;
								assign node8 = (inp[5]) ? node10 : 3'b001;
									assign node10 = (inp[10]) ? 3'b001 : node11;
										assign node11 = (inp[1]) ? 3'b000 : node12;
											assign node12 = (inp[0]) ? 3'b000 : 3'b001;
						assign node18 = (inp[10]) ? node50 : node19;
							assign node19 = (inp[5]) ? node37 : node20;
								assign node20 = (inp[8]) ? node30 : node21;
									assign node21 = (inp[11]) ? node25 : node22;
										assign node22 = (inp[2]) ? 3'b100 : 3'b000;
										assign node25 = (inp[1]) ? node27 : 3'b101;
											assign node27 = (inp[0]) ? 3'b001 : 3'b101;
									assign node30 = (inp[2]) ? node32 : 3'b000;
										assign node32 = (inp[1]) ? node34 : 3'b000;
											assign node34 = (inp[0]) ? 3'b100 : 3'b000;
								assign node37 = (inp[8]) ? node43 : node38;
									assign node38 = (inp[0]) ? node40 : 3'b000;
										assign node40 = (inp[1]) ? 3'b100 : 3'b000;
									assign node43 = (inp[0]) ? node45 : 3'b100;
										assign node45 = (inp[2]) ? node47 : 3'b100;
											assign node47 = (inp[11]) ? 3'b000 : 3'b100;
							assign node50 = (inp[5]) ? node68 : node51;
								assign node51 = (inp[8]) ? node61 : node52;
									assign node52 = (inp[11]) ? node56 : node53;
										assign node53 = (inp[0]) ? 3'b001 : 3'b101;
										assign node56 = (inp[0]) ? node58 : 3'b100;
											assign node58 = (inp[2]) ? 3'b100 : 3'b000;
									assign node61 = (inp[11]) ? node63 : 3'b001;
										assign node63 = (inp[0]) ? 3'b001 : node64;
											assign node64 = (inp[1]) ? 3'b001 : 3'b000;
								assign node68 = (inp[8]) ? node74 : node69;
									assign node69 = (inp[0]) ? node71 : 3'b001;
										assign node71 = (inp[1]) ? 3'b101 : 3'b001;
									assign node74 = (inp[11]) ? node80 : node75;
										assign node75 = (inp[2]) ? node77 : 3'b100;
											assign node77 = (inp[1]) ? 3'b000 : 3'b100;
										assign node80 = (inp[1]) ? node82 : 3'b101;
											assign node82 = (inp[2]) ? 3'b001 : 3'b101;
					assign node85 = (inp[7]) ? node149 : node86;
						assign node86 = (inp[10]) ? node124 : node87;
							assign node87 = (inp[8]) ? node105 : node88;
								assign node88 = (inp[11]) ? node94 : node89;
									assign node89 = (inp[0]) ? node91 : 3'b100;
										assign node91 = (inp[5]) ? 3'b010 : 3'b110;
									assign node94 = (inp[5]) ? node100 : node95;
										assign node95 = (inp[1]) ? 3'b001 : node96;
											assign node96 = (inp[0]) ? 3'b001 : 3'b100;
										assign node100 = (inp[0]) ? 3'b110 : node101;
											assign node101 = (inp[1]) ? 3'b100 : 3'b001;
								assign node105 = (inp[5]) ? node115 : node106;
									assign node106 = (inp[11]) ? node108 : 3'b010;
										assign node108 = (inp[0]) ? node112 : node109;
											assign node109 = (inp[1]) ? 3'b100 : 3'b001;
											assign node112 = (inp[1]) ? 3'b110 : 3'b100;
									assign node115 = (inp[11]) ? node121 : node116;
										assign node116 = (inp[0]) ? 3'b100 : node117;
											assign node117 = (inp[2]) ? 3'b110 : 3'b010;
										assign node121 = (inp[0]) ? 3'b010 : 3'b110;
							assign node124 = (inp[8]) ? node132 : node125;
								assign node125 = (inp[5]) ? node129 : node126;
									assign node126 = (inp[11]) ? 3'b011 : 3'b101;
									assign node129 = (inp[11]) ? 3'b101 : 3'b001;
								assign node132 = (inp[5]) ? node140 : node133;
									assign node133 = (inp[11]) ? 3'b101 : node134;
										assign node134 = (inp[1]) ? 3'b001 : node135;
											assign node135 = (inp[0]) ? 3'b001 : 3'b000;
									assign node140 = (inp[11]) ? node146 : node141;
										assign node141 = (inp[0]) ? 3'b110 : node142;
											assign node142 = (inp[1]) ? 3'b110 : 3'b001;
										assign node146 = (inp[0]) ? 3'b001 : 3'b101;
						assign node149 = (inp[10]) ? node163 : node150;
							assign node150 = (inp[8]) ? node158 : node151;
								assign node151 = (inp[5]) ? node155 : node152;
									assign node152 = (inp[11]) ? 3'b010 : 3'b100;
									assign node155 = (inp[11]) ? 3'b100 : 3'b000;
								assign node158 = (inp[11]) ? node160 : 3'b000;
									assign node160 = (inp[5]) ? 3'b000 : 3'b100;
							assign node163 = (inp[5]) ? node175 : node164;
								assign node164 = (inp[8]) ? node168 : node165;
									assign node165 = (inp[11]) ? 3'b001 : 3'b110;
									assign node168 = (inp[11]) ? node170 : 3'b010;
										assign node170 = (inp[0]) ? 3'b110 : node171;
											assign node171 = (inp[1]) ? 3'b110 : 3'b000;
								assign node175 = (inp[11]) ? node179 : node176;
									assign node176 = (inp[8]) ? 3'b100 : 3'b010;
									assign node179 = (inp[8]) ? 3'b010 : node180;
										assign node180 = (inp[2]) ? 3'b110 : node181;
											assign node181 = (inp[1]) ? 3'b110 : 3'b010;
				assign node186 = (inp[4]) ? node240 : node187;
					assign node187 = (inp[10]) ? node203 : node188;
						assign node188 = (inp[7]) ? 3'b000 : node189;
							assign node189 = (inp[8]) ? node197 : node190;
								assign node190 = (inp[5]) ? node194 : node191;
									assign node191 = (inp[11]) ? 3'b010 : 3'b100;
									assign node194 = (inp[11]) ? 3'b100 : 3'b000;
								assign node197 = (inp[11]) ? node199 : 3'b000;
									assign node199 = (inp[5]) ? 3'b000 : 3'b100;
						assign node203 = (inp[7]) ? node227 : node204;
							assign node204 = (inp[11]) ? node214 : node205;
								assign node205 = (inp[8]) ? node209 : node206;
									assign node206 = (inp[5]) ? 3'b010 : 3'b110;
									assign node209 = (inp[5]) ? node211 : 3'b010;
										assign node211 = (inp[1]) ? 3'b100 : 3'b110;
								assign node214 = (inp[5]) ? node222 : node215;
									assign node215 = (inp[8]) ? node217 : 3'b001;
										assign node217 = (inp[0]) ? 3'b110 : node218;
											assign node218 = (inp[2]) ? 3'b100 : 3'b000;
									assign node222 = (inp[8]) ? node224 : 3'b110;
										assign node224 = (inp[2]) ? 3'b010 : 3'b110;
							assign node227 = (inp[8]) ? node235 : node228;
								assign node228 = (inp[5]) ? node232 : node229;
									assign node229 = (inp[11]) ? 3'b010 : 3'b100;
									assign node232 = (inp[11]) ? 3'b100 : 3'b000;
								assign node235 = (inp[2]) ? node237 : 3'b000;
									assign node237 = (inp[11]) ? 3'b100 : 3'b000;
					assign node240 = (inp[10]) ? node242 : 3'b000;
						assign node242 = (inp[7]) ? 3'b000 : node243;
							assign node243 = (inp[11]) ? node249 : node244;
								assign node244 = (inp[8]) ? 3'b000 : node245;
									assign node245 = (inp[5]) ? 3'b000 : 3'b100;
								assign node249 = (inp[1]) ? 3'b100 : node250;
									assign node250 = (inp[0]) ? node254 : node251;
										assign node251 = (inp[5]) ? 3'b000 : 3'b100;
										assign node254 = (inp[5]) ? 3'b100 : node255;
											assign node255 = (inp[8]) ? 3'b100 : 3'b010;
			assign node261 = (inp[3]) ? 3'b000 : node262;
				assign node262 = (inp[7]) ? node342 : node263;
					assign node263 = (inp[10]) ? node295 : node264;
						assign node264 = (inp[4]) ? 3'b000 : node265;
							assign node265 = (inp[11]) ? node275 : node266;
								assign node266 = (inp[2]) ? 3'b000 : node267;
									assign node267 = (inp[5]) ? 3'b000 : node268;
										assign node268 = (inp[0]) ? 3'b100 : node269;
											assign node269 = (inp[8]) ? 3'b000 : 3'b000;
								assign node275 = (inp[8]) ? node283 : node276;
									assign node276 = (inp[5]) ? node280 : node277;
										assign node277 = (inp[0]) ? 3'b010 : 3'b110;
										assign node280 = (inp[0]) ? 3'b100 : 3'b000;
									assign node283 = (inp[2]) ? node289 : node284;
										assign node284 = (inp[0]) ? node286 : 3'b000;
											assign node286 = (inp[5]) ? 3'b000 : 3'b100;
										assign node289 = (inp[5]) ? node291 : 3'b100;
											assign node291 = (inp[0]) ? 3'b000 : 3'b100;
						assign node295 = (inp[4]) ? node329 : node296;
							assign node296 = (inp[11]) ? node314 : node297;
								assign node297 = (inp[8]) ? node305 : node298;
									assign node298 = (inp[0]) ? node302 : node299;
										assign node299 = (inp[2]) ? 3'b110 : 3'b011;
										assign node302 = (inp[2]) ? 3'b010 : 3'b110;
									assign node305 = (inp[5]) ? node309 : node306;
										assign node306 = (inp[2]) ? 3'b010 : 3'b110;
										assign node309 = (inp[1]) ? node311 : 3'b000;
											assign node311 = (inp[0]) ? 3'b100 : 3'b000;
								assign node314 = (inp[5]) ? node320 : node315;
									assign node315 = (inp[8]) ? 3'b011 : node316;
										assign node316 = (inp[0]) ? 3'b001 : 3'b101;
									assign node320 = (inp[8]) ? node326 : node321;
										assign node321 = (inp[0]) ? node323 : 3'b011;
											assign node323 = (inp[1]) ? 3'b110 : 3'b011;
										assign node326 = (inp[0]) ? 3'b010 : 3'b110;
							assign node329 = (inp[11]) ? node335 : node330;
								assign node330 = (inp[8]) ? 3'b000 : node331;
									assign node331 = (inp[5]) ? 3'b000 : 3'b100;
								assign node335 = (inp[8]) ? node339 : node336;
									assign node336 = (inp[5]) ? 3'b100 : 3'b010;
									assign node339 = (inp[5]) ? 3'b000 : 3'b100;
					assign node342 = (inp[4]) ? 3'b000 : node343;
						assign node343 = (inp[10]) ? node345 : 3'b000;
							assign node345 = (inp[11]) ? node351 : node346;
								assign node346 = (inp[8]) ? 3'b000 : node347;
									assign node347 = (inp[5]) ? 3'b000 : 3'b100;
								assign node351 = (inp[1]) ? node359 : node352;
									assign node352 = (inp[5]) ? node356 : node353;
										assign node353 = (inp[8]) ? 3'b100 : 3'b010;
										assign node356 = (inp[8]) ? 3'b000 : 3'b100;
									assign node359 = (inp[5]) ? node361 : 3'b100;
										assign node361 = (inp[0]) ? 3'b100 : 3'b000;
		assign node366 = (inp[3]) ? node778 : node367;
			assign node367 = (inp[6]) ? node503 : node368;
				assign node368 = (inp[10]) ? node478 : node369;
					assign node369 = (inp[7]) ? node407 : node370;
						assign node370 = (inp[4]) ? node372 : 3'b111;
							assign node372 = (inp[0]) ? node392 : node373;
								assign node373 = (inp[1]) ? node387 : node374;
									assign node374 = (inp[11]) ? node380 : node375;
										assign node375 = (inp[8]) ? node377 : 3'b111;
											assign node377 = (inp[2]) ? 3'b101 : 3'b011;
										assign node380 = (inp[5]) ? node384 : node381;
											assign node381 = (inp[8]) ? 3'b001 : 3'b101;
											assign node384 = (inp[8]) ? 3'b111 : 3'b011;
									assign node387 = (inp[11]) ? 3'b111 : node388;
										assign node388 = (inp[2]) ? 3'b111 : 3'b101;
								assign node392 = (inp[5]) ? node400 : node393;
									assign node393 = (inp[11]) ? node397 : node394;
										assign node394 = (inp[8]) ? 3'b011 : 3'b111;
										assign node397 = (inp[8]) ? 3'b111 : 3'b001;
									assign node400 = (inp[11]) ? node404 : node401;
										assign node401 = (inp[8]) ? 3'b101 : 3'b011;
										assign node404 = (inp[8]) ? 3'b011 : 3'b111;
						assign node407 = (inp[4]) ? node443 : node408;
							assign node408 = (inp[11]) ? node428 : node409;
								assign node409 = (inp[5]) ? node419 : node410;
									assign node410 = (inp[0]) ? node414 : node411;
										assign node411 = (inp[8]) ? 3'b111 : 3'b001;
										assign node414 = (inp[8]) ? node416 : 3'b111;
											assign node416 = (inp[1]) ? 3'b011 : 3'b111;
									assign node419 = (inp[8]) ? node423 : node420;
										assign node420 = (inp[0]) ? 3'b011 : 3'b111;
										assign node423 = (inp[2]) ? 3'b101 : node424;
											assign node424 = (inp[1]) ? 3'b101 : 3'b011;
								assign node428 = (inp[8]) ? node434 : node429;
									assign node429 = (inp[5]) ? 3'b001 : node430;
										assign node430 = (inp[0]) ? 3'b001 : 3'b101;
									assign node434 = (inp[5]) ? node438 : node435;
										assign node435 = (inp[1]) ? 3'b111 : 3'b001;
										assign node438 = (inp[1]) ? node440 : 3'b111;
											assign node440 = (inp[0]) ? 3'b011 : 3'b111;
							assign node443 = (inp[2]) ? node463 : node444;
								assign node444 = (inp[1]) ? node454 : node445;
									assign node445 = (inp[11]) ? 3'b101 : node446;
										assign node446 = (inp[8]) ? node450 : node447;
											assign node447 = (inp[5]) ? 3'b001 : 3'b101;
											assign node450 = (inp[5]) ? 3'b101 : 3'b001;
									assign node454 = (inp[11]) ? node458 : node455;
										assign node455 = (inp[5]) ? 3'b110 : 3'b101;
										assign node458 = (inp[5]) ? node460 : 3'b011;
											assign node460 = (inp[0]) ? 3'b001 : 3'b101;
								assign node463 = (inp[11]) ? node471 : node464;
									assign node464 = (inp[0]) ? 3'b001 : node465;
										assign node465 = (inp[8]) ? 3'b001 : node466;
											assign node466 = (inp[5]) ? 3'b001 : 3'b101;
									assign node471 = (inp[5]) ? node475 : node472;
										assign node472 = (inp[8]) ? 3'b101 : 3'b011;
										assign node475 = (inp[8]) ? 3'b001 : 3'b101;
					assign node478 = (inp[7]) ? node480 : 3'b111;
						assign node480 = (inp[4]) ? node482 : 3'b111;
							assign node482 = (inp[0]) ? node492 : node483;
								assign node483 = (inp[5]) ? node485 : 3'b111;
									assign node485 = (inp[11]) ? 3'b111 : node486;
										assign node486 = (inp[1]) ? node488 : 3'b111;
											assign node488 = (inp[8]) ? 3'b001 : 3'b011;
								assign node492 = (inp[11]) ? node498 : node493;
									assign node493 = (inp[2]) ? 3'b011 : node494;
										assign node494 = (inp[5]) ? 3'b011 : 3'b111;
									assign node498 = (inp[8]) ? node500 : 3'b111;
										assign node500 = (inp[5]) ? 3'b011 : 3'b111;
				assign node503 = (inp[10]) ? node641 : node504;
					assign node504 = (inp[7]) ? node574 : node505;
						assign node505 = (inp[4]) ? node545 : node506;
							assign node506 = (inp[11]) ? node526 : node507;
								assign node507 = (inp[5]) ? node515 : node508;
									assign node508 = (inp[8]) ? node510 : 3'b101;
										assign node510 = (inp[0]) ? 3'b001 : node511;
											assign node511 = (inp[1]) ? 3'b001 : 3'b101;
									assign node515 = (inp[8]) ? node519 : node516;
										assign node516 = (inp[0]) ? 3'b001 : 3'b101;
										assign node519 = (inp[0]) ? node523 : node520;
											assign node520 = (inp[2]) ? 3'b011 : 3'b001;
											assign node523 = (inp[1]) ? 3'b110 : 3'b111;
								assign node526 = (inp[8]) ? node534 : node527;
									assign node527 = (inp[5]) ? node531 : node528;
										assign node528 = (inp[0]) ? 3'b010 : 3'b110;
										assign node531 = (inp[0]) ? 3'b100 : 3'b000;
									assign node534 = (inp[5]) ? node540 : node535;
										assign node535 = (inp[0]) ? node537 : 3'b000;
											assign node537 = (inp[1]) ? 3'b101 : 3'b000;
										assign node540 = (inp[1]) ? node542 : 3'b101;
											assign node542 = (inp[0]) ? 3'b001 : 3'b101;
							assign node545 = (inp[11]) ? node555 : node546;
								assign node546 = (inp[8]) ? node552 : node547;
									assign node547 = (inp[0]) ? node549 : 3'b110;
										assign node549 = (inp[5]) ? 3'b010 : 3'b110;
									assign node552 = (inp[5]) ? 3'b100 : 3'b010;
								assign node555 = (inp[8]) ? node567 : node556;
									assign node556 = (inp[5]) ? node562 : node557;
										assign node557 = (inp[2]) ? 3'b001 : node558;
											assign node558 = (inp[0]) ? 3'b001 : 3'b111;
										assign node562 = (inp[0]) ? 3'b110 : node563;
											assign node563 = (inp[1]) ? 3'b000 : 3'b001;
									assign node567 = (inp[1]) ? 3'b110 : node568;
										assign node568 = (inp[5]) ? node570 : 3'b001;
											assign node570 = (inp[0]) ? 3'b010 : 3'b110;
						assign node574 = (inp[4]) ? node606 : node575;
							assign node575 = (inp[11]) ? node591 : node576;
								assign node576 = (inp[0]) ? node586 : node577;
									assign node577 = (inp[8]) ? 3'b010 : node578;
										assign node578 = (inp[1]) ? node582 : node579;
											assign node579 = (inp[5]) ? 3'b110 : 3'b010;
											assign node582 = (inp[2]) ? 3'b010 : 3'b110;
									assign node586 = (inp[5]) ? 3'b100 : node587;
										assign node587 = (inp[8]) ? 3'b010 : 3'b110;
								assign node591 = (inp[5]) ? node599 : node592;
									assign node592 = (inp[2]) ? 3'b001 : node593;
										assign node593 = (inp[1]) ? node595 : 3'b110;
											assign node595 = (inp[0]) ? 3'b001 : 3'b101;
									assign node599 = (inp[0]) ? node603 : node600;
										assign node600 = (inp[8]) ? 3'b110 : 3'b001;
										assign node603 = (inp[8]) ? 3'b010 : 3'b110;
							assign node606 = (inp[11]) ? node624 : node607;
								assign node607 = (inp[5]) ? node617 : node608;
									assign node608 = (inp[0]) ? 3'b100 : node609;
										assign node609 = (inp[2]) ? node613 : node610;
											assign node610 = (inp[8]) ? 3'b100 : 3'b000;
											assign node613 = (inp[8]) ? 3'b000 : 3'b000;
									assign node617 = (inp[8]) ? 3'b000 : node618;
										assign node618 = (inp[0]) ? 3'b000 : node619;
											assign node619 = (inp[2]) ? 3'b000 : 3'b100;
								assign node624 = (inp[5]) ? node630 : node625;
									assign node625 = (inp[2]) ? 3'b010 : node626;
										assign node626 = (inp[1]) ? 3'b100 : 3'b010;
									assign node630 = (inp[1]) ? node636 : node631;
										assign node631 = (inp[8]) ? 3'b100 : node632;
											assign node632 = (inp[0]) ? 3'b100 : 3'b010;
										assign node636 = (inp[0]) ? node638 : 3'b100;
											assign node638 = (inp[8]) ? 3'b000 : 3'b100;
					assign node641 = (inp[7]) ? node705 : node642;
						assign node642 = (inp[4]) ? node668 : node643;
							assign node643 = (inp[11]) ? 3'b111 : node644;
								assign node644 = (inp[8]) ? node654 : node645;
									assign node645 = (inp[5]) ? node649 : node646;
										assign node646 = (inp[1]) ? 3'b111 : 3'b011;
										assign node649 = (inp[0]) ? node651 : 3'b111;
											assign node651 = (inp[1]) ? 3'b011 : 3'b111;
									assign node654 = (inp[5]) ? node660 : node655;
										assign node655 = (inp[0]) ? node657 : 3'b111;
											assign node657 = (inp[1]) ? 3'b011 : 3'b111;
										assign node660 = (inp[0]) ? node664 : node661;
											assign node661 = (inp[2]) ? 3'b001 : 3'b011;
											assign node664 = (inp[1]) ? 3'b101 : 3'b001;
							assign node668 = (inp[5]) ? node690 : node669;
								assign node669 = (inp[0]) ? node681 : node670;
									assign node670 = (inp[1]) ? node678 : node671;
										assign node671 = (inp[8]) ? node675 : node672;
											assign node672 = (inp[11]) ? 3'b111 : 3'b011;
											assign node675 = (inp[11]) ? 3'b011 : 3'b111;
										assign node678 = (inp[11]) ? 3'b111 : 3'b101;
									assign node681 = (inp[11]) ? node685 : node682;
										assign node682 = (inp[8]) ? 3'b001 : 3'b101;
										assign node685 = (inp[8]) ? 3'b101 : node686;
											assign node686 = (inp[1]) ? 3'b011 : 3'b111;
								assign node690 = (inp[8]) ? node700 : node691;
									assign node691 = (inp[11]) ? node695 : node692;
										assign node692 = (inp[0]) ? 3'b001 : 3'b101;
										assign node695 = (inp[0]) ? node697 : 3'b011;
											assign node697 = (inp[1]) ? 3'b101 : 3'b001;
									assign node700 = (inp[11]) ? 3'b101 : node701;
										assign node701 = (inp[2]) ? 3'b001 : 3'b110;
						assign node705 = (inp[4]) ? node737 : node706;
							assign node706 = (inp[11]) ? node726 : node707;
								assign node707 = (inp[8]) ? node715 : node708;
									assign node708 = (inp[0]) ? node712 : node709;
										assign node709 = (inp[5]) ? 3'b101 : 3'b010;
										assign node712 = (inp[5]) ? 3'b001 : 3'b101;
									assign node715 = (inp[5]) ? node721 : node716;
										assign node716 = (inp[0]) ? node718 : 3'b101;
											assign node718 = (inp[1]) ? 3'b001 : 3'b101;
										assign node721 = (inp[0]) ? node723 : 3'b001;
											assign node723 = (inp[2]) ? 3'b110 : 3'b001;
								assign node726 = (inp[2]) ? 3'b011 : node727;
									assign node727 = (inp[5]) ? 3'b101 : node728;
										assign node728 = (inp[8]) ? node732 : node729;
											assign node729 = (inp[0]) ? 3'b011 : 3'b111;
											assign node732 = (inp[1]) ? 3'b101 : 3'b011;
							assign node737 = (inp[11]) ? node757 : node738;
								assign node738 = (inp[0]) ? node744 : node739;
									assign node739 = (inp[8]) ? node741 : 3'b001;
										assign node741 = (inp[5]) ? 3'b010 : 3'b110;
									assign node744 = (inp[5]) ? node750 : node745;
										assign node745 = (inp[8]) ? node747 : 3'b110;
											assign node747 = (inp[1]) ? 3'b010 : 3'b110;
										assign node750 = (inp[1]) ? node754 : node751;
											assign node751 = (inp[8]) ? 3'b010 : 3'b010;
											assign node754 = (inp[8]) ? 3'b100 : 3'b010;
								assign node757 = (inp[1]) ? node765 : node758;
									assign node758 = (inp[8]) ? node762 : node759;
										assign node759 = (inp[5]) ? 3'b001 : 3'b101;
										assign node762 = (inp[5]) ? 3'b110 : 3'b001;
									assign node765 = (inp[5]) ? node771 : node766;
										assign node766 = (inp[2]) ? node768 : 3'b001;
											assign node768 = (inp[0]) ? 3'b110 : 3'b001;
										assign node771 = (inp[8]) ? node775 : node772;
											assign node772 = (inp[0]) ? 3'b110 : 3'b001;
											assign node775 = (inp[0]) ? 3'b010 : 3'b110;
			assign node778 = (inp[6]) ? node1022 : node779;
				assign node779 = (inp[10]) ? node903 : node780;
					assign node780 = (inp[7]) ? node844 : node781;
						assign node781 = (inp[4]) ? node805 : node782;
							assign node782 = (inp[11]) ? node790 : node783;
								assign node783 = (inp[5]) ? node787 : node784;
									assign node784 = (inp[8]) ? 3'b001 : 3'b101;
									assign node787 = (inp[8]) ? 3'b110 : 3'b001;
								assign node790 = (inp[5]) ? node794 : node791;
									assign node791 = (inp[8]) ? 3'b101 : 3'b011;
									assign node794 = (inp[8]) ? node800 : node795;
										assign node795 = (inp[2]) ? 3'b101 : node796;
											assign node796 = (inp[1]) ? 3'b101 : 3'b001;
										assign node800 = (inp[2]) ? 3'b001 : node801;
											assign node801 = (inp[1]) ? 3'b001 : 3'b001;
							assign node805 = (inp[0]) ? node823 : node806;
								assign node806 = (inp[11]) ? node814 : node807;
									assign node807 = (inp[8]) ? node811 : node808;
										assign node808 = (inp[5]) ? 3'b010 : 3'b110;
										assign node811 = (inp[5]) ? 3'b100 : 3'b010;
									assign node814 = (inp[1]) ? node816 : 3'b001;
										assign node816 = (inp[5]) ? node820 : node817;
											assign node817 = (inp[8]) ? 3'b110 : 3'b001;
											assign node820 = (inp[8]) ? 3'b010 : 3'b110;
								assign node823 = (inp[2]) ? node835 : node824;
									assign node824 = (inp[8]) ? node830 : node825;
										assign node825 = (inp[11]) ? 3'b110 : node826;
											assign node826 = (inp[5]) ? 3'b010 : 3'b110;
										assign node830 = (inp[1]) ? node832 : 3'b010;
											assign node832 = (inp[11]) ? 3'b010 : 3'b100;
									assign node835 = (inp[11]) ? node839 : node836;
										assign node836 = (inp[5]) ? 3'b100 : 3'b110;
										assign node839 = (inp[1]) ? 3'b110 : node840;
											assign node840 = (inp[5]) ? 3'b010 : 3'b110;
						assign node844 = (inp[4]) ? node870 : node845;
							assign node845 = (inp[11]) ? node861 : node846;
								assign node846 = (inp[8]) ? node850 : node847;
									assign node847 = (inp[5]) ? 3'b010 : 3'b110;
									assign node850 = (inp[5]) ? node856 : node851;
										assign node851 = (inp[1]) ? 3'b010 : node852;
											assign node852 = (inp[0]) ? 3'b010 : 3'b010;
										assign node856 = (inp[0]) ? 3'b100 : node857;
											assign node857 = (inp[2]) ? 3'b100 : 3'b010;
								assign node861 = (inp[5]) ? node865 : node862;
									assign node862 = (inp[8]) ? 3'b110 : 3'b001;
									assign node865 = (inp[8]) ? node867 : 3'b110;
										assign node867 = (inp[0]) ? 3'b010 : 3'b110;
							assign node870 = (inp[11]) ? node882 : node871;
								assign node871 = (inp[8]) ? 3'b000 : node872;
									assign node872 = (inp[5]) ? node876 : node873;
										assign node873 = (inp[2]) ? 3'b100 : 3'b000;
										assign node876 = (inp[1]) ? 3'b000 : node877;
											assign node877 = (inp[2]) ? 3'b000 : 3'b000;
								assign node882 = (inp[5]) ? node894 : node883;
									assign node883 = (inp[8]) ? node889 : node884;
										assign node884 = (inp[0]) ? 3'b010 : node885;
											assign node885 = (inp[1]) ? 3'b010 : 3'b100;
										assign node889 = (inp[0]) ? 3'b100 : node890;
											assign node890 = (inp[1]) ? 3'b000 : 3'b010;
									assign node894 = (inp[8]) ? node900 : node895;
										assign node895 = (inp[1]) ? 3'b100 : node896;
											assign node896 = (inp[0]) ? 3'b100 : 3'b010;
										assign node900 = (inp[1]) ? 3'b000 : 3'b100;
					assign node903 = (inp[4]) ? node957 : node904;
						assign node904 = (inp[7]) ? node930 : node905;
							assign node905 = (inp[8]) ? node915 : node906;
								assign node906 = (inp[5]) ? node908 : 3'b111;
									assign node908 = (inp[11]) ? 3'b111 : node909;
										assign node909 = (inp[0]) ? 3'b011 : node910;
											assign node910 = (inp[1]) ? 3'b011 : 3'b111;
								assign node915 = (inp[5]) ? node923 : node916;
									assign node916 = (inp[11]) ? 3'b111 : node917;
										assign node917 = (inp[0]) ? 3'b011 : node918;
											assign node918 = (inp[2]) ? 3'b011 : 3'b111;
									assign node923 = (inp[11]) ? 3'b011 : node924;
										assign node924 = (inp[0]) ? 3'b101 : node925;
											assign node925 = (inp[1]) ? 3'b001 : 3'b011;
							assign node930 = (inp[11]) ? node946 : node931;
								assign node931 = (inp[8]) ? node939 : node932;
									assign node932 = (inp[0]) ? node936 : node933;
										assign node933 = (inp[5]) ? 3'b101 : 3'b011;
										assign node936 = (inp[5]) ? 3'b001 : 3'b101;
									assign node939 = (inp[5]) ? node943 : node940;
										assign node940 = (inp[0]) ? 3'b001 : 3'b101;
										assign node943 = (inp[0]) ? 3'b110 : 3'b001;
								assign node946 = (inp[5]) ? node948 : 3'b011;
									assign node948 = (inp[8]) ? node952 : node949;
										assign node949 = (inp[0]) ? 3'b101 : 3'b011;
										assign node952 = (inp[0]) ? node954 : 3'b101;
											assign node954 = (inp[1]) ? 3'b001 : 3'b101;
						assign node957 = (inp[7]) ? node983 : node958;
							assign node958 = (inp[0]) ? node974 : node959;
								assign node959 = (inp[11]) ? node969 : node960;
									assign node960 = (inp[2]) ? node966 : node961;
										assign node961 = (inp[5]) ? node963 : 3'b111;
											assign node963 = (inp[8]) ? 3'b001 : 3'b101;
										assign node966 = (inp[8]) ? 3'b110 : 3'b101;
									assign node969 = (inp[8]) ? 3'b011 : node970;
										assign node970 = (inp[1]) ? 3'b011 : 3'b111;
								assign node974 = (inp[8]) ? node976 : 3'b101;
									assign node976 = (inp[5]) ? node980 : node977;
										assign node977 = (inp[11]) ? 3'b101 : 3'b001;
										assign node980 = (inp[11]) ? 3'b001 : 3'b110;
							assign node983 = (inp[8]) ? node1001 : node984;
								assign node984 = (inp[0]) ? node992 : node985;
									assign node985 = (inp[11]) ? node989 : node986;
										assign node986 = (inp[5]) ? 3'b110 : 3'b001;
										assign node989 = (inp[5]) ? 3'b001 : 3'b101;
									assign node992 = (inp[11]) ? node996 : node993;
										assign node993 = (inp[5]) ? 3'b010 : 3'b110;
										assign node996 = (inp[5]) ? 3'b110 : node997;
											assign node997 = (inp[2]) ? 3'b001 : 3'b101;
								assign node1001 = (inp[1]) ? node1013 : node1002;
									assign node1002 = (inp[5]) ? node1010 : node1003;
										assign node1003 = (inp[0]) ? node1007 : node1004;
											assign node1004 = (inp[11]) ? 3'b001 : 3'b100;
											assign node1007 = (inp[2]) ? 3'b010 : 3'b000;
										assign node1010 = (inp[11]) ? 3'b110 : 3'b100;
									assign node1013 = (inp[5]) ? 3'b010 : node1014;
										assign node1014 = (inp[11]) ? node1018 : node1015;
											assign node1015 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1018 = (inp[0]) ? 3'b110 : 3'b001;
				assign node1022 = (inp[10]) ? node1080 : node1023;
					assign node1023 = (inp[4]) ? node1067 : node1024;
						assign node1024 = (inp[7]) ? node1058 : node1025;
							assign node1025 = (inp[11]) ? node1039 : node1026;
								assign node1026 = (inp[8]) ? 3'b000 : node1027;
									assign node1027 = (inp[2]) ? node1033 : node1028;
										assign node1028 = (inp[5]) ? node1030 : 3'b100;
											assign node1030 = (inp[0]) ? 3'b000 : 3'b100;
										assign node1033 = (inp[0]) ? 3'b100 : node1034;
											assign node1034 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1039 = (inp[5]) ? node1047 : node1040;
									assign node1040 = (inp[2]) ? 3'b010 : node1041;
										assign node1041 = (inp[0]) ? 3'b100 : node1042;
											assign node1042 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1047 = (inp[1]) ? node1053 : node1048;
										assign node1048 = (inp[0]) ? node1050 : 3'b100;
											assign node1050 = (inp[2]) ? 3'b110 : 3'b100;
										assign node1053 = (inp[2]) ? 3'b100 : node1054;
											assign node1054 = (inp[8]) ? 3'b000 : 3'b010;
							assign node1058 = (inp[5]) ? 3'b000 : node1059;
								assign node1059 = (inp[11]) ? node1061 : 3'b000;
									assign node1061 = (inp[0]) ? 3'b000 : node1062;
										assign node1062 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1067 = (inp[5]) ? 3'b000 : node1068;
							assign node1068 = (inp[1]) ? node1070 : 3'b000;
								assign node1070 = (inp[11]) ? node1072 : 3'b000;
									assign node1072 = (inp[2]) ? 3'b000 : node1073;
										assign node1073 = (inp[7]) ? 3'b000 : node1074;
											assign node1074 = (inp[0]) ? 3'b000 : 3'b100;
					assign node1080 = (inp[4]) ? node1146 : node1081;
						assign node1081 = (inp[7]) ? node1121 : node1082;
							assign node1082 = (inp[8]) ? node1096 : node1083;
								assign node1083 = (inp[0]) ? node1089 : node1084;
									assign node1084 = (inp[11]) ? node1086 : 3'b001;
										assign node1086 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1089 = (inp[11]) ? node1093 : node1090;
										assign node1090 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1093 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1096 = (inp[2]) ? node1108 : node1097;
									assign node1097 = (inp[1]) ? node1103 : node1098;
										assign node1098 = (inp[5]) ? 3'b110 : node1099;
											assign node1099 = (inp[11]) ? 3'b001 : 3'b110;
										assign node1103 = (inp[0]) ? node1105 : 3'b110;
											assign node1105 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1108 = (inp[11]) ? node1116 : node1109;
										assign node1109 = (inp[5]) ? node1113 : node1110;
											assign node1110 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1113 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1116 = (inp[1]) ? node1118 : 3'b001;
											assign node1118 = (inp[0]) ? 3'b110 : 3'b001;
							assign node1121 = (inp[11]) ? node1135 : node1122;
								assign node1122 = (inp[5]) ? node1128 : node1123;
									assign node1123 = (inp[8]) ? 3'b100 : node1124;
										assign node1124 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1128 = (inp[8]) ? 3'b000 : node1129;
										assign node1129 = (inp[0]) ? node1131 : 3'b100;
											assign node1131 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1135 = (inp[5]) ? node1143 : node1136;
									assign node1136 = (inp[8]) ? 3'b010 : node1137;
										assign node1137 = (inp[0]) ? node1139 : 3'b110;
											assign node1139 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1143 = (inp[8]) ? 3'b100 : 3'b010;
						assign node1146 = (inp[7]) ? node1170 : node1147;
							assign node1147 = (inp[11]) ? node1159 : node1148;
								assign node1148 = (inp[2]) ? node1154 : node1149;
									assign node1149 = (inp[8]) ? node1151 : 3'b100;
										assign node1151 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1154 = (inp[8]) ? node1156 : 3'b010;
										assign node1156 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1159 = (inp[8]) ? node1167 : node1160;
									assign node1160 = (inp[5]) ? 3'b010 : node1161;
										assign node1161 = (inp[1]) ? node1163 : 3'b110;
											assign node1163 = (inp[0]) ? 3'b010 : 3'b110;
									assign node1167 = (inp[5]) ? 3'b100 : 3'b010;
							assign node1170 = (inp[5]) ? 3'b000 : node1171;
								assign node1171 = (inp[11]) ? node1173 : 3'b000;
									assign node1173 = (inp[8]) ? 3'b000 : node1174;
										assign node1174 = (inp[0]) ? node1176 : 3'b100;
											assign node1176 = (inp[2]) ? 3'b000 : 3'b100;

endmodule