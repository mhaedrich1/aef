module dtc_split75_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node3;
	wire [40-1:0] node4;
	wire [40-1:0] node6;
	wire [40-1:0] node8;
	wire [40-1:0] node10;
	wire [40-1:0] node15;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node50;
	wire [40-1:0] node52;
	wire [40-1:0] node54;
	wire [40-1:0] node55;
	wire [40-1:0] node56;
	wire [40-1:0] node58;
	wire [40-1:0] node61;
	wire [40-1:0] node62;
	wire [40-1:0] node65;
	wire [40-1:0] node69;
	wire [40-1:0] node70;
	wire [40-1:0] node72;
	wire [40-1:0] node74;
	wire [40-1:0] node75;
	wire [40-1:0] node77;
	wire [40-1:0] node80;
	wire [40-1:0] node81;
	wire [40-1:0] node84;
	wire [40-1:0] node87;
	wire [40-1:0] node88;
	wire [40-1:0] node89;
	wire [40-1:0] node91;
	wire [40-1:0] node93;
	wire [40-1:0] node97;
	wire [40-1:0] node99;
	wire [40-1:0] node101;
	wire [40-1:0] node102;
	wire [40-1:0] node106;
	wire [40-1:0] node107;
	wire [40-1:0] node110;
	wire [40-1:0] node111;
	wire [40-1:0] node113;
	wire [40-1:0] node115;
	wire [40-1:0] node117;
	wire [40-1:0] node119;
	wire [40-1:0] node121;
	wire [40-1:0] node124;
	wire [40-1:0] node125;
	wire [40-1:0] node127;
	wire [40-1:0] node129;
	wire [40-1:0] node130;
	wire [40-1:0] node132;
	wire [40-1:0] node135;
	wire [40-1:0] node136;
	wire [40-1:0] node139;
	wire [40-1:0] node142;
	wire [40-1:0] node143;
	wire [40-1:0] node145;
	wire [40-1:0] node147;
	wire [40-1:0] node148;
	wire [40-1:0] node151;
	wire [40-1:0] node154;
	wire [40-1:0] node157;
	wire [40-1:0] node158;
	wire [40-1:0] node160;
	wire [40-1:0] node161;
	wire [40-1:0] node163;
	wire [40-1:0] node164;
	wire [40-1:0] node166;
	wire [40-1:0] node168;
	wire [40-1:0] node170;
	wire [40-1:0] node171;
	wire [40-1:0] node175;
	wire [40-1:0] node176;
	wire [40-1:0] node178;
	wire [40-1:0] node180;
	wire [40-1:0] node181;
	wire [40-1:0] node184;
	wire [40-1:0] node187;
	wire [40-1:0] node188;
	wire [40-1:0] node190;
	wire [40-1:0] node192;
	wire [40-1:0] node197;
	wire [40-1:0] node198;
	wire [40-1:0] node200;
	wire [40-1:0] node202;
	wire [40-1:0] node203;
	wire [40-1:0] node205;
	wire [40-1:0] node208;
	wire [40-1:0] node209;
	wire [40-1:0] node212;
	wire [40-1:0] node215;
	wire [40-1:0] node216;
	wire [40-1:0] node219;
	wire [40-1:0] node220;
	wire [40-1:0] node222;
	wire [40-1:0] node224;
	wire [40-1:0] node226;
	wire [40-1:0] node228;
	wire [40-1:0] node229;
	wire [40-1:0] node232;
	wire [40-1:0] node235;
	wire [40-1:0] node236;
	wire [40-1:0] node238;
	wire [40-1:0] node240;
	wire [40-1:0] node241;
	wire [40-1:0] node243;
	wire [40-1:0] node246;
	wire [40-1:0] node247;
	wire [40-1:0] node250;
	wire [40-1:0] node253;
	wire [40-1:0] node254;
	wire [40-1:0] node256;
	wire [40-1:0] node258;
	wire [40-1:0] node259;
	wire [40-1:0] node262;
	wire [40-1:0] node265;
	wire [40-1:0] node268;
	wire [40-1:0] node269;
	wire [40-1:0] node270;
	wire [40-1:0] node273;
	wire [40-1:0] node274;
	wire [40-1:0] node275;
	wire [40-1:0] node276;
	wire [40-1:0] node277;
	wire [40-1:0] node280;
	wire [40-1:0] node283;
	wire [40-1:0] node284;
	wire [40-1:0] node287;
	wire [40-1:0] node290;
	wire [40-1:0] node291;
	wire [40-1:0] node292;
	wire [40-1:0] node295;
	wire [40-1:0] node298;
	wire [40-1:0] node299;
	wire [40-1:0] node302;
	wire [40-1:0] node305;
	wire [40-1:0] node306;
	wire [40-1:0] node307;
	wire [40-1:0] node308;
	wire [40-1:0] node311;
	wire [40-1:0] node314;
	wire [40-1:0] node315;
	wire [40-1:0] node318;
	wire [40-1:0] node321;
	wire [40-1:0] node322;
	wire [40-1:0] node323;
	wire [40-1:0] node326;
	wire [40-1:0] node329;
	wire [40-1:0] node330;
	wire [40-1:0] node333;
	wire [40-1:0] node336;
	wire [40-1:0] node337;
	wire [40-1:0] node340;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node344;
	wire [40-1:0] node345;
	wire [40-1:0] node346;
	wire [40-1:0] node347;
	wire [40-1:0] node348;
	wire [40-1:0] node349;
	wire [40-1:0] node350;
	wire [40-1:0] node351;
	wire [40-1:0] node354;
	wire [40-1:0] node357;
	wire [40-1:0] node358;
	wire [40-1:0] node361;
	wire [40-1:0] node364;
	wire [40-1:0] node365;
	wire [40-1:0] node366;
	wire [40-1:0] node369;
	wire [40-1:0] node372;
	wire [40-1:0] node373;
	wire [40-1:0] node376;
	wire [40-1:0] node379;
	wire [40-1:0] node380;
	wire [40-1:0] node381;
	wire [40-1:0] node382;
	wire [40-1:0] node385;
	wire [40-1:0] node388;
	wire [40-1:0] node389;
	wire [40-1:0] node392;
	wire [40-1:0] node395;
	wire [40-1:0] node396;
	wire [40-1:0] node397;
	wire [40-1:0] node400;
	wire [40-1:0] node403;
	wire [40-1:0] node404;
	wire [40-1:0] node407;
	wire [40-1:0] node410;
	wire [40-1:0] node411;
	wire [40-1:0] node412;
	wire [40-1:0] node413;
	wire [40-1:0] node414;
	wire [40-1:0] node417;
	wire [40-1:0] node420;
	wire [40-1:0] node421;
	wire [40-1:0] node424;
	wire [40-1:0] node427;
	wire [40-1:0] node428;
	wire [40-1:0] node429;
	wire [40-1:0] node432;
	wire [40-1:0] node435;
	wire [40-1:0] node436;
	wire [40-1:0] node439;
	wire [40-1:0] node442;
	wire [40-1:0] node443;
	wire [40-1:0] node444;
	wire [40-1:0] node445;
	wire [40-1:0] node448;
	wire [40-1:0] node451;
	wire [40-1:0] node452;
	wire [40-1:0] node455;
	wire [40-1:0] node458;
	wire [40-1:0] node459;
	wire [40-1:0] node460;
	wire [40-1:0] node463;
	wire [40-1:0] node466;
	wire [40-1:0] node467;
	wire [40-1:0] node470;
	wire [40-1:0] node473;
	wire [40-1:0] node474;
	wire [40-1:0] node475;
	wire [40-1:0] node476;
	wire [40-1:0] node477;
	wire [40-1:0] node478;
	wire [40-1:0] node481;
	wire [40-1:0] node484;
	wire [40-1:0] node485;
	wire [40-1:0] node488;
	wire [40-1:0] node491;
	wire [40-1:0] node492;
	wire [40-1:0] node493;
	wire [40-1:0] node496;
	wire [40-1:0] node499;
	wire [40-1:0] node500;
	wire [40-1:0] node503;
	wire [40-1:0] node506;
	wire [40-1:0] node507;
	wire [40-1:0] node508;
	wire [40-1:0] node509;
	wire [40-1:0] node512;
	wire [40-1:0] node515;
	wire [40-1:0] node516;
	wire [40-1:0] node519;
	wire [40-1:0] node522;
	wire [40-1:0] node523;
	wire [40-1:0] node524;
	wire [40-1:0] node527;
	wire [40-1:0] node530;
	wire [40-1:0] node531;
	wire [40-1:0] node534;
	wire [40-1:0] node537;
	wire [40-1:0] node538;
	wire [40-1:0] node539;
	wire [40-1:0] node540;
	wire [40-1:0] node541;
	wire [40-1:0] node544;
	wire [40-1:0] node547;
	wire [40-1:0] node548;
	wire [40-1:0] node551;
	wire [40-1:0] node554;
	wire [40-1:0] node555;
	wire [40-1:0] node556;
	wire [40-1:0] node559;
	wire [40-1:0] node562;
	wire [40-1:0] node563;
	wire [40-1:0] node566;
	wire [40-1:0] node569;
	wire [40-1:0] node570;
	wire [40-1:0] node571;
	wire [40-1:0] node572;
	wire [40-1:0] node575;
	wire [40-1:0] node578;
	wire [40-1:0] node579;
	wire [40-1:0] node582;
	wire [40-1:0] node585;
	wire [40-1:0] node586;
	wire [40-1:0] node587;
	wire [40-1:0] node590;
	wire [40-1:0] node593;
	wire [40-1:0] node594;
	wire [40-1:0] node597;
	wire [40-1:0] node600;
	wire [40-1:0] node601;
	wire [40-1:0] node602;
	wire [40-1:0] node604;
	wire [40-1:0] node605;
	wire [40-1:0] node606;
	wire [40-1:0] node607;
	wire [40-1:0] node610;
	wire [40-1:0] node616;
	wire [40-1:0] node617;
	wire [40-1:0] node618;
	wire [40-1:0] node619;
	wire [40-1:0] node620;
	wire [40-1:0] node621;
	wire [40-1:0] node624;
	wire [40-1:0] node627;
	wire [40-1:0] node628;
	wire [40-1:0] node631;
	wire [40-1:0] node634;
	wire [40-1:0] node635;
	wire [40-1:0] node636;
	wire [40-1:0] node639;
	wire [40-1:0] node642;
	wire [40-1:0] node643;
	wire [40-1:0] node646;
	wire [40-1:0] node649;
	wire [40-1:0] node650;
	wire [40-1:0] node651;
	wire [40-1:0] node652;
	wire [40-1:0] node655;
	wire [40-1:0] node658;
	wire [40-1:0] node659;
	wire [40-1:0] node662;
	wire [40-1:0] node665;
	wire [40-1:0] node666;
	wire [40-1:0] node667;
	wire [40-1:0] node670;
	wire [40-1:0] node673;
	wire [40-1:0] node674;
	wire [40-1:0] node677;
	wire [40-1:0] node680;
	wire [40-1:0] node681;
	wire [40-1:0] node682;
	wire [40-1:0] node683;
	wire [40-1:0] node684;
	wire [40-1:0] node687;
	wire [40-1:0] node690;
	wire [40-1:0] node691;
	wire [40-1:0] node694;
	wire [40-1:0] node697;
	wire [40-1:0] node698;
	wire [40-1:0] node699;
	wire [40-1:0] node702;
	wire [40-1:0] node705;
	wire [40-1:0] node706;
	wire [40-1:0] node709;
	wire [40-1:0] node712;
	wire [40-1:0] node713;
	wire [40-1:0] node714;
	wire [40-1:0] node715;
	wire [40-1:0] node718;
	wire [40-1:0] node721;
	wire [40-1:0] node722;
	wire [40-1:0] node725;
	wire [40-1:0] node728;
	wire [40-1:0] node729;
	wire [40-1:0] node730;
	wire [40-1:0] node733;
	wire [40-1:0] node736;
	wire [40-1:0] node737;
	wire [40-1:0] node740;
	wire [40-1:0] node743;
	wire [40-1:0] node744;
	wire [40-1:0] node745;
	wire [40-1:0] node746;
	wire [40-1:0] node748;
	wire [40-1:0] node749;
	wire [40-1:0] node750;
	wire [40-1:0] node751;
	wire [40-1:0] node754;
	wire [40-1:0] node757;
	wire [40-1:0] node758;
	wire [40-1:0] node761;
	wire [40-1:0] node764;
	wire [40-1:0] node765;
	wire [40-1:0] node766;
	wire [40-1:0] node771;
	wire [40-1:0] node772;
	wire [40-1:0] node773;
	wire [40-1:0] node775;
	wire [40-1:0] node776;
	wire [40-1:0] node780;
	wire [40-1:0] node781;
	wire [40-1:0] node782;
	wire [40-1:0] node785;
	wire [40-1:0] node788;
	wire [40-1:0] node789;
	wire [40-1:0] node795;
	wire [40-1:0] node796;
	wire [40-1:0] node798;
	wire [40-1:0] node799;
	wire [40-1:0] node801;
	wire [40-1:0] node803;
	wire [40-1:0] node804;
	wire [40-1:0] node807;
	wire [40-1:0] node811;
	wire [40-1:0] node812;
	wire [40-1:0] node813;
	wire [40-1:0] node814;
	wire [40-1:0] node815;
	wire [40-1:0] node816;
	wire [40-1:0] node819;
	wire [40-1:0] node822;
	wire [40-1:0] node823;
	wire [40-1:0] node826;
	wire [40-1:0] node829;
	wire [40-1:0] node830;
	wire [40-1:0] node831;
	wire [40-1:0] node834;
	wire [40-1:0] node837;
	wire [40-1:0] node838;
	wire [40-1:0] node841;
	wire [40-1:0] node844;
	wire [40-1:0] node845;
	wire [40-1:0] node846;
	wire [40-1:0] node847;
	wire [40-1:0] node850;
	wire [40-1:0] node853;
	wire [40-1:0] node854;
	wire [40-1:0] node857;
	wire [40-1:0] node860;
	wire [40-1:0] node861;
	wire [40-1:0] node862;
	wire [40-1:0] node865;
	wire [40-1:0] node868;
	wire [40-1:0] node869;
	wire [40-1:0] node872;
	wire [40-1:0] node875;
	wire [40-1:0] node876;
	wire [40-1:0] node877;
	wire [40-1:0] node878;
	wire [40-1:0] node879;
	wire [40-1:0] node882;
	wire [40-1:0] node885;
	wire [40-1:0] node886;
	wire [40-1:0] node889;
	wire [40-1:0] node892;
	wire [40-1:0] node893;
	wire [40-1:0] node894;
	wire [40-1:0] node897;
	wire [40-1:0] node900;
	wire [40-1:0] node901;
	wire [40-1:0] node904;
	wire [40-1:0] node907;
	wire [40-1:0] node908;
	wire [40-1:0] node909;
	wire [40-1:0] node910;
	wire [40-1:0] node913;
	wire [40-1:0] node916;
	wire [40-1:0] node917;
	wire [40-1:0] node920;
	wire [40-1:0] node923;
	wire [40-1:0] node924;
	wire [40-1:0] node925;
	wire [40-1:0] node928;
	wire [40-1:0] node931;
	wire [40-1:0] node932;
	wire [40-1:0] node935;
	wire [40-1:0] node938;
	wire [40-1:0] node939;
	wire [40-1:0] node940;
	wire [40-1:0] node942;
	wire [40-1:0] node943;
	wire [40-1:0] node945;
	wire [40-1:0] node947;
	wire [40-1:0] node949;
	wire [40-1:0] node950;
	wire [40-1:0] node953;
	wire [40-1:0] node956;
	wire [40-1:0] node957;
	wire [40-1:0] node959;
	wire [40-1:0] node961;
	wire [40-1:0] node962;
	wire [40-1:0] node965;
	wire [40-1:0] node968;
	wire [40-1:0] node969;
	wire [40-1:0] node971;
	wire [40-1:0] node972;
	wire [40-1:0] node975;
	wire [40-1:0] node978;
	wire [40-1:0] node979;
	wire [40-1:0] node980;
	wire [40-1:0] node983;
	wire [40-1:0] node987;
	wire [40-1:0] node988;
	wire [40-1:0] node989;
	wire [40-1:0] node990;
	wire [40-1:0] node992;
	wire [40-1:0] node995;
	wire [40-1:0] node996;
	wire [40-1:0] node1000;
	wire [40-1:0] node1001;
	wire [40-1:0] node1003;
	wire [40-1:0] node1006;
	wire [40-1:0] node1007;
	wire [40-1:0] node1012;
	wire [40-1:0] node1013;
	wire [40-1:0] node1014;
	wire [40-1:0] node1016;
	wire [40-1:0] node1017;
	wire [40-1:0] node1018;
	wire [40-1:0] node1019;
	wire [40-1:0] node1020;
	wire [40-1:0] node1023;
	wire [40-1:0] node1026;
	wire [40-1:0] node1027;
	wire [40-1:0] node1030;
	wire [40-1:0] node1033;
	wire [40-1:0] node1034;
	wire [40-1:0] node1035;
	wire [40-1:0] node1038;
	wire [40-1:0] node1041;
	wire [40-1:0] node1042;
	wire [40-1:0] node1045;
	wire [40-1:0] node1048;
	wire [40-1:0] node1049;
	wire [40-1:0] node1050;
	wire [40-1:0] node1051;
	wire [40-1:0] node1054;
	wire [40-1:0] node1057;
	wire [40-1:0] node1058;
	wire [40-1:0] node1061;
	wire [40-1:0] node1064;
	wire [40-1:0] node1065;
	wire [40-1:0] node1066;
	wire [40-1:0] node1069;
	wire [40-1:0] node1072;
	wire [40-1:0] node1073;
	wire [40-1:0] node1076;
	wire [40-1:0] node1079;
	wire [40-1:0] node1080;
	wire [40-1:0] node1081;
	wire [40-1:0] node1082;
	wire [40-1:0] node1083;
	wire [40-1:0] node1084;
	wire [40-1:0] node1087;
	wire [40-1:0] node1090;
	wire [40-1:0] node1091;
	wire [40-1:0] node1094;
	wire [40-1:0] node1097;
	wire [40-1:0] node1098;
	wire [40-1:0] node1099;
	wire [40-1:0] node1102;
	wire [40-1:0] node1105;
	wire [40-1:0] node1106;
	wire [40-1:0] node1109;
	wire [40-1:0] node1112;
	wire [40-1:0] node1113;
	wire [40-1:0] node1114;
	wire [40-1:0] node1115;
	wire [40-1:0] node1118;
	wire [40-1:0] node1121;
	wire [40-1:0] node1122;
	wire [40-1:0] node1125;
	wire [40-1:0] node1128;
	wire [40-1:0] node1129;
	wire [40-1:0] node1130;
	wire [40-1:0] node1133;
	wire [40-1:0] node1136;
	wire [40-1:0] node1137;
	wire [40-1:0] node1140;
	wire [40-1:0] node1144;
	wire [40-1:0] node1145;
	wire [40-1:0] node1146;
	wire [40-1:0] node1147;
	wire [40-1:0] node1149;
	wire [40-1:0] node1150;
	wire [40-1:0] node1151;
	wire [40-1:0] node1154;
	wire [40-1:0] node1157;
	wire [40-1:0] node1158;
	wire [40-1:0] node1161;
	wire [40-1:0] node1164;
	wire [40-1:0] node1165;
	wire [40-1:0] node1166;
	wire [40-1:0] node1167;
	wire [40-1:0] node1170;
	wire [40-1:0] node1173;
	wire [40-1:0] node1174;
	wire [40-1:0] node1177;
	wire [40-1:0] node1181;
	wire [40-1:0] node1182;
	wire [40-1:0] node1183;
	wire [40-1:0] node1185;
	wire [40-1:0] node1186;
	wire [40-1:0] node1189;
	wire [40-1:0] node1192;
	wire [40-1:0] node1193;
	wire [40-1:0] node1194;
	wire [40-1:0] node1197;
	wire [40-1:0] node1201;
	wire [40-1:0] node1202;
	wire [40-1:0] node1204;
	wire [40-1:0] node1205;
	wire [40-1:0] node1208;
	wire [40-1:0] node1211;
	wire [40-1:0] node1212;
	wire [40-1:0] node1213;
	wire [40-1:0] node1216;
	wire [40-1:0] node1220;
	wire [40-1:0] node1221;
	wire [40-1:0] node1223;
	wire [40-1:0] node1224;
	wire [40-1:0] node1225;
	wire [40-1:0] node1226;
	wire [40-1:0] node1229;
	wire [40-1:0] node1232;
	wire [40-1:0] node1233;
	wire [40-1:0] node1236;
	wire [40-1:0] node1239;
	wire [40-1:0] node1240;
	wire [40-1:0] node1241;
	wire [40-1:0] node1244;
	wire [40-1:0] node1247;
	wire [40-1:0] node1248;
	wire [40-1:0] node1251;
	wire [40-1:0] node1254;
	wire [40-1:0] node1255;
	wire [40-1:0] node1256;
	wire [40-1:0] node1257;
	wire [40-1:0] node1258;
	wire [40-1:0] node1261;
	wire [40-1:0] node1264;
	wire [40-1:0] node1265;
	wire [40-1:0] node1268;
	wire [40-1:0] node1271;
	wire [40-1:0] node1272;
	wire [40-1:0] node1273;
	wire [40-1:0] node1276;
	wire [40-1:0] node1279;
	wire [40-1:0] node1280;
	wire [40-1:0] node1283;

	assign outp = (inp[9]) ? node268 : node1;
		assign node1 = (inp[1]) ? node15 : node2;
			assign node2 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node3;
				assign node3 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node4;
					assign node4 = (inp[7]) ? node6 : 40'b0000000000000000000000000000000000000000;
						assign node6 = (inp[8]) ? node8 : 40'b0000000000000000000000000000000000000000;
							assign node8 = (inp[4]) ? node10 : 40'b0000000000000000000000000000000000000000;
								assign node10 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
			assign node15 = (inp[4]) ? node17 : 40'b0000000001000000000000000000000000000000;
				assign node17 = (inp[7]) ? node157 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[3]) ? node24 : node21;
								assign node21 = (inp[11]) ? 40'b0000000000000010000001000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[11]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000100010000000000000000000000000;
							assign node27 = (inp[3]) ? node31 : node28;
								assign node28 = (inp[11]) ? 40'b0000000000000000000001000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[11]) ? node33 : 40'b0000000000100000000000000000000010000000;
									assign node33 = (inp[10]) ? node39 : node34;
										assign node34 = (inp[13]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[0]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[13]) ? node43 : node40;
											assign node40 = (inp[0]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000010000000;
						assign node46 = (inp[14]) ? node106 : node47;
							assign node47 = (inp[0]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[3]) ? node69 : node50;
									assign node50 = (inp[12]) ? node52 : 40'b0000000000000000000000000000000000000000;
										assign node52 = (inp[15]) ? node54 : 40'b0000000000000000000000000000000000000000;
											assign node54 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node55;
												assign node55 = (inp[6]) ? node61 : node56;
													assign node56 = (inp[5]) ? node58 : 40'b0000000000000000000000000000000000000000;
														assign node58 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node61 = (inp[10]) ? node65 : node62;
														assign node62 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node65 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node69 = (inp[13]) ? node87 : node70;
										assign node70 = (inp[12]) ? node72 : 40'b0000000000000000000000000000000000000000;
											assign node72 = (inp[15]) ? node74 : 40'b0000000000000000000000000000000000000000;
												assign node74 = (inp[2]) ? node80 : node75;
													assign node75 = (inp[5]) ? node77 : 40'b0000000000000000000000000000000000000000;
														assign node77 = (inp[6]) ? 40'b0000000010000000010000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node80 = (inp[10]) ? node84 : node81;
														assign node81 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000000000000010;
														assign node84 = (inp[6]) ? 40'b0000000000000000010000100000000010000010 : 40'b0000000000000000000000000000000000000000;
										assign node87 = (inp[11]) ? node97 : node88;
											assign node88 = (inp[10]) ? 40'b0000000000000000000000000000001000000000 : node89;
												assign node89 = (inp[15]) ? node91 : 40'b0000000000000000000000000000000000000000;
													assign node91 = (inp[12]) ? node93 : 40'b0000000000000000000000000000000000000000;
														assign node93 = (inp[2]) ? 40'b0000000000000010010000100000000000000000 : 40'b0000000010000010010000100000000000000000;
											assign node97 = (inp[15]) ? node99 : 40'b0000000000000000000000000000000000000000;
												assign node99 = (inp[12]) ? node101 : 40'b0000000000000000000000000000000000000000;
													assign node101 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node102;
														assign node102 = (inp[2]) ? 40'b0000000000000010010000100000010000000000 : 40'b0000000000000000000000000000000000000000;
							assign node106 = (inp[3]) ? node110 : node107;
								assign node107 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node110 = (inp[0]) ? node124 : node111;
									assign node111 = (inp[15]) ? node113 : 40'b0000000000000000000000000000000000000000;
										assign node113 = (inp[12]) ? node115 : 40'b0000000000000000000000000000000000000000;
											assign node115 = (inp[6]) ? node117 : 40'b0000000000000000000000000000000000000000;
												assign node117 = (inp[5]) ? node119 : 40'b0000000000000000000000000000000000000000;
													assign node119 = (inp[2]) ? node121 : 40'b0000000000000000000000000000000000000000;
														assign node121 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node124 = (inp[10]) ? node142 : node125;
										assign node125 = (inp[15]) ? node127 : 40'b0000000000000000000000000000000000000000;
											assign node127 = (inp[12]) ? node129 : 40'b0000000000000000000000000000000000000000;
												assign node129 = (inp[2]) ? node135 : node130;
													assign node130 = (inp[5]) ? node132 : 40'b0000000000000000000000000000000000000000;
														assign node132 = (inp[6]) ? 40'b0000000010001010010000100000000001000000 : 40'b0000000000000000000000000000000000000000;
													assign node135 = (inp[13]) ? node139 : node136;
														assign node136 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000000001000010;
														assign node139 = (inp[11]) ? 40'b0000000000001010010000100000000001000000 : 40'b0000000000000010010100100000000001000000;
										assign node142 = (inp[13]) ? node154 : node143;
											assign node143 = (inp[12]) ? node145 : 40'b0000000000000000000000000000000000000000;
												assign node145 = (inp[15]) ? node147 : 40'b0000000000000000000000000000000000000000;
													assign node147 = (inp[2]) ? node151 : node148;
														assign node148 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node151 = (inp[11]) ? 40'b0000000000001000010000100000000011000000 : 40'b0000000000000000010100100000000011000000;
											assign node154 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node157 = (inp[14]) ? node197 : node158;
						assign node158 = (inp[8]) ? node160 : 40'b0000000000000000000000000000000000000000;
							assign node160 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node161;
								assign node161 = (inp[0]) ? node163 : 40'b0000000000000000000000000000000000000000;
									assign node163 = (inp[3]) ? node175 : node164;
										assign node164 = (inp[12]) ? node166 : 40'b0000000000000000000000000000000000000000;
											assign node166 = (inp[13]) ? node168 : 40'b0000000000000000000000000000000000000000;
												assign node168 = (inp[15]) ? node170 : 40'b0000000000000000000000000000000000000000;
													assign node170 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node171;
														assign node171 = (inp[6]) ? 40'b0000000000000010000000100000000100000000 : 40'b0000000000000010000000100000001100000000;
										assign node175 = (inp[10]) ? node187 : node176;
											assign node176 = (inp[12]) ? node178 : 40'b0000000000000000000000000000000000000000;
												assign node178 = (inp[15]) ? node180 : 40'b0000000000000000000000000000000000000000;
													assign node180 = (inp[13]) ? node184 : node181;
														assign node181 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node184 = (inp[6]) ? 40'b0000000000000010000000100000000100000000 : 40'b0000000000000000000000000000000000000000;
											assign node187 = (inp[13]) ? 40'b0000000000000000000000010000000100000000 : node188;
												assign node188 = (inp[15]) ? node190 : 40'b0000000000000000000000000000000000000000;
													assign node190 = (inp[12]) ? node192 : 40'b0000000000000000000000000000000000000000;
														assign node192 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
						assign node197 = (inp[8]) ? node215 : node198;
							assign node198 = (inp[11]) ? node200 : 40'b0000000000000000000000000000000000000000;
								assign node200 = (inp[3]) ? node202 : 40'b0000000000000000000000000000000000000000;
									assign node202 = (inp[10]) ? node208 : node203;
										assign node203 = (inp[13]) ? node205 : 40'b0000000000000000000000000000000000000000;
											assign node205 = (inp[0]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node208 = (inp[13]) ? node212 : node209;
											assign node209 = (inp[0]) ? 40'b0000000000000000000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node212 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000110000000;
							assign node215 = (inp[3]) ? node219 : node216;
								assign node216 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node219 = (inp[0]) ? node235 : node220;
									assign node220 = (inp[5]) ? node222 : 40'b0000000000000000000000000000000000000000;
										assign node222 = (inp[12]) ? node224 : 40'b0000000000000000000000000000000000000000;
											assign node224 = (inp[15]) ? node226 : 40'b0000000000000000000000000000000000000000;
												assign node226 = (inp[2]) ? node228 : 40'b0000000000000000000000000000000000000000;
													assign node228 = (inp[11]) ? node232 : node229;
														assign node229 = (inp[6]) ? 40'b0100000000000000000000001000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node232 = (inp[10]) ? 40'b0100000000000000000000000000000000000001 : 40'b0000000000000000000000000000000000000000;
									assign node235 = (inp[13]) ? node253 : node236;
										assign node236 = (inp[15]) ? node238 : 40'b0000000000000000000000000000000000000000;
											assign node238 = (inp[12]) ? node240 : 40'b0000000000000000000000000000000000000000;
												assign node240 = (inp[6]) ? node246 : node241;
													assign node241 = (inp[5]) ? node243 : 40'b0000000000000000000000000000000000000000;
														assign node243 = (inp[2]) ? 40'b0100000000000000000000000000001100000001 : 40'b0000000000000000000000000000000000000000;
													assign node246 = (inp[10]) ? node250 : node247;
														assign node247 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000010000001000000000000000100000000;
														assign node250 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node253 = (inp[10]) ? node265 : node254;
											assign node254 = (inp[15]) ? node256 : 40'b0000000000000000000000000000000000000000;
												assign node256 = (inp[12]) ? node258 : 40'b0000000000000000000000000000000000000000;
													assign node258 = (inp[5]) ? node262 : node259;
														assign node259 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node262 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000010000010000000100000000100000000;
											assign node265 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node268 = (inp[1]) ? node336 : node269;
			assign node269 = (inp[8]) ? node273 : node270;
				assign node270 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node273 = (inp[7]) ? node305 : node274;
					assign node274 = (inp[3]) ? node290 : node275;
						assign node275 = (inp[11]) ? node283 : node276;
							assign node276 = (inp[14]) ? node280 : node277;
								assign node277 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node280 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
							assign node283 = (inp[14]) ? node287 : node284;
								assign node284 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node287 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
						assign node290 = (inp[11]) ? node298 : node291;
							assign node291 = (inp[14]) ? node295 : node292;
								assign node292 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node295 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
							assign node298 = (inp[14]) ? node302 : node299;
								assign node299 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
								assign node302 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node305 = (inp[14]) ? node321 : node306;
						assign node306 = (inp[3]) ? node314 : node307;
							assign node307 = (inp[11]) ? node311 : node308;
								assign node308 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node311 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
							assign node314 = (inp[11]) ? node318 : node315;
								assign node315 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node318 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
						assign node321 = (inp[11]) ? node329 : node322;
							assign node322 = (inp[3]) ? node326 : node323;
								assign node323 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node326 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
							assign node329 = (inp[3]) ? node333 : node330;
								assign node330 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
								assign node333 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node336 = (inp[4]) ? node340 : node337;
				assign node337 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node340 = (inp[8]) ? node342 : 40'b0000100000000000000000000000000000000000;
					assign node342 = (inp[7]) ? node938 : node343;
						assign node343 = (inp[3]) ? node743 : node344;
							assign node344 = (inp[14]) ? node600 : node345;
								assign node345 = (inp[13]) ? node473 : node346;
									assign node346 = (inp[0]) ? node410 : node347;
										assign node347 = (inp[15]) ? node379 : node348;
											assign node348 = (inp[10]) ? node364 : node349;
												assign node349 = (inp[11]) ? node357 : node350;
													assign node350 = (inp[2]) ? node354 : node351;
														assign node351 = (inp[5]) ? 40'b0001000000011101010110000010101000010000 : 40'b1001000000011101010010000010101000010000;
														assign node354 = (inp[12]) ? 40'b0001000000010101010010000001101000010000 : 40'b0001000000010101010110000010101000010000;
													assign node357 = (inp[5]) ? node361 : node358;
														assign node358 = (inp[6]) ? 40'b0001000000011101010010000010101000000000 : 40'b1001000000010101010010000000101000000000;
														assign node361 = (inp[6]) ? 40'b0001000000010101010010000011101000000000 : 40'b0001000000010101010110000010101000000000;
												assign node364 = (inp[11]) ? node372 : node365;
													assign node365 = (inp[6]) ? node369 : node366;
														assign node366 = (inp[5]) ? 40'b0001000000010001010110000010101000010000 : 40'b1001000000010001010010000000101000010000;
														assign node369 = (inp[12]) ? 40'b0001000000011001010010000011101000010000 : 40'b0001000000011001010010000010101000010000;
													assign node372 = (inp[6]) ? node376 : node373;
														assign node373 = (inp[5]) ? 40'b0001000000010001010110000010101000000000 : 40'b1001000000010001010010000000101000000000;
														assign node376 = (inp[5]) ? 40'b0001000000010001010010000011101000000000 : 40'b0001000000011001010010000010101000000000;
											assign node379 = (inp[10]) ? node395 : node380;
												assign node380 = (inp[11]) ? node388 : node381;
													assign node381 = (inp[12]) ? node385 : node382;
														assign node382 = (inp[6]) ? 40'b1001000000001101010010000010101000010000 : 40'b1001000000000101010110000010101000010000;
														assign node385 = (inp[2]) ? 40'b0001000000000101010010000001101000010000 : 40'b0001000000001101010010000010101000010000;
													assign node388 = (inp[12]) ? node392 : node389;
														assign node389 = (inp[2]) ? 40'b0001000000000101010110000010101000000000 : 40'b1001000000000101010010000000101000000000;
														assign node392 = (inp[2]) ? 40'b0001000000000101010010000011101000000000 : 40'b0001000000001101010010000010101000000000;
												assign node395 = (inp[11]) ? node403 : node396;
													assign node396 = (inp[2]) ? node400 : node397;
														assign node397 = (inp[12]) ? 40'b0001000000001001010010000010101000010000 : 40'b1001000000000001010010000010101000010000;
														assign node400 = (inp[12]) ? 40'b0001000000000001010010000001101000010000 : 40'b0001000000000001010110000010101000010000;
													assign node403 = (inp[12]) ? node407 : node404;
														assign node404 = (inp[2]) ? 40'b0001000000000001010110000010101000000000 : 40'b1001000000000001010010000000101000000000;
														assign node407 = (inp[2]) ? 40'b0001000000000001010010000001101000000000 : 40'b0001000000001001010010000010101000000000;
										assign node410 = (inp[15]) ? node442 : node411;
											assign node411 = (inp[11]) ? node427 : node412;
												assign node412 = (inp[10]) ? node420 : node413;
													assign node413 = (inp[2]) ? node417 : node414;
														assign node414 = (inp[12]) ? 40'b0000000000011101010010000010101000010000 : 40'b1000000000010101010010000010101000010000;
														assign node417 = (inp[12]) ? 40'b0000000000010101010010000001101000010000 : 40'b0000000000010101010110000010101000010000;
													assign node420 = (inp[12]) ? node424 : node421;
														assign node421 = (inp[2]) ? 40'b0000000000010001010110000010101000010000 : 40'b1000000000010001010010000000101000010000;
														assign node424 = (inp[2]) ? 40'b0000000000010001010010000001101000010000 : 40'b0000000000011001010010000010101000010000;
												assign node427 = (inp[10]) ? node435 : node428;
													assign node428 = (inp[2]) ? node432 : node429;
														assign node429 = (inp[12]) ? 40'b0000000000011101010010000010101000000000 : 40'b1000000000010101010010000000101000000000;
														assign node432 = (inp[12]) ? 40'b0000000000010101010010000001101000000000 : 40'b0000000000010101010110000010101000000000;
													assign node435 = (inp[6]) ? node439 : node436;
														assign node436 = (inp[5]) ? 40'b0000000000010001010110000010101000000000 : 40'b1000000000010001010010000000101000000000;
														assign node439 = (inp[5]) ? 40'b0000000000010001010010000001101000000000 : 40'b0000000000011001010010000010101000000000;
											assign node442 = (inp[11]) ? node458 : node443;
												assign node443 = (inp[10]) ? node451 : node444;
													assign node444 = (inp[12]) ? node448 : node445;
														assign node445 = (inp[6]) ? 40'b1000000000000101010010000001101000010000 : 40'b1000000000000101010110000010101000010000;
														assign node448 = (inp[2]) ? 40'b0000000000000101010010000001101000010000 : 40'b0000000000001101010010000010101000010000;
													assign node451 = (inp[12]) ? node455 : node452;
														assign node452 = (inp[2]) ? 40'b0000000000000001010110000010101000010000 : 40'b1000000000000001010010000000101000010000;
														assign node455 = (inp[2]) ? 40'b0000000000000001010010000011101000010000 : 40'b0000000000001001010010000010101000010000;
												assign node458 = (inp[10]) ? node466 : node459;
													assign node459 = (inp[12]) ? node463 : node460;
														assign node460 = (inp[2]) ? 40'b0000000000000101010110000010101000000000 : 40'b1000000000000101010010000000101000000000;
														assign node463 = (inp[6]) ? 40'b0000000000001101010010000011101000000000 : 40'b0000000000001101010110000010101000000000;
													assign node466 = (inp[12]) ? node470 : node467;
														assign node467 = (inp[2]) ? 40'b0000000000000001010110000010101000000000 : 40'b1000000000000001010010000010101000000000;
														assign node470 = (inp[2]) ? 40'b0000000000000001010010000001101000000000 : 40'b0000000000001001010010000010101000000000;
									assign node473 = (inp[11]) ? node537 : node474;
										assign node474 = (inp[15]) ? node506 : node475;
											assign node475 = (inp[10]) ? node491 : node476;
												assign node476 = (inp[0]) ? node484 : node477;
													assign node477 = (inp[2]) ? node481 : node478;
														assign node478 = (inp[12]) ? 40'b0001000000011101010010000010001000010000 : 40'b1001000000010101010010000000001000010000;
														assign node481 = (inp[12]) ? 40'b0001000000010101010010000001001000010000 : 40'b0001000000010101010110000010001000010000;
													assign node484 = (inp[5]) ? node488 : node485;
														assign node485 = (inp[6]) ? 40'b0000000000011101010010000010001000010000 : 40'b1000000000010101010010000000001000010000;
														assign node488 = (inp[2]) ? 40'b0000000000010101010110000011001000010000 : 40'b0000000000011101010110000010001000010000;
												assign node491 = (inp[0]) ? node499 : node492;
													assign node492 = (inp[6]) ? node496 : node493;
														assign node493 = (inp[5]) ? 40'b0001000000010001010110000010001000010000 : 40'b1001000000010001010010000000001000010000;
														assign node496 = (inp[12]) ? 40'b0001000000011001010010000011001000010000 : 40'b1001000000011001010010000010001000010000;
													assign node499 = (inp[2]) ? node503 : node500;
														assign node500 = (inp[12]) ? 40'b0000000000011001010010000010001000010000 : 40'b1000000000010001010010000000001000010000;
														assign node503 = (inp[12]) ? 40'b0000000000010001010010000001001000010000 : 40'b0000000000010001010110000010001000010000;
											assign node506 = (inp[10]) ? node522 : node507;
												assign node507 = (inp[0]) ? node515 : node508;
													assign node508 = (inp[12]) ? node512 : node509;
														assign node509 = (inp[2]) ? 40'b0001000000000101010110000010001000010000 : 40'b1001000000000101010010000000001000010000;
														assign node512 = (inp[2]) ? 40'b0001000000000101010010000001001000010000 : 40'b0001000000001101010010000010001000010000;
													assign node515 = (inp[5]) ? node519 : node516;
														assign node516 = (inp[12]) ? 40'b0000000000001101010010000010001000010000 : 40'b1000000000000101010010000000001000010000;
														assign node519 = (inp[2]) ? 40'b0000000000000101010110000011001000010000 : 40'b0000000000001101010110000010001000010000;
												assign node522 = (inp[0]) ? node530 : node523;
													assign node523 = (inp[12]) ? node527 : node524;
														assign node524 = (inp[2]) ? 40'b0001000000000001010110000010001000010000 : 40'b1001000000000001010010000000001000010000;
														assign node527 = (inp[2]) ? 40'b0001000000000001010010000001001000010000 : 40'b0001000000001001010010000010001000010000;
													assign node530 = (inp[12]) ? node534 : node531;
														assign node531 = (inp[6]) ? 40'b1000000000000001010010000000001000010000 : 40'b1000000000000001010110000010001000010000;
														assign node534 = (inp[6]) ? 40'b0000000000001001010010000011001000010000 : 40'b0000000000001001010010000010001000010000;
										assign node537 = (inp[10]) ? node569 : node538;
											assign node538 = (inp[0]) ? node554 : node539;
												assign node539 = (inp[15]) ? node547 : node540;
													assign node540 = (inp[5]) ? node544 : node541;
														assign node541 = (inp[6]) ? 40'b0001000000011101010010000010001000000000 : 40'b1001000000010101010010000010001000000000;
														assign node544 = (inp[6]) ? 40'b0001000000010101010010000001001000000000 : 40'b0001000000010101010110000010001000000000;
													assign node547 = (inp[5]) ? node551 : node548;
														assign node548 = (inp[6]) ? 40'b0001000000001101010010000010001000000000 : 40'b1001000000000101010010000000001000000000;
														assign node551 = (inp[6]) ? 40'b0001000000000101010010000001001000000000 : 40'b0001000000000101010110000010001000000000;
												assign node554 = (inp[15]) ? node562 : node555;
													assign node555 = (inp[5]) ? node559 : node556;
														assign node556 = (inp[6]) ? 40'b0000000000011101010010000010001000000000 : 40'b1000000000010101010010000000001000000000;
														assign node559 = (inp[6]) ? 40'b0000000000010101010010000001001000000000 : 40'b0000000000010101010110000010001000000000;
													assign node562 = (inp[6]) ? node566 : node563;
														assign node563 = (inp[5]) ? 40'b0000000000000101010110000010001000000000 : 40'b1000000000000101010010000000001000000000;
														assign node566 = (inp[2]) ? 40'b0000000000000101010010000011001000000000 : 40'b0000000000001101010010000010001000000000;
											assign node569 = (inp[0]) ? node585 : node570;
												assign node570 = (inp[15]) ? node578 : node571;
													assign node571 = (inp[2]) ? node575 : node572;
														assign node572 = (inp[12]) ? 40'b0001000000011001010010000010001000000000 : 40'b1001000000010001010010000000001000000000;
														assign node575 = (inp[12]) ? 40'b0001000000010001010010000011001000000000 : 40'b0001000000010001010110000010001000000000;
													assign node578 = (inp[6]) ? node582 : node579;
														assign node579 = (inp[5]) ? 40'b0001000000000001010110000010001000000000 : 40'b1001000000000001010010000000001000000000;
														assign node582 = (inp[5]) ? 40'b0001000000000001010010000001001000000000 : 40'b0001000000001001010010000010001000000000;
												assign node585 = (inp[15]) ? node593 : node586;
													assign node586 = (inp[12]) ? node590 : node587;
														assign node587 = (inp[6]) ? 40'b0000000000010001010110000010001000000000 : 40'b0000000000010001010110000010001000000000;
														assign node590 = (inp[2]) ? 40'b0000000000010001010010000001001000000000 : 40'b0000000000011001010010000010001000000000;
													assign node593 = (inp[5]) ? node597 : node594;
														assign node594 = (inp[6]) ? 40'b0000000000001001010010000010001000000000 : 40'b1000000000000001010010000000001000000000;
														assign node597 = (inp[6]) ? 40'b0000000000000001010010000001001000000000 : 40'b0000000000000001010110000010001000000000;
								assign node600 = (inp[11]) ? node616 : node601;
									assign node601 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node602;
										assign node602 = (inp[2]) ? node604 : 40'b0000000000000000000000000000000000000000;
											assign node604 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node605;
												assign node605 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node606;
													assign node606 = (inp[15]) ? node610 : node607;
														assign node607 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b1001000000010000001000000000000000000000;
														assign node610 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0001000000000000001100000010000000000000;
									assign node616 = (inp[13]) ? node680 : node617;
										assign node617 = (inp[10]) ? node649 : node618;
											assign node618 = (inp[15]) ? node634 : node619;
												assign node619 = (inp[0]) ? node627 : node620;
													assign node620 = (inp[5]) ? node624 : node621;
														assign node621 = (inp[6]) ? 40'b0001010000011100000000000010100000000000 : 40'b1001010000010100000000000000100000000000;
														assign node624 = (inp[6]) ? 40'b0001010000010100000000000001100000000000 : 40'b0001010000010100000100000010100000000000;
													assign node627 = (inp[6]) ? node631 : node628;
														assign node628 = (inp[5]) ? 40'b0000010000010100000100000010100000000000 : 40'b1000010000010100000000000000100000000000;
														assign node631 = (inp[12]) ? 40'b0000010000011100000000000011100000000000 : 40'b0000010000010100000100000010100000000000;
												assign node634 = (inp[0]) ? node642 : node635;
													assign node635 = (inp[12]) ? node639 : node636;
														assign node636 = (inp[2]) ? 40'b0001010000000100000100000010100000000000 : 40'b1001010000000100000000000000100000000000;
														assign node639 = (inp[2]) ? 40'b0001010000000100000000000011100000000000 : 40'b0001010000001100000000000010100000000000;
													assign node642 = (inp[6]) ? node646 : node643;
														assign node643 = (inp[5]) ? 40'b0000010000000100000100000010100000000000 : 40'b1000010000000100000000000000100000000000;
														assign node646 = (inp[12]) ? 40'b0000010000001100000000000011100000000000 : 40'b0000010000001100000000000010100000000000;
											assign node649 = (inp[15]) ? node665 : node650;
												assign node650 = (inp[0]) ? node658 : node651;
													assign node651 = (inp[5]) ? node655 : node652;
														assign node652 = (inp[6]) ? 40'b0001010000011000000000000010100000000000 : 40'b1001010000010000000000000000100000000000;
														assign node655 = (inp[6]) ? 40'b0001010000010000000000000001100000000000 : 40'b0001010000010000000100000010100000000000;
													assign node658 = (inp[5]) ? node662 : node659;
														assign node659 = (inp[2]) ? 40'b0000010000010000000100000010100000000000 : 40'b1000010000011000000000000010100000000000;
														assign node662 = (inp[6]) ? 40'b0000010000010000000000000001100000000000 : 40'b0000010000010000000100000010100000000000;
												assign node665 = (inp[0]) ? node673 : node666;
													assign node666 = (inp[5]) ? node670 : node667;
														assign node667 = (inp[6]) ? 40'b0001010000001000000000000010100000000000 : 40'b1001010000000000000000000000100000000000;
														assign node670 = (inp[6]) ? 40'b0001010000000000000000000001100000000000 : 40'b0001010000000000000100000010100000000000;
													assign node673 = (inp[2]) ? node677 : node674;
														assign node674 = (inp[12]) ? 40'b0000010000001000000000000010100000000000 : 40'b1000010000000000000000000000100000000000;
														assign node677 = (inp[12]) ? 40'b0000010000000000000000000001100000000000 : 40'b0000010000000000000100000010100000000000;
										assign node680 = (inp[10]) ? node712 : node681;
											assign node681 = (inp[0]) ? node697 : node682;
												assign node682 = (inp[15]) ? node690 : node683;
													assign node683 = (inp[2]) ? node687 : node684;
														assign node684 = (inp[5]) ? 40'b1001010000010100000000000011000000000000 : 40'b1001010000011100000000000010000000000000;
														assign node687 = (inp[12]) ? 40'b0001010000010100000000000001000000000000 : 40'b0001010000010100000100000010000000000000;
													assign node690 = (inp[5]) ? node694 : node691;
														assign node691 = (inp[6]) ? 40'b1001010000001100000000000010000000000000 : 40'b1001010000000100000000000000000000000000;
														assign node694 = (inp[6]) ? 40'b0001010000000100000000000001000000000000 : 40'b0001010000000100000100000010000000000000;
												assign node697 = (inp[15]) ? node705 : node698;
													assign node698 = (inp[12]) ? node702 : node699;
														assign node699 = (inp[2]) ? 40'b0000010000010100000100000010000000000000 : 40'b1000010000010100000000000000000000000000;
														assign node702 = (inp[2]) ? 40'b0000010000010100000000000001000000000000 : 40'b0000010000011100000000000010000000000000;
													assign node705 = (inp[5]) ? node709 : node706;
														assign node706 = (inp[6]) ? 40'b0000010000001100000000000010000000000000 : 40'b1000010000000100000000000000000000000000;
														assign node709 = (inp[6]) ? 40'b0000010000000100000000000001000000000000 : 40'b0000010000000100000100000010000000000000;
											assign node712 = (inp[0]) ? node728 : node713;
												assign node713 = (inp[15]) ? node721 : node714;
													assign node714 = (inp[5]) ? node718 : node715;
														assign node715 = (inp[6]) ? 40'b0001010000011000000000000010000000000000 : 40'b1001010000010000000000000000000000000000;
														assign node718 = (inp[6]) ? 40'b0001010000010000000000000001000000000000 : 40'b0001010000010000000100000010000000000000;
													assign node721 = (inp[5]) ? node725 : node722;
														assign node722 = (inp[6]) ? 40'b0001010000001000000000000010000000000000 : 40'b1001010000000000000000000000000000000000;
														assign node725 = (inp[6]) ? 40'b0001010000000000000000000001000000000000 : 40'b0001010000000000000100000010000000000000;
												assign node728 = (inp[15]) ? node736 : node729;
													assign node729 = (inp[2]) ? node733 : node730;
														assign node730 = (inp[5]) ? 40'b0000010000010000000000000001000000000000 : 40'b1000010000011000000000000010000000000000;
														assign node733 = (inp[12]) ? 40'b0000010000010000000000000001000000000000 : 40'b0000010000010000000100000010000000000000;
													assign node736 = (inp[12]) ? node740 : node737;
														assign node737 = (inp[2]) ? 40'b0000010000000000000100000010000000000000 : 40'b1000010000000000000000000000000000000000;
														assign node740 = (inp[6]) ? 40'b0000010000001000000000000011000000000000 : 40'b0000010000000000000000000001000000000000;
							assign node743 = (inp[11]) ? node795 : node744;
								assign node744 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node745;
									assign node745 = (inp[15]) ? node771 : node746;
										assign node746 = (inp[13]) ? node748 : 40'b0000000000000000000000000000000000000000;
											assign node748 = (inp[2]) ? node764 : node749;
												assign node749 = (inp[0]) ? node757 : node750;
													assign node750 = (inp[10]) ? node754 : node751;
														assign node751 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node754 = (inp[5]) ? 40'b1001000000010000000000000000000000100000 : 40'b1001000000011000000000000010000000100000;
													assign node757 = (inp[10]) ? node761 : node758;
														assign node758 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100000000000000000000100000;
														assign node761 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node764 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node765;
													assign node765 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node766;
														assign node766 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node771 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node772;
											assign node772 = (inp[2]) ? node780 : node773;
												assign node773 = (inp[5]) ? node775 : 40'b0000000000000000000000000000000000000000;
													assign node775 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node776;
														assign node776 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node780 = (inp[12]) ? node788 : node781;
													assign node781 = (inp[0]) ? node785 : node782;
														assign node782 = (inp[10]) ? 40'b0001000000000000000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
														assign node785 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000100000100000010100000100000;
													assign node788 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node789;
														assign node789 = (inp[10]) ? 40'b0001000000000000000100000011100000100000 : 40'b0000000000000000000000000000000000000000;
								assign node795 = (inp[14]) ? node811 : node796;
									assign node796 = (inp[2]) ? node798 : 40'b0000000000000000000000000000000000000000;
										assign node798 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node799;
											assign node799 = (inp[5]) ? node801 : 40'b0000000000000000000000000000000000000000;
												assign node801 = (inp[12]) ? node803 : 40'b0000000000000000000000000000000000000000;
													assign node803 = (inp[15]) ? node807 : node804;
														assign node804 = (inp[0]) ? 40'b1000000000010100001000000000000000010000 : 40'b0000000000000000000000000000000000000000;
														assign node807 = (inp[10]) ? 40'b0001000000000000001100000010000000010000 : 40'b0000000000000000000000000000000000000000;
									assign node811 = (inp[10]) ? node875 : node812;
										assign node812 = (inp[13]) ? node844 : node813;
											assign node813 = (inp[0]) ? node829 : node814;
												assign node814 = (inp[15]) ? node822 : node815;
													assign node815 = (inp[2]) ? node819 : node816;
														assign node816 = (inp[12]) ? 40'b0011000000011100000000000010100000000000 : 40'b1011000000010100000000000000100000000000;
														assign node819 = (inp[12]) ? 40'b0011000000010100000000000001100000000000 : 40'b0011000000010100000100000010100000000000;
													assign node822 = (inp[5]) ? node826 : node823;
														assign node823 = (inp[6]) ? 40'b0011000000001100000000000010100000000000 : 40'b1011000000000100000000000000100000000000;
														assign node826 = (inp[6]) ? 40'b0011000000000100000000000001100000000000 : 40'b0011000000000100000100000010100000000000;
												assign node829 = (inp[15]) ? node837 : node830;
													assign node830 = (inp[2]) ? node834 : node831;
														assign node831 = (inp[12]) ? 40'b0010000000011100000000000010100000000000 : 40'b1010000000010100000000000000100000000000;
														assign node834 = (inp[12]) ? 40'b0010000000010100000000000011100000000000 : 40'b0010000000010100000100000010100000000000;
													assign node837 = (inp[6]) ? node841 : node838;
														assign node838 = (inp[5]) ? 40'b0010000000000100000100000010100000000000 : 40'b1010000000000100000000000000100000000000;
														assign node841 = (inp[5]) ? 40'b0010000000000100000000000001100000000000 : 40'b0010000000001100000000000010100000000000;
											assign node844 = (inp[15]) ? node860 : node845;
												assign node845 = (inp[0]) ? node853 : node846;
													assign node846 = (inp[12]) ? node850 : node847;
														assign node847 = (inp[2]) ? 40'b0011000000010100000100000010000000000000 : 40'b1011000000010100000000000010000000000000;
														assign node850 = (inp[2]) ? 40'b0011000000010100000000000001000000000000 : 40'b0011000000011100000000000010000000000000;
													assign node853 = (inp[2]) ? node857 : node854;
														assign node854 = (inp[12]) ? 40'b0010000000011100000000000010000000000000 : 40'b1010000000010100000000000000000000000000;
														assign node857 = (inp[12]) ? 40'b0010000000010100000000000001000000000000 : 40'b0010000000010100000100000010000000000000;
												assign node860 = (inp[0]) ? node868 : node861;
													assign node861 = (inp[5]) ? node865 : node862;
														assign node862 = (inp[6]) ? 40'b0011000000001100000000000010000000000000 : 40'b1011000000000100000000000000000000000000;
														assign node865 = (inp[2]) ? 40'b0011000000000100000100000011000000000000 : 40'b0011000000001100000000000010000000000000;
													assign node868 = (inp[6]) ? node872 : node869;
														assign node869 = (inp[5]) ? 40'b0010000000000100000100000010000000000000 : 40'b1010000000000100000100000010000000000000;
														assign node872 = (inp[5]) ? 40'b0010000000000100000000000001000000000000 : 40'b0010000000001100000000000010000000000000;
										assign node875 = (inp[0]) ? node907 : node876;
											assign node876 = (inp[13]) ? node892 : node877;
												assign node877 = (inp[15]) ? node885 : node878;
													assign node878 = (inp[5]) ? node882 : node879;
														assign node879 = (inp[12]) ? 40'b0011000000011000000000000010100000000000 : 40'b0011000000011000000000000010100000000000;
														assign node882 = (inp[6]) ? 40'b0011000000010000000000000001100000000000 : 40'b0011000000010000000100000010100000000000;
													assign node885 = (inp[5]) ? node889 : node886;
														assign node886 = (inp[6]) ? 40'b0011000000001000000000000010100000000000 : 40'b1011000000000000000000000000100000000000;
														assign node889 = (inp[6]) ? 40'b0011000000000000000000000001100000000000 : 40'b0011000000000000000100000010100000000000;
												assign node892 = (inp[15]) ? node900 : node893;
													assign node893 = (inp[5]) ? node897 : node894;
														assign node894 = (inp[6]) ? 40'b0011000000011000000000000010000000000000 : 40'b1011000000010000000000000000000000000000;
														assign node897 = (inp[6]) ? 40'b0011000000010000000000000011000000000000 : 40'b0011000000010000000100000010000000000000;
													assign node900 = (inp[12]) ? node904 : node901;
														assign node901 = (inp[2]) ? 40'b0011000000000000000100000010000000000000 : 40'b1011000000000000000000000000000000000000;
														assign node904 = (inp[2]) ? 40'b0011000000000000000000000001000000000000 : 40'b0011000000001000000000000010000000000000;
											assign node907 = (inp[15]) ? node923 : node908;
												assign node908 = (inp[13]) ? node916 : node909;
													assign node909 = (inp[6]) ? node913 : node910;
														assign node910 = (inp[5]) ? 40'b0010000000010000000100000010100000000000 : 40'b1010000000010000000000000000100000000000;
														assign node913 = (inp[12]) ? 40'b0010000000011000000000000011100000000000 : 40'b1010000000010000000000000000100000000000;
													assign node916 = (inp[6]) ? node920 : node917;
														assign node917 = (inp[5]) ? 40'b0010000000010000000100000010000000000000 : 40'b1010000000010000000000000000000000000000;
														assign node920 = (inp[5]) ? 40'b0010000000010000000000000001000000000000 : 40'b0010000000011000000000000010000000000000;
												assign node923 = (inp[13]) ? node931 : node924;
													assign node924 = (inp[12]) ? node928 : node925;
														assign node925 = (inp[2]) ? 40'b0010000000000000000100000010100000000000 : 40'b1010000000000000000000000000100000000000;
														assign node928 = (inp[2]) ? 40'b0010000000000000000000000001100000000000 : 40'b0010000000001000000000000010100000000000;
													assign node931 = (inp[6]) ? node935 : node932;
														assign node932 = (inp[12]) ? 40'b0010000000001000000000000010000000000000 : 40'b1010000000000000000100000010000000000000;
														assign node935 = (inp[5]) ? 40'b0010000000000000000000000001000000000000 : 40'b0010000000001000000000000010000000000000;
						assign node938 = (inp[3]) ? node1012 : node939;
							assign node939 = (inp[11]) ? node987 : node940;
								assign node940 = (inp[14]) ? node942 : 40'b0000000000000000000000000000000000000000;
									assign node942 = (inp[0]) ? node956 : node943;
										assign node943 = (inp[13]) ? node945 : 40'b0000000000000000000000000000000000000000;
											assign node945 = (inp[10]) ? node947 : 40'b0000000000000000000000000000000000000000;
												assign node947 = (inp[15]) ? node949 : 40'b0000000000000000000000000000000000000000;
													assign node949 = (inp[2]) ? node953 : node950;
														assign node950 = (inp[5]) ? 40'b1001001100000000000000000001000000000000 : 40'b1001001100001000000000000010000000000000;
														assign node953 = (inp[5]) ? 40'b0001001100000000000100000011000000000000 : 40'b0001001100000000000100000010000000000000;
										assign node956 = (inp[10]) ? node968 : node957;
											assign node957 = (inp[15]) ? node959 : 40'b0000000000000000000000000000000000000000;
												assign node959 = (inp[13]) ? node961 : 40'b0000000000000000000000000000000000000000;
													assign node961 = (inp[2]) ? node965 : node962;
														assign node962 = (inp[5]) ? 40'b1000001100000100000000000000000000000000 : 40'b1000001100001100000000000010000000000000;
														assign node965 = (inp[5]) ? 40'b0000001100000100000100000011000000000000 : 40'b0000001100000100000100000010000000000000;
											assign node968 = (inp[13]) ? node978 : node969;
												assign node969 = (inp[15]) ? node971 : 40'b0000000000000000000000000000000000000000;
													assign node971 = (inp[6]) ? node975 : node972;
														assign node972 = (inp[5]) ? 40'b0000001100000000000100000010100000000000 : 40'b1000001100000000000000000000100000000000;
														assign node975 = (inp[5]) ? 40'b0000001100000000000000000001100000000000 : 40'b0000001100001000000000000010100000000000;
												assign node978 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node979;
													assign node979 = (inp[5]) ? node983 : node980;
														assign node980 = (inp[6]) ? 40'b0000001100011000000000000010000000000000 : 40'b1000001100010000000000000010000000000000;
														assign node983 = (inp[6]) ? 40'b0000001100010000000000000001000000000000 : 40'b0000001100010000000100000010000000000000;
								assign node987 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node988;
									assign node988 = (inp[15]) ? node1000 : node989;
										assign node989 = (inp[10]) ? node995 : node990;
											assign node990 = (inp[0]) ? node992 : 40'b0000000000000000000000000000000000000000;
												assign node992 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
											assign node995 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node996;
												assign node996 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
										assign node1000 = (inp[0]) ? node1006 : node1001;
											assign node1001 = (inp[10]) ? node1003 : 40'b0000000000000000000000000000000000000000;
												assign node1003 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
											assign node1006 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node1007;
												assign node1007 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
							assign node1012 = (inp[0]) ? node1144 : node1013;
								assign node1013 = (inp[11]) ? node1079 : node1014;
									assign node1014 = (inp[14]) ? node1016 : 40'b0000000000000000000000000000000000000000;
										assign node1016 = (inp[15]) ? node1048 : node1017;
											assign node1017 = (inp[10]) ? node1033 : node1018;
												assign node1018 = (inp[13]) ? node1026 : node1019;
													assign node1019 = (inp[6]) ? node1023 : node1020;
														assign node1020 = (inp[5]) ? 40'b0001001000010100000100000010100000000000 : 40'b1001001000010100000000000000100000000000;
														assign node1023 = (inp[5]) ? 40'b0001001000010100000000000001100000000000 : 40'b0001001000011100000000000010100000000000;
													assign node1026 = (inp[2]) ? node1030 : node1027;
														assign node1027 = (inp[5]) ? 40'b0001001000011100000000000011000000000000 : 40'b1001001000011100000000000010000000000000;
														assign node1030 = (inp[12]) ? 40'b0001001000010100000000000011000000000000 : 40'b0001001000010100000100000010000000000000;
												assign node1033 = (inp[13]) ? node1041 : node1034;
													assign node1034 = (inp[12]) ? node1038 : node1035;
														assign node1035 = (inp[2]) ? 40'b0001001000010000000100000010100000000000 : 40'b1001001000010000000000000000100000000000;
														assign node1038 = (inp[2]) ? 40'b0001001000010000000000000011100000000000 : 40'b0001001000011000000000000010100000000000;
													assign node1041 = (inp[5]) ? node1045 : node1042;
														assign node1042 = (inp[2]) ? 40'b0001001000011000000100000010000000000000 : 40'b1001001000011000000000000010000000000000;
														assign node1045 = (inp[6]) ? 40'b0001001000010000000000000001000000000000 : 40'b0001001000010000000100000010000000000000;
											assign node1048 = (inp[13]) ? node1064 : node1049;
												assign node1049 = (inp[10]) ? node1057 : node1050;
													assign node1050 = (inp[2]) ? node1054 : node1051;
														assign node1051 = (inp[5]) ? 40'b0001001000001100000100000010100000000000 : 40'b1001001000001100000000000010100000000000;
														assign node1054 = (inp[12]) ? 40'b0001001000000100000000000001100000000000 : 40'b0001001000000100000100000010100000000000;
													assign node1057 = (inp[2]) ? node1061 : node1058;
														assign node1058 = (inp[12]) ? 40'b0001001000001000000000000010100000000000 : 40'b1001001000000000000000000000100000000000;
														assign node1061 = (inp[12]) ? 40'b0001001000000000000000000001100000000000 : 40'b0001001000000000000100000010100000000000;
												assign node1064 = (inp[10]) ? node1072 : node1065;
													assign node1065 = (inp[12]) ? node1069 : node1066;
														assign node1066 = (inp[2]) ? 40'b0001001000000100000100000010000000000000 : 40'b1001001000000100000000000000000000000000;
														assign node1069 = (inp[2]) ? 40'b0001001000000100000000000001000000000000 : 40'b0001001000001100000000000010000000000000;
													assign node1072 = (inp[2]) ? node1076 : node1073;
														assign node1073 = (inp[12]) ? 40'b0001001000001000000000000010000000000000 : 40'b1001001000000000000000000000000000000000;
														assign node1076 = (inp[12]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000000000000100000010000000000000;
									assign node1079 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node1080;
										assign node1080 = (inp[15]) ? node1112 : node1081;
											assign node1081 = (inp[13]) ? node1097 : node1082;
												assign node1082 = (inp[10]) ? node1090 : node1083;
													assign node1083 = (inp[5]) ? node1087 : node1084;
														assign node1084 = (inp[6]) ? 40'b0001001000011100000000000010100000001000 : 40'b1001001000010100000000000000100000001000;
														assign node1087 = (inp[6]) ? 40'b0001001000010100000000000001100000001000 : 40'b0001001000010100000100000010100000001000;
													assign node1090 = (inp[12]) ? node1094 : node1091;
														assign node1091 = (inp[2]) ? 40'b0001001000010000000100000010100000001000 : 40'b1001001000010000000000000000100000001000;
														assign node1094 = (inp[2]) ? 40'b0001001000010000000000000011100000001000 : 40'b0001001000011000000000000010100000001000;
												assign node1097 = (inp[10]) ? node1105 : node1098;
													assign node1098 = (inp[2]) ? node1102 : node1099;
														assign node1099 = (inp[12]) ? 40'b0001001000011100000000000010000000001000 : 40'b1001001000010100000000000000000000001000;
														assign node1102 = (inp[12]) ? 40'b0001001000010100000000000001000000001000 : 40'b0001001000010100000100000010000000001000;
													assign node1105 = (inp[2]) ? node1109 : node1106;
														assign node1106 = (inp[12]) ? 40'b0001001000011000000000000010000000001000 : 40'b1001001000010000000000000000000000001000;
														assign node1109 = (inp[12]) ? 40'b0001001000010000000000000001000000001000 : 40'b0001001000010000000100000010000000001000;
											assign node1112 = (inp[13]) ? node1128 : node1113;
												assign node1113 = (inp[10]) ? node1121 : node1114;
													assign node1114 = (inp[2]) ? node1118 : node1115;
														assign node1115 = (inp[12]) ? 40'b0001001000001100000000000010100000001000 : 40'b1001001000000100000000000000100000001000;
														assign node1118 = (inp[12]) ? 40'b0001001000000100000000000011100000001000 : 40'b0001001000000100000100000010100000001000;
													assign node1121 = (inp[5]) ? node1125 : node1122;
														assign node1122 = (inp[6]) ? 40'b0001001000001000000000000010100000001000 : 40'b1001001000000000000000000010100000001000;
														assign node1125 = (inp[6]) ? 40'b0001001000000000000000000001100000001000 : 40'b0001001000000000000100000010100000001000;
												assign node1128 = (inp[10]) ? node1136 : node1129;
													assign node1129 = (inp[12]) ? node1133 : node1130;
														assign node1130 = (inp[2]) ? 40'b0001001000000100000100000010000000001000 : 40'b1001001000000100000000000000000000001000;
														assign node1133 = (inp[2]) ? 40'b0001001000000100000000000001000000001000 : 40'b0001001000001100000000000010000000001000;
													assign node1136 = (inp[6]) ? node1140 : node1137;
														assign node1137 = (inp[5]) ? 40'b0001001000000000000100000010000000001000 : 40'b1001001000000000000000000000000000001000;
														assign node1140 = (inp[5]) ? 40'b0001001000000000000000000011000000001000 : 40'b0001001000001000000000000010000000001000;
								assign node1144 = (inp[10]) ? node1220 : node1145;
									assign node1145 = (inp[15]) ? node1181 : node1146;
										assign node1146 = (inp[14]) ? node1164 : node1147;
											assign node1147 = (inp[11]) ? node1149 : 40'b0000000000000000000000000000000000000000;
												assign node1149 = (inp[13]) ? node1157 : node1150;
													assign node1150 = (inp[2]) ? node1154 : node1151;
														assign node1151 = (inp[12]) ? 40'b0000001000011100000000000010100000001000 : 40'b1000001000010100000000000000100000001000;
														assign node1154 = (inp[12]) ? 40'b0000001000010100000000000001100000001000 : 40'b0000001000010100000100000010100000001000;
													assign node1157 = (inp[5]) ? node1161 : node1158;
														assign node1158 = (inp[6]) ? 40'b0000001000011100000000000010000000001000 : 40'b1000001000010100000000000000000000001000;
														assign node1161 = (inp[6]) ? 40'b0000001000010100000000000001000000001000 : 40'b0000001000010100000100000010000000001000;
											assign node1164 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1165;
												assign node1165 = (inp[13]) ? node1173 : node1166;
													assign node1166 = (inp[5]) ? node1170 : node1167;
														assign node1167 = (inp[6]) ? 40'b0000001000011100000000000010100000000000 : 40'b1000001000010100000000000000100000000000;
														assign node1170 = (inp[6]) ? 40'b0000001000010100000000000001100000000000 : 40'b0000001000010100000100000010100000000000;
													assign node1173 = (inp[12]) ? node1177 : node1174;
														assign node1174 = (inp[2]) ? 40'b0000001000010100000100000010000000000000 : 40'b1000001000010100000000000000000000000000;
														assign node1177 = (inp[2]) ? 40'b0000001000010100000000000001000000000000 : 40'b0000001000011100000000000010000000000000;
										assign node1181 = (inp[13]) ? node1201 : node1182;
											assign node1182 = (inp[14]) ? node1192 : node1183;
												assign node1183 = (inp[11]) ? node1185 : 40'b0000000000000000000000000000000000000000;
													assign node1185 = (inp[2]) ? node1189 : node1186;
														assign node1186 = (inp[12]) ? 40'b0000001000001100000000000010100000001000 : 40'b1000001000000100000000000000100000001000;
														assign node1189 = (inp[5]) ? 40'b0000001000000100000100000011100000001000 : 40'b0000001000000100000100000010100000001000;
												assign node1192 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1193;
													assign node1193 = (inp[6]) ? node1197 : node1194;
														assign node1194 = (inp[5]) ? 40'b0000001000000100000100000010100000000000 : 40'b1000001000000100000000000010100000000000;
														assign node1197 = (inp[5]) ? 40'b0000001000000100000000000001100000000000 : 40'b0000001000001100000000000010100000000000;
											assign node1201 = (inp[14]) ? node1211 : node1202;
												assign node1202 = (inp[11]) ? node1204 : 40'b0000000000000000000000000000000000000000;
													assign node1204 = (inp[2]) ? node1208 : node1205;
														assign node1205 = (inp[12]) ? 40'b0000001000001100000100000010000000001000 : 40'b1000001000000100000000000000000000001000;
														assign node1208 = (inp[12]) ? 40'b0000001000000100000000000011000000001000 : 40'b0000001000000100000100000010000000001000;
												assign node1211 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1212;
													assign node1212 = (inp[2]) ? node1216 : node1213;
														assign node1213 = (inp[12]) ? 40'b0000001000001100000000000010000000000000 : 40'b1000001000000100000000000000000000000000;
														assign node1216 = (inp[12]) ? 40'b0000001000000100000000000011000000000000 : 40'b0000001000000100000100000010000000000000;
									assign node1220 = (inp[14]) ? node1254 : node1221;
										assign node1221 = (inp[11]) ? node1223 : 40'b0000000000000000000000000000000000000000;
											assign node1223 = (inp[15]) ? node1239 : node1224;
												assign node1224 = (inp[13]) ? node1232 : node1225;
													assign node1225 = (inp[12]) ? node1229 : node1226;
														assign node1226 = (inp[2]) ? 40'b0000001000010000000100000010100000001000 : 40'b1000001000010000000000000000100000001000;
														assign node1229 = (inp[5]) ? 40'b0000001000010000000000000001100000001000 : 40'b0000001000011000000000000010100000001000;
													assign node1232 = (inp[6]) ? node1236 : node1233;
														assign node1233 = (inp[5]) ? 40'b0000001000010000000100000010000000001000 : 40'b1000001000010000000000000000000000001000;
														assign node1236 = (inp[5]) ? 40'b0000001000010000000000000001000000001000 : 40'b0000001000011000000000000010000000001000;
												assign node1239 = (inp[13]) ? node1247 : node1240;
													assign node1240 = (inp[2]) ? node1244 : node1241;
														assign node1241 = (inp[12]) ? 40'b0000001000001000000000000010100000001000 : 40'b1000001000000000000000000000100000001000;
														assign node1244 = (inp[5]) ? 40'b0000001000000000000100000011100000001000 : 40'b1000001000000000000000000000100000001000;
													assign node1247 = (inp[2]) ? node1251 : node1248;
														assign node1248 = (inp[12]) ? 40'b0000001000001000000000000010000000001000 : 40'b1000001000000000000000000000000000001000;
														assign node1251 = (inp[12]) ? 40'b0000001000000000000000000001000000001000 : 40'b0000001000000000000100000010000000001000;
										assign node1254 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1255;
											assign node1255 = (inp[15]) ? node1271 : node1256;
												assign node1256 = (inp[13]) ? node1264 : node1257;
													assign node1257 = (inp[6]) ? node1261 : node1258;
														assign node1258 = (inp[5]) ? 40'b0000001000010000000100000010100000000000 : 40'b1000001000010000000000000000100000000000;
														assign node1261 = (inp[12]) ? 40'b0000001000011000000000000011100000000000 : 40'b0000001000010000000000000001100000000000;
													assign node1264 = (inp[2]) ? node1268 : node1265;
														assign node1265 = (inp[5]) ? 40'b1000001000010000000000000000000000000000 : 40'b1000001000011000000000000010000000000000;
														assign node1268 = (inp[12]) ? 40'b0000001000010000000000000001000000000000 : 40'b0000001000010000000100000010000000000000;
												assign node1271 = (inp[13]) ? node1279 : node1272;
													assign node1272 = (inp[6]) ? node1276 : node1273;
														assign node1273 = (inp[12]) ? 40'b0000001000001000000100000010100000000000 : 40'b1000001000000000000100000010100000000000;
														assign node1276 = (inp[5]) ? 40'b0000001000001000000000000011100000000000 : 40'b0000001000001000000000000010100000000000;
													assign node1279 = (inp[6]) ? node1283 : node1280;
														assign node1280 = (inp[5]) ? 40'b1000001000000000000100000010000000000000 : 40'b1000001000000000000000000000000000000000;
														assign node1283 = (inp[12]) ? 40'b0000001000001000000000000011000000000000 : 40'b0000001000000000000100000010000000000000;

endmodule