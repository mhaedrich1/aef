module dtc_split5_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node25;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node33;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node39;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node57;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node67;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node81;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node95;
	wire [1-1:0] node97;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node103;
	wire [1-1:0] node105;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node121;
	wire [1-1:0] node123;
	wire [1-1:0] node125;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node131;
	wire [1-1:0] node134;
	wire [1-1:0] node135;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node143;
	wire [1-1:0] node146;
	wire [1-1:0] node147;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node158;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node167;
	wire [1-1:0] node170;
	wire [1-1:0] node171;
	wire [1-1:0] node173;
	wire [1-1:0] node175;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node181;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node193;
	wire [1-1:0] node195;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node203;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node226;
	wire [1-1:0] node227;
	wire [1-1:0] node229;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node241;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node249;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node261;
	wire [1-1:0] node263;
	wire [1-1:0] node265;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node271;
	wire [1-1:0] node273;
	wire [1-1:0] node276;
	wire [1-1:0] node277;
	wire [1-1:0] node279;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node295;
	wire [1-1:0] node297;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node317;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node324;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node329;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node335;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node343;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node347;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node361;
	wire [1-1:0] node364;
	wire [1-1:0] node365;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node371;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node383;
	wire [1-1:0] node385;
	wire [1-1:0] node387;
	wire [1-1:0] node389;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node395;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node401;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node411;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node417;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node427;
	wire [1-1:0] node429;
	wire [1-1:0] node431;
	wire [1-1:0] node433;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node439;
	wire [1-1:0] node441;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node447;
	wire [1-1:0] node450;
	wire [1-1:0] node451;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node459;
	wire [1-1:0] node461;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node467;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node475;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node487;
	wire [1-1:0] node488;
	wire [1-1:0] node489;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node501;
	wire [1-1:0] node504;
	wire [1-1:0] node505;
	wire [1-1:0] node507;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node515;
	wire [1-1:0] node516;
	wire [1-1:0] node517;
	wire [1-1:0] node519;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node525;
	wire [1-1:0] node528;
	wire [1-1:0] node529;
	wire [1-1:0] node533;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node557;
	wire [1-1:0] node559;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node565;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node573;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node577;
	wire [1-1:0] node580;
	wire [1-1:0] node581;
	wire [1-1:0] node585;
	wire [1-1:0] node586;
	wire [1-1:0] node587;
	wire [1-1:0] node592;
	wire [1-1:0] node593;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node597;
	wire [1-1:0] node600;
	wire [1-1:0] node601;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node607;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node627;
	wire [1-1:0] node629;
	wire [1-1:0] node631;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node637;
	wire [1-1:0] node639;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node645;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node662;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node671;
	wire [1-1:0] node673;
	wire [1-1:0] node676;
	wire [1-1:0] node677;
	wire [1-1:0] node681;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node691;
	wire [1-1:0] node693;
	wire [1-1:0] node695;
	wire [1-1:0] node698;
	wire [1-1:0] node699;
	wire [1-1:0] node701;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node713;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node722;
	wire [1-1:0] node723;
	wire [1-1:0] node724;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node731;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node741;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node751;
	wire [1-1:0] node753;
	wire [1-1:0] node755;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node761;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node769;
	wire [1-1:0] node770;
	wire [1-1:0] node771;
	wire [1-1:0] node773;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node781;
	wire [1-1:0] node782;
	wire [1-1:0] node783;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node793;
	wire [1-1:0] node796;
	wire [1-1:0] node797;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node804;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node828;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node844;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node855;
	wire [1-1:0] node857;
	wire [1-1:0] node860;
	wire [1-1:0] node861;
	wire [1-1:0] node863;
	wire [1-1:0] node865;
	wire [1-1:0] node867;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node877;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node893;
	wire [1-1:0] node895;
	wire [1-1:0] node897;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node903;
	wire [1-1:0] node905;
	wire [1-1:0] node908;
	wire [1-1:0] node909;
	wire [1-1:0] node911;
	wire [1-1:0] node914;
	wire [1-1:0] node915;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node923;
	wire [1-1:0] node924;
	wire [1-1:0] node928;
	wire [1-1:0] node929;
	wire [1-1:0] node931;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node939;
	wire [1-1:0] node940;
	wire [1-1:0] node941;
	wire [1-1:0] node943;
	wire [1-1:0] node946;
	wire [1-1:0] node947;
	wire [1-1:0] node951;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node958;
	wire [1-1:0] node959;
	wire [1-1:0] node960;
	wire [1-1:0] node961;
	wire [1-1:0] node963;
	wire [1-1:0] node965;
	wire [1-1:0] node967;
	wire [1-1:0] node970;
	wire [1-1:0] node971;
	wire [1-1:0] node973;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node979;
	wire [1-1:0] node982;
	wire [1-1:0] node983;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node993;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node999;
	wire [1-1:0] node1002;
	wire [1-1:0] node1003;
	wire [1-1:0] node1007;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1014;
	wire [1-1:0] node1015;
	wire [1-1:0] node1019;
	wire [1-1:0] node1020;
	wire [1-1:0] node1021;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1028;
	wire [1-1:0] node1029;
	wire [1-1:0] node1031;
	wire [1-1:0] node1033;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1039;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1047;
	wire [1-1:0] node1048;
	wire [1-1:0] node1049;
	wire [1-1:0] node1051;
	wire [1-1:0] node1054;
	wire [1-1:0] node1056;
	wire [1-1:0] node1059;
	wire [1-1:0] node1060;
	wire [1-1:0] node1061;
	wire [1-1:0] node1066;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1071;
	wire [1-1:0] node1074;
	wire [1-1:0] node1075;
	wire [1-1:0] node1080;
	wire [1-1:0] node1081;
	wire [1-1:0] node1082;
	wire [1-1:0] node1083;
	wire [1-1:0] node1089;
	wire [1-1:0] node1090;
	wire [1-1:0] node1091;
	wire [1-1:0] node1092;
	wire [1-1:0] node1094;
	wire [1-1:0] node1095;
	wire [1-1:0] node1097;
	wire [1-1:0] node1099;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1105;
	wire [1-1:0] node1108;
	wire [1-1:0] node1109;
	wire [1-1:0] node1113;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1117;
	wire [1-1:0] node1119;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1125;
	wire [1-1:0] node1128;
	wire [1-1:0] node1129;
	wire [1-1:0] node1133;
	wire [1-1:0] node1134;
	wire [1-1:0] node1135;
	wire [1-1:0] node1137;
	wire [1-1:0] node1140;
	wire [1-1:0] node1141;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1151;
	wire [1-1:0] node1153;
	wire [1-1:0] node1156;
	wire [1-1:0] node1157;
	wire [1-1:0] node1159;
	wire [1-1:0] node1162;
	wire [1-1:0] node1163;
	wire [1-1:0] node1167;
	wire [1-1:0] node1168;
	wire [1-1:0] node1169;
	wire [1-1:0] node1171;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1180;
	wire [1-1:0] node1181;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1185;
	wire [1-1:0] node1188;
	wire [1-1:0] node1189;
	wire [1-1:0] node1193;
	wire [1-1:0] node1194;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1200;
	wire [1-1:0] node1201;
	wire [1-1:0] node1207;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1210;
	wire [1-1:0] node1211;
	wire [1-1:0] node1213;
	wire [1-1:0] node1215;
	wire [1-1:0] node1218;
	wire [1-1:0] node1219;
	wire [1-1:0] node1221;
	wire [1-1:0] node1224;
	wire [1-1:0] node1225;
	wire [1-1:0] node1229;
	wire [1-1:0] node1230;
	wire [1-1:0] node1231;
	wire [1-1:0] node1233;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1240;
	wire [1-1:0] node1243;
	wire [1-1:0] node1244;
	wire [1-1:0] node1245;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1252;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1262;
	wire [1-1:0] node1263;
	wire [1-1:0] node1269;
	wire [1-1:0] node1270;
	wire [1-1:0] node1271;
	wire [1-1:0] node1272;
	wire [1-1:0] node1273;
	wire [1-1:0] node1275;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1290;
	wire [1-1:0] node1291;
	wire [1-1:0] node1292;
	wire [1-1:0] node1293;
	wire [1-1:0] node1299;
	wire [1-1:0] node1300;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1308;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1311;
	wire [1-1:0] node1312;
	wire [1-1:0] node1313;
	wire [1-1:0] node1315;
	wire [1-1:0] node1317;
	wire [1-1:0] node1319;
	wire [1-1:0] node1322;
	wire [1-1:0] node1323;
	wire [1-1:0] node1325;
	wire [1-1:0] node1327;
	wire [1-1:0] node1330;
	wire [1-1:0] node1331;
	wire [1-1:0] node1333;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1341;
	wire [1-1:0] node1342;
	wire [1-1:0] node1343;
	wire [1-1:0] node1345;
	wire [1-1:0] node1347;
	wire [1-1:0] node1350;
	wire [1-1:0] node1351;
	wire [1-1:0] node1353;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1361;
	wire [1-1:0] node1362;
	wire [1-1:0] node1363;
	wire [1-1:0] node1365;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1373;
	wire [1-1:0] node1374;
	wire [1-1:0] node1375;
	wire [1-1:0] node1380;
	wire [1-1:0] node1381;
	wire [1-1:0] node1382;
	wire [1-1:0] node1383;
	wire [1-1:0] node1385;
	wire [1-1:0] node1387;
	wire [1-1:0] node1390;
	wire [1-1:0] node1391;
	wire [1-1:0] node1393;
	wire [1-1:0] node1396;
	wire [1-1:0] node1397;
	wire [1-1:0] node1401;
	wire [1-1:0] node1402;
	wire [1-1:0] node1403;
	wire [1-1:0] node1405;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1413;
	wire [1-1:0] node1414;
	wire [1-1:0] node1415;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1425;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1438;
	wire [1-1:0] node1439;
	wire [1-1:0] node1440;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1449;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1452;
	wire [1-1:0] node1453;
	wire [1-1:0] node1455;
	wire [1-1:0] node1457;
	wire [1-1:0] node1460;
	wire [1-1:0] node1461;
	wire [1-1:0] node1463;
	wire [1-1:0] node1466;
	wire [1-1:0] node1467;
	wire [1-1:0] node1471;
	wire [1-1:0] node1472;
	wire [1-1:0] node1473;
	wire [1-1:0] node1475;
	wire [1-1:0] node1480;
	wire [1-1:0] node1481;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1485;
	wire [1-1:0] node1488;
	wire [1-1:0] node1489;
	wire [1-1:0] node1494;
	wire [1-1:0] node1495;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1505;
	wire [1-1:0] node1506;
	wire [1-1:0] node1507;
	wire [1-1:0] node1509;
	wire [1-1:0] node1512;
	wire [1-1:0] node1513;
	wire [1-1:0] node1517;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1522;
	wire [1-1:0] node1526;
	wire [1-1:0] node1527;
	wire [1-1:0] node1528;
	wire [1-1:0] node1529;
	wire [1-1:0] node1532;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1541;
	wire [1-1:0] node1548;
	wire [1-1:0] node1549;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1555;
	wire [1-1:0] node1557;
	wire [1-1:0] node1560;
	wire [1-1:0] node1561;
	wire [1-1:0] node1563;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1571;
	wire [1-1:0] node1572;
	wire [1-1:0] node1573;
	wire [1-1:0] node1575;
	wire [1-1:0] node1578;
	wire [1-1:0] node1579;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1590;
	wire [1-1:0] node1591;
	wire [1-1:0] node1592;
	wire [1-1:0] node1594;
	wire [1-1:0] node1595;
	wire [1-1:0] node1599;
	wire [1-1:0] node1600;
	wire [1-1:0] node1604;
	wire [1-1:0] node1605;
	wire [1-1:0] node1606;
	wire [1-1:0] node1607;
	wire [1-1:0] node1613;
	wire [1-1:0] node1614;
	wire [1-1:0] node1615;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1619;
	wire [1-1:0] node1622;
	wire [1-1:0] node1623;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1629;
	wire [1-1:0] node1634;
	wire [1-1:0] node1635;
	wire [1-1:0] node1636;
	wire [1-1:0] node1637;
	wire [1-1:0] node1643;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1654;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1657;
	wire [1-1:0] node1658;
	wire [1-1:0] node1659;
	wire [1-1:0] node1661;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1676;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1679;
	wire [1-1:0] node1685;
	wire [1-1:0] node1687;
	wire [1-1:0] node1688;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1696;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1699;
	wire [1-1:0] node1700;
	wire [1-1:0] node1701;

	assign outp = (inp[4]) ? node844 : node1;
		assign node1 = (inp[10]) ? node377 : node2;
			assign node2 = (inp[5]) ? node156 : node3;
				assign node3 = (inp[0]) ? node47 : node4;
					assign node4 = (inp[12]) ? node6 : 1'b1;
						assign node6 = (inp[2]) ? node18 : node7;
							assign node7 = (inp[3]) ? node9 : 1'b1;
								assign node9 = (inp[6]) ? node11 : 1'b1;
									assign node11 = (inp[7]) ? node13 : 1'b1;
										assign node13 = (inp[11]) ? node15 : 1'b1;
											assign node15 = (inp[8]) ? 1'b0 : 1'b1;
							assign node18 = (inp[1]) ? node28 : node19;
								assign node19 = (inp[3]) ? node21 : 1'b1;
									assign node21 = (inp[8]) ? node23 : 1'b1;
										assign node23 = (inp[9]) ? node25 : 1'b1;
											assign node25 = (inp[7]) ? 1'b0 : 1'b1;
								assign node28 = (inp[6]) ? node36 : node29;
									assign node29 = (inp[7]) ? node31 : 1'b1;
										assign node31 = (inp[3]) ? node33 : 1'b1;
											assign node33 = (inp[9]) ? 1'b0 : 1'b1;
									assign node36 = (inp[8]) ? node42 : node37;
										assign node37 = (inp[11]) ? node39 : 1'b1;
											assign node39 = (inp[9]) ? 1'b0 : 1'b1;
										assign node42 = (inp[3]) ? 1'b0 : node43;
											assign node43 = (inp[9]) ? 1'b0 : 1'b1;
					assign node47 = (inp[1]) ? node89 : node48;
						assign node48 = (inp[2]) ? node60 : node49;
							assign node49 = (inp[3]) ? node51 : 1'b1;
								assign node51 = (inp[7]) ? node53 : 1'b1;
									assign node53 = (inp[12]) ? node55 : 1'b1;
										assign node55 = (inp[9]) ? node57 : 1'b1;
											assign node57 = (inp[6]) ? 1'b0 : 1'b1;
							assign node60 = (inp[6]) ? node70 : node61;
								assign node61 = (inp[12]) ? node63 : 1'b1;
									assign node63 = (inp[7]) ? node65 : 1'b1;
										assign node65 = (inp[3]) ? node67 : 1'b1;
											assign node67 = (inp[9]) ? 1'b0 : 1'b1;
								assign node70 = (inp[3]) ? node78 : node71;
									assign node71 = (inp[8]) ? node73 : 1'b1;
										assign node73 = (inp[9]) ? node75 : 1'b1;
											assign node75 = (inp[7]) ? 1'b0 : 1'b1;
									assign node78 = (inp[12]) ? node84 : node79;
										assign node79 = (inp[11]) ? node81 : 1'b1;
											assign node81 = (inp[8]) ? 1'b1 : 1'b0;
										assign node84 = (inp[9]) ? 1'b0 : node85;
											assign node85 = (inp[8]) ? 1'b0 : 1'b1;
						assign node89 = (inp[8]) ? node119 : node90;
							assign node90 = (inp[11]) ? node100 : node91;
								assign node91 = (inp[12]) ? node93 : 1'b1;
									assign node93 = (inp[6]) ? node95 : 1'b1;
										assign node95 = (inp[7]) ? node97 : 1'b1;
											assign node97 = (inp[9]) ? 1'b0 : 1'b1;
								assign node100 = (inp[9]) ? node108 : node101;
									assign node101 = (inp[3]) ? node103 : 1'b1;
										assign node103 = (inp[6]) ? node105 : 1'b1;
											assign node105 = (inp[2]) ? 1'b0 : 1'b0;
									assign node108 = (inp[3]) ? node114 : node109;
										assign node109 = (inp[6]) ? 1'b0 : node110;
											assign node110 = (inp[12]) ? 1'b1 : 1'b1;
										assign node114 = (inp[2]) ? 1'b0 : node115;
											assign node115 = (inp[6]) ? 1'b0 : 1'b1;
							assign node119 = (inp[12]) ? node139 : node120;
								assign node120 = (inp[6]) ? node128 : node121;
									assign node121 = (inp[2]) ? node123 : 1'b1;
										assign node123 = (inp[9]) ? node125 : 1'b1;
											assign node125 = (inp[3]) ? 1'b0 : 1'b1;
									assign node128 = (inp[7]) ? node134 : node129;
										assign node129 = (inp[3]) ? node131 : 1'b1;
											assign node131 = (inp[11]) ? 1'b0 : 1'b1;
										assign node134 = (inp[11]) ? 1'b0 : node135;
											assign node135 = (inp[3]) ? 1'b0 : 1'b1;
								assign node139 = (inp[3]) ? node151 : node140;
									assign node140 = (inp[9]) ? node146 : node141;
										assign node141 = (inp[2]) ? node143 : 1'b1;
											assign node143 = (inp[6]) ? 1'b0 : 1'b1;
										assign node146 = (inp[6]) ? 1'b0 : node147;
											assign node147 = (inp[7]) ? 1'b0 : 1'b1;
									assign node151 = (inp[11]) ? 1'b0 : node152;
										assign node152 = (inp[6]) ? 1'b0 : 1'b1;
				assign node156 = (inp[6]) ? node256 : node157;
					assign node157 = (inp[2]) ? node189 : node158;
						assign node158 = (inp[3]) ? node160 : 1'b1;
							assign node160 = (inp[11]) ? node170 : node161;
								assign node161 = (inp[8]) ? node163 : 1'b1;
									assign node163 = (inp[0]) ? node165 : 1'b1;
										assign node165 = (inp[12]) ? node167 : 1'b1;
											assign node167 = (inp[7]) ? 1'b0 : 1'b1;
								assign node170 = (inp[1]) ? node178 : node171;
									assign node171 = (inp[9]) ? node173 : 1'b1;
										assign node173 = (inp[7]) ? node175 : 1'b1;
											assign node175 = (inp[12]) ? 1'b0 : 1'b1;
									assign node178 = (inp[7]) ? node184 : node179;
										assign node179 = (inp[0]) ? node181 : 1'b1;
											assign node181 = (inp[8]) ? 1'b0 : 1'b1;
										assign node184 = (inp[0]) ? 1'b0 : node185;
											assign node185 = (inp[12]) ? 1'b0 : 1'b1;
						assign node189 = (inp[9]) ? node217 : node190;
							assign node190 = (inp[7]) ? node198 : node191;
								assign node191 = (inp[8]) ? node193 : 1'b1;
									assign node193 = (inp[0]) ? node195 : 1'b1;
										assign node195 = (inp[1]) ? 1'b0 : 1'b1;
								assign node198 = (inp[12]) ? node206 : node199;
									assign node199 = (inp[11]) ? node201 : 1'b1;
										assign node201 = (inp[3]) ? node203 : 1'b1;
											assign node203 = (inp[8]) ? 1'b0 : 1'b1;
									assign node206 = (inp[8]) ? node212 : node207;
										assign node207 = (inp[0]) ? node209 : 1'b1;
											assign node209 = (inp[11]) ? 1'b0 : 1'b1;
										assign node212 = (inp[3]) ? 1'b0 : node213;
											assign node213 = (inp[11]) ? 1'b0 : 1'b1;
							assign node217 = (inp[8]) ? node237 : node218;
								assign node218 = (inp[12]) ? node226 : node219;
									assign node219 = (inp[1]) ? node221 : 1'b1;
										assign node221 = (inp[7]) ? node223 : 1'b1;
											assign node223 = (inp[0]) ? 1'b0 : 1'b1;
									assign node226 = (inp[0]) ? node232 : node227;
										assign node227 = (inp[3]) ? node229 : 1'b1;
											assign node229 = (inp[11]) ? 1'b0 : 1'b1;
										assign node232 = (inp[11]) ? 1'b0 : node233;
											assign node233 = (inp[7]) ? 1'b0 : 1'b1;
								assign node237 = (inp[1]) ? node249 : node238;
									assign node238 = (inp[11]) ? node244 : node239;
										assign node239 = (inp[0]) ? node241 : 1'b1;
											assign node241 = (inp[7]) ? 1'b0 : 1'b1;
										assign node244 = (inp[7]) ? 1'b0 : node245;
											assign node245 = (inp[3]) ? 1'b0 : 1'b1;
									assign node249 = (inp[0]) ? 1'b0 : node250;
										assign node250 = (inp[7]) ? 1'b0 : node251;
											assign node251 = (inp[11]) ? 1'b0 : 1'b0;
					assign node256 = (inp[2]) ? node324 : node257;
						assign node257 = (inp[0]) ? node287 : node258;
							assign node258 = (inp[8]) ? node268 : node259;
								assign node259 = (inp[7]) ? node261 : 1'b1;
									assign node261 = (inp[12]) ? node263 : 1'b1;
										assign node263 = (inp[11]) ? node265 : 1'b1;
											assign node265 = (inp[3]) ? 1'b0 : 1'b1;
								assign node268 = (inp[3]) ? node276 : node269;
									assign node269 = (inp[12]) ? node271 : 1'b1;
										assign node271 = (inp[7]) ? node273 : 1'b1;
											assign node273 = (inp[1]) ? 1'b0 : 1'b1;
									assign node276 = (inp[7]) ? node282 : node277;
										assign node277 = (inp[1]) ? node279 : 1'b1;
											assign node279 = (inp[12]) ? 1'b0 : 1'b1;
										assign node282 = (inp[9]) ? 1'b0 : node283;
											assign node283 = (inp[12]) ? 1'b0 : 1'b1;
							assign node287 = (inp[9]) ? node305 : node288;
								assign node288 = (inp[11]) ? node294 : node289;
									assign node289 = (inp[3]) ? node291 : 1'b1;
										assign node291 = (inp[1]) ? 1'b0 : 1'b1;
									assign node294 = (inp[8]) ? node300 : node295;
										assign node295 = (inp[1]) ? node297 : 1'b1;
											assign node297 = (inp[3]) ? 1'b0 : 1'b1;
										assign node300 = (inp[12]) ? 1'b0 : node301;
											assign node301 = (inp[3]) ? 1'b0 : 1'b1;
								assign node305 = (inp[11]) ? node317 : node306;
									assign node306 = (inp[12]) ? node312 : node307;
										assign node307 = (inp[1]) ? node309 : 1'b1;
											assign node309 = (inp[8]) ? 1'b0 : 1'b1;
										assign node312 = (inp[1]) ? 1'b0 : node313;
											assign node313 = (inp[7]) ? 1'b0 : 1'b1;
									assign node317 = (inp[8]) ? 1'b0 : node318;
										assign node318 = (inp[7]) ? 1'b0 : node319;
											assign node319 = (inp[1]) ? 1'b0 : 1'b0;
						assign node324 = (inp[3]) ? node356 : node325;
							assign node325 = (inp[0]) ? node343 : node326;
								assign node326 = (inp[1]) ? node332 : node327;
									assign node327 = (inp[12]) ? node329 : 1'b1;
										assign node329 = (inp[7]) ? 1'b0 : 1'b1;
									assign node332 = (inp[7]) ? node338 : node333;
										assign node333 = (inp[12]) ? node335 : 1'b1;
											assign node335 = (inp[11]) ? 1'b0 : 1'b1;
										assign node338 = (inp[9]) ? 1'b0 : node339;
											assign node339 = (inp[8]) ? 1'b0 : 1'b1;
								assign node343 = (inp[9]) ? 1'b0 : node344;
									assign node344 = (inp[11]) ? node350 : node345;
										assign node345 = (inp[8]) ? node347 : 1'b1;
											assign node347 = (inp[7]) ? 1'b0 : 1'b1;
										assign node350 = (inp[12]) ? 1'b0 : node351;
											assign node351 = (inp[1]) ? 1'b0 : 1'b1;
							assign node356 = (inp[7]) ? 1'b0 : node357;
								assign node357 = (inp[0]) ? node369 : node358;
									assign node358 = (inp[8]) ? node364 : node359;
										assign node359 = (inp[1]) ? node361 : 1'b1;
											assign node361 = (inp[9]) ? 1'b0 : 1'b1;
										assign node364 = (inp[11]) ? 1'b0 : node365;
											assign node365 = (inp[12]) ? 1'b0 : 1'b0;
									assign node369 = (inp[1]) ? 1'b0 : node370;
										assign node370 = (inp[12]) ? 1'b0 : node371;
											assign node371 = (inp[9]) ? 1'b0 : 1'b1;
			assign node377 = (inp[3]) ? node621 : node378;
				assign node378 = (inp[0]) ? node494 : node379;
					assign node379 = (inp[8]) ? node425 : node380;
						assign node380 = (inp[7]) ? node392 : node381;
							assign node381 = (inp[11]) ? node383 : 1'b1;
								assign node383 = (inp[1]) ? node385 : 1'b1;
									assign node385 = (inp[5]) ? node387 : 1'b1;
										assign node387 = (inp[2]) ? node389 : 1'b1;
											assign node389 = (inp[6]) ? 1'b0 : 1'b1;
							assign node392 = (inp[9]) ? node404 : node393;
								assign node393 = (inp[2]) ? node395 : 1'b1;
									assign node395 = (inp[1]) ? node397 : 1'b1;
										assign node397 = (inp[11]) ? node401 : node398;
											assign node398 = (inp[5]) ? 1'b1 : 1'b1;
											assign node401 = (inp[12]) ? 1'b0 : 1'b1;
								assign node404 = (inp[12]) ? node414 : node405;
									assign node405 = (inp[5]) ? node407 : 1'b1;
										assign node407 = (inp[6]) ? node411 : node408;
											assign node408 = (inp[2]) ? 1'b1 : 1'b1;
											assign node411 = (inp[1]) ? 1'b0 : 1'b0;
									assign node414 = (inp[11]) ? node420 : node415;
										assign node415 = (inp[2]) ? node417 : 1'b1;
											assign node417 = (inp[1]) ? 1'b0 : 1'b1;
										assign node420 = (inp[1]) ? 1'b0 : node421;
											assign node421 = (inp[6]) ? 1'b0 : 1'b1;
						assign node425 = (inp[9]) ? node455 : node426;
							assign node426 = (inp[12]) ? node436 : node427;
								assign node427 = (inp[5]) ? node429 : 1'b1;
									assign node429 = (inp[1]) ? node431 : 1'b1;
										assign node431 = (inp[6]) ? node433 : 1'b1;
											assign node433 = (inp[2]) ? 1'b0 : 1'b1;
								assign node436 = (inp[2]) ? node444 : node437;
									assign node437 = (inp[11]) ? node439 : 1'b1;
										assign node439 = (inp[6]) ? node441 : 1'b1;
											assign node441 = (inp[1]) ? 1'b0 : 1'b1;
									assign node444 = (inp[6]) ? node450 : node445;
										assign node445 = (inp[11]) ? node447 : 1'b1;
											assign node447 = (inp[1]) ? 1'b0 : 1'b1;
										assign node450 = (inp[7]) ? 1'b0 : node451;
											assign node451 = (inp[1]) ? 1'b0 : 1'b1;
							assign node455 = (inp[6]) ? node475 : node456;
								assign node456 = (inp[5]) ? node464 : node457;
									assign node457 = (inp[11]) ? node459 : 1'b1;
										assign node459 = (inp[7]) ? node461 : 1'b1;
											assign node461 = (inp[2]) ? 1'b0 : 1'b1;
									assign node464 = (inp[1]) ? node470 : node465;
										assign node465 = (inp[2]) ? node467 : 1'b1;
											assign node467 = (inp[7]) ? 1'b0 : 1'b1;
										assign node470 = (inp[11]) ? 1'b0 : node471;
											assign node471 = (inp[7]) ? 1'b0 : 1'b1;
								assign node475 = (inp[1]) ? node487 : node476;
									assign node476 = (inp[2]) ? node482 : node477;
										assign node477 = (inp[11]) ? node479 : 1'b1;
											assign node479 = (inp[7]) ? 1'b0 : 1'b1;
										assign node482 = (inp[12]) ? 1'b0 : node483;
											assign node483 = (inp[7]) ? 1'b0 : 1'b1;
									assign node487 = (inp[12]) ? 1'b0 : node488;
										assign node488 = (inp[5]) ? 1'b0 : node489;
											assign node489 = (inp[7]) ? 1'b0 : 1'b1;
					assign node494 = (inp[6]) ? node552 : node495;
						assign node495 = (inp[5]) ? node515 : node496;
							assign node496 = (inp[11]) ? node498 : 1'b1;
								assign node498 = (inp[9]) ? node504 : node499;
									assign node499 = (inp[1]) ? node501 : 1'b1;
										assign node501 = (inp[12]) ? 1'b0 : 1'b1;
									assign node504 = (inp[7]) ? node510 : node505;
										assign node505 = (inp[2]) ? node507 : 1'b1;
											assign node507 = (inp[8]) ? 1'b0 : 1'b1;
										assign node510 = (inp[12]) ? 1'b0 : node511;
											assign node511 = (inp[8]) ? 1'b0 : 1'b1;
							assign node515 = (inp[2]) ? node533 : node516;
								assign node516 = (inp[12]) ? node522 : node517;
									assign node517 = (inp[7]) ? node519 : 1'b1;
										assign node519 = (inp[1]) ? 1'b0 : 1'b1;
									assign node522 = (inp[11]) ? node528 : node523;
										assign node523 = (inp[8]) ? node525 : 1'b1;
											assign node525 = (inp[7]) ? 1'b0 : 1'b1;
										assign node528 = (inp[9]) ? 1'b0 : node529;
											assign node529 = (inp[7]) ? 1'b0 : 1'b1;
								assign node533 = (inp[1]) ? node545 : node534;
									assign node534 = (inp[7]) ? node540 : node535;
										assign node535 = (inp[12]) ? node537 : 1'b1;
											assign node537 = (inp[11]) ? 1'b0 : 1'b1;
										assign node540 = (inp[9]) ? 1'b0 : node541;
											assign node541 = (inp[8]) ? 1'b0 : 1'b1;
									assign node545 = (inp[8]) ? 1'b0 : node546;
										assign node546 = (inp[9]) ? 1'b0 : node547;
											assign node547 = (inp[12]) ? 1'b0 : 1'b1;
						assign node552 = (inp[11]) ? node592 : node553;
							assign node553 = (inp[1]) ? node573 : node554;
								assign node554 = (inp[12]) ? node562 : node555;
									assign node555 = (inp[9]) ? node557 : 1'b1;
										assign node557 = (inp[2]) ? node559 : 1'b1;
											assign node559 = (inp[5]) ? 1'b0 : 1'b1;
									assign node562 = (inp[9]) ? node568 : node563;
										assign node563 = (inp[8]) ? node565 : 1'b1;
											assign node565 = (inp[7]) ? 1'b0 : 1'b1;
										assign node568 = (inp[2]) ? 1'b0 : node569;
											assign node569 = (inp[5]) ? 1'b0 : 1'b1;
								assign node573 = (inp[8]) ? node585 : node574;
									assign node574 = (inp[2]) ? node580 : node575;
										assign node575 = (inp[7]) ? node577 : 1'b1;
											assign node577 = (inp[12]) ? 1'b0 : 1'b1;
										assign node580 = (inp[9]) ? 1'b0 : node581;
											assign node581 = (inp[7]) ? 1'b0 : 1'b1;
									assign node585 = (inp[2]) ? 1'b0 : node586;
										assign node586 = (inp[12]) ? 1'b0 : node587;
											assign node587 = (inp[9]) ? 1'b0 : 1'b1;
							assign node592 = (inp[5]) ? node612 : node593;
								assign node593 = (inp[12]) ? node605 : node594;
									assign node594 = (inp[7]) ? node600 : node595;
										assign node595 = (inp[9]) ? node597 : 1'b1;
											assign node597 = (inp[8]) ? 1'b0 : 1'b1;
										assign node600 = (inp[2]) ? 1'b0 : node601;
											assign node601 = (inp[1]) ? 1'b0 : 1'b1;
									assign node605 = (inp[9]) ? 1'b0 : node606;
										assign node606 = (inp[8]) ? 1'b0 : node607;
											assign node607 = (inp[2]) ? 1'b0 : 1'b1;
								assign node612 = (inp[2]) ? 1'b0 : node613;
									assign node613 = (inp[9]) ? 1'b0 : node614;
										assign node614 = (inp[8]) ? 1'b0 : node615;
											assign node615 = (inp[7]) ? 1'b0 : 1'b1;
				assign node621 = (inp[11]) ? node747 : node622;
					assign node622 = (inp[5]) ? node688 : node623;
						assign node623 = (inp[2]) ? node653 : node624;
							assign node624 = (inp[6]) ? node634 : node625;
								assign node625 = (inp[1]) ? node627 : 1'b1;
									assign node627 = (inp[8]) ? node629 : 1'b1;
										assign node629 = (inp[9]) ? node631 : 1'b1;
											assign node631 = (inp[12]) ? 1'b0 : 1'b1;
								assign node634 = (inp[0]) ? node642 : node635;
									assign node635 = (inp[12]) ? node637 : 1'b1;
										assign node637 = (inp[1]) ? node639 : 1'b1;
											assign node639 = (inp[8]) ? 1'b0 : 1'b1;
									assign node642 = (inp[8]) ? node648 : node643;
										assign node643 = (inp[12]) ? node645 : 1'b1;
											assign node645 = (inp[9]) ? 1'b0 : 1'b1;
										assign node648 = (inp[7]) ? 1'b0 : node649;
											assign node649 = (inp[1]) ? 1'b0 : 1'b1;
							assign node653 = (inp[6]) ? node669 : node654;
								assign node654 = (inp[1]) ? node662 : node655;
									assign node655 = (inp[7]) ? node657 : 1'b1;
										assign node657 = (inp[0]) ? node659 : 1'b1;
											assign node659 = (inp[9]) ? 1'b0 : 1'b1;
									assign node662 = (inp[8]) ? 1'b0 : node663;
										assign node663 = (inp[7]) ? node665 : 1'b1;
											assign node665 = (inp[0]) ? 1'b0 : 1'b1;
								assign node669 = (inp[8]) ? node681 : node670;
									assign node670 = (inp[1]) ? node676 : node671;
										assign node671 = (inp[12]) ? node673 : 1'b1;
											assign node673 = (inp[7]) ? 1'b0 : 1'b1;
										assign node676 = (inp[9]) ? 1'b0 : node677;
											assign node677 = (inp[0]) ? 1'b0 : 1'b1;
									assign node681 = (inp[0]) ? 1'b0 : node682;
										assign node682 = (inp[1]) ? 1'b0 : node683;
											assign node683 = (inp[7]) ? 1'b0 : 1'b1;
						assign node688 = (inp[1]) ? node722 : node689;
							assign node689 = (inp[7]) ? node709 : node690;
								assign node690 = (inp[2]) ? node698 : node691;
									assign node691 = (inp[0]) ? node693 : 1'b1;
										assign node693 = (inp[6]) ? node695 : 1'b1;
											assign node695 = (inp[12]) ? 1'b0 : 1'b1;
									assign node698 = (inp[12]) ? node704 : node699;
										assign node699 = (inp[6]) ? node701 : 1'b1;
											assign node701 = (inp[9]) ? 1'b0 : 1'b1;
										assign node704 = (inp[9]) ? 1'b0 : node705;
											assign node705 = (inp[6]) ? 1'b0 : 1'b1;
								assign node709 = (inp[6]) ? 1'b0 : node710;
									assign node710 = (inp[9]) ? node716 : node711;
										assign node711 = (inp[2]) ? node713 : 1'b1;
											assign node713 = (inp[0]) ? 1'b0 : 1'b1;
										assign node716 = (inp[2]) ? 1'b0 : node717;
											assign node717 = (inp[12]) ? 1'b0 : 1'b1;
							assign node722 = (inp[2]) ? node738 : node723;
								assign node723 = (inp[0]) ? node731 : node724;
									assign node724 = (inp[6]) ? node726 : 1'b1;
										assign node726 = (inp[8]) ? 1'b0 : node727;
											assign node727 = (inp[12]) ? 1'b0 : 1'b1;
									assign node731 = (inp[12]) ? 1'b0 : node732;
										assign node732 = (inp[7]) ? 1'b0 : node733;
											assign node733 = (inp[8]) ? 1'b0 : 1'b1;
								assign node738 = (inp[9]) ? 1'b0 : node739;
									assign node739 = (inp[12]) ? 1'b0 : node740;
										assign node740 = (inp[7]) ? 1'b0 : node741;
											assign node741 = (inp[8]) ? 1'b0 : 1'b1;
					assign node747 = (inp[7]) ? node809 : node748;
						assign node748 = (inp[9]) ? node788 : node749;
							assign node749 = (inp[2]) ? node769 : node750;
								assign node750 = (inp[12]) ? node758 : node751;
									assign node751 = (inp[0]) ? node753 : 1'b1;
										assign node753 = (inp[1]) ? node755 : 1'b1;
											assign node755 = (inp[6]) ? 1'b0 : 1'b1;
									assign node758 = (inp[5]) ? node764 : node759;
										assign node759 = (inp[6]) ? node761 : 1'b1;
											assign node761 = (inp[8]) ? 1'b0 : 1'b1;
										assign node764 = (inp[8]) ? 1'b0 : node765;
											assign node765 = (inp[0]) ? 1'b0 : 1'b1;
								assign node769 = (inp[8]) ? node781 : node770;
									assign node770 = (inp[6]) ? node776 : node771;
										assign node771 = (inp[0]) ? node773 : 1'b1;
											assign node773 = (inp[1]) ? 1'b0 : 1'b1;
										assign node776 = (inp[1]) ? 1'b0 : node777;
											assign node777 = (inp[0]) ? 1'b0 : 1'b1;
									assign node781 = (inp[12]) ? 1'b0 : node782;
										assign node782 = (inp[1]) ? 1'b0 : node783;
											assign node783 = (inp[0]) ? 1'b0 : 1'b1;
							assign node788 = (inp[8]) ? node802 : node789;
								assign node789 = (inp[1]) ? 1'b0 : node790;
									assign node790 = (inp[2]) ? node796 : node791;
										assign node791 = (inp[6]) ? node793 : 1'b1;
											assign node793 = (inp[12]) ? 1'b0 : 1'b1;
										assign node796 = (inp[5]) ? 1'b0 : node797;
											assign node797 = (inp[6]) ? 1'b0 : 1'b1;
								assign node802 = (inp[5]) ? 1'b0 : node803;
									assign node803 = (inp[6]) ? 1'b0 : node804;
										assign node804 = (inp[12]) ? 1'b0 : 1'b1;
						assign node809 = (inp[2]) ? node833 : node810;
							assign node810 = (inp[8]) ? node826 : node811;
								assign node811 = (inp[12]) ? node819 : node812;
									assign node812 = (inp[6]) ? node814 : 1'b1;
										assign node814 = (inp[0]) ? 1'b0 : node815;
											assign node815 = (inp[1]) ? 1'b0 : 1'b1;
									assign node819 = (inp[1]) ? 1'b0 : node820;
										assign node820 = (inp[0]) ? 1'b0 : node821;
											assign node821 = (inp[6]) ? 1'b0 : 1'b1;
								assign node826 = (inp[9]) ? 1'b0 : node827;
									assign node827 = (inp[5]) ? 1'b0 : node828;
										assign node828 = (inp[0]) ? 1'b0 : 1'b1;
							assign node833 = (inp[6]) ? 1'b0 : node834;
								assign node834 = (inp[1]) ? 1'b0 : node835;
									assign node835 = (inp[0]) ? 1'b0 : node836;
										assign node836 = (inp[12]) ? 1'b0 : node837;
											assign node837 = (inp[5]) ? 1'b0 : 1'b0;
		assign node844 = (inp[8]) ? node1308 : node845;
			assign node845 = (inp[0]) ? node1089 : node846;
				assign node846 = (inp[1]) ? node958 : node847;
					assign node847 = (inp[5]) ? node889 : node848;
						assign node848 = (inp[9]) ? node860 : node849;
							assign node849 = (inp[11]) ? node851 : 1'b1;
								assign node851 = (inp[10]) ? node853 : 1'b1;
									assign node853 = (inp[12]) ? node855 : 1'b1;
										assign node855 = (inp[2]) ? node857 : 1'b1;
											assign node857 = (inp[6]) ? 1'b0 : 1'b1;
							assign node860 = (inp[12]) ? node870 : node861;
								assign node861 = (inp[10]) ? node863 : 1'b1;
									assign node863 = (inp[7]) ? node865 : 1'b1;
										assign node865 = (inp[2]) ? node867 : 1'b1;
											assign node867 = (inp[11]) ? 1'b0 : 1'b1;
								assign node870 = (inp[11]) ? node880 : node871;
									assign node871 = (inp[6]) ? node873 : 1'b1;
										assign node873 = (inp[3]) ? node877 : node874;
											assign node874 = (inp[2]) ? 1'b1 : 1'b1;
											assign node877 = (inp[2]) ? 1'b0 : 1'b0;
									assign node880 = (inp[7]) ? node884 : node881;
										assign node881 = (inp[3]) ? 1'b0 : 1'b1;
										assign node884 = (inp[2]) ? 1'b0 : node885;
											assign node885 = (inp[6]) ? 1'b0 : 1'b1;
						assign node889 = (inp[6]) ? node919 : node890;
							assign node890 = (inp[12]) ? node900 : node891;
								assign node891 = (inp[2]) ? node893 : 1'b1;
									assign node893 = (inp[11]) ? node895 : 1'b1;
										assign node895 = (inp[7]) ? node897 : 1'b1;
											assign node897 = (inp[3]) ? 1'b0 : 1'b1;
								assign node900 = (inp[9]) ? node908 : node901;
									assign node901 = (inp[11]) ? node903 : 1'b1;
										assign node903 = (inp[7]) ? node905 : 1'b1;
											assign node905 = (inp[10]) ? 1'b0 : 1'b1;
									assign node908 = (inp[10]) ? node914 : node909;
										assign node909 = (inp[11]) ? node911 : 1'b1;
											assign node911 = (inp[3]) ? 1'b0 : 1'b1;
										assign node914 = (inp[7]) ? 1'b0 : node915;
											assign node915 = (inp[2]) ? 1'b0 : 1'b1;
							assign node919 = (inp[10]) ? node939 : node920;
								assign node920 = (inp[11]) ? node928 : node921;
									assign node921 = (inp[3]) ? node923 : 1'b1;
										assign node923 = (inp[7]) ? 1'b1 : node924;
											assign node924 = (inp[2]) ? 1'b0 : 1'b1;
									assign node928 = (inp[2]) ? node934 : node929;
										assign node929 = (inp[7]) ? node931 : 1'b1;
											assign node931 = (inp[9]) ? 1'b0 : 1'b1;
										assign node934 = (inp[7]) ? 1'b0 : node935;
											assign node935 = (inp[3]) ? 1'b0 : 1'b1;
								assign node939 = (inp[12]) ? node951 : node940;
									assign node940 = (inp[7]) ? node946 : node941;
										assign node941 = (inp[3]) ? node943 : 1'b1;
											assign node943 = (inp[11]) ? 1'b0 : 1'b1;
										assign node946 = (inp[9]) ? 1'b0 : node947;
											assign node947 = (inp[3]) ? 1'b0 : 1'b1;
									assign node951 = (inp[11]) ? 1'b0 : node952;
										assign node952 = (inp[2]) ? 1'b0 : node953;
											assign node953 = (inp[7]) ? 1'b0 : 1'b1;
					assign node958 = (inp[2]) ? node1026 : node959;
						assign node959 = (inp[9]) ? node987 : node960;
							assign node960 = (inp[11]) ? node970 : node961;
								assign node961 = (inp[6]) ? node963 : 1'b1;
									assign node963 = (inp[7]) ? node965 : 1'b1;
										assign node965 = (inp[12]) ? node967 : 1'b1;
											assign node967 = (inp[10]) ? 1'b0 : 1'b1;
								assign node970 = (inp[3]) ? node976 : node971;
									assign node971 = (inp[7]) ? node973 : 1'b1;
										assign node973 = (inp[5]) ? 1'b0 : 1'b1;
									assign node976 = (inp[12]) ? node982 : node977;
										assign node977 = (inp[10]) ? node979 : 1'b1;
											assign node979 = (inp[6]) ? 1'b0 : 1'b1;
										assign node982 = (inp[10]) ? 1'b0 : node983;
											assign node983 = (inp[5]) ? 1'b0 : 1'b0;
							assign node987 = (inp[10]) ? node1007 : node988;
								assign node988 = (inp[7]) ? node996 : node989;
									assign node989 = (inp[5]) ? node991 : 1'b1;
										assign node991 = (inp[3]) ? node993 : 1'b1;
											assign node993 = (inp[12]) ? 1'b0 : 1'b1;
									assign node996 = (inp[12]) ? node1002 : node997;
										assign node997 = (inp[5]) ? node999 : 1'b1;
											assign node999 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1002 = (inp[3]) ? 1'b0 : node1003;
											assign node1003 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1007 = (inp[3]) ? node1019 : node1008;
									assign node1008 = (inp[5]) ? node1014 : node1009;
										assign node1009 = (inp[11]) ? node1011 : 1'b1;
											assign node1011 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1014 = (inp[12]) ? 1'b0 : node1015;
											assign node1015 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1019 = (inp[6]) ? 1'b0 : node1020;
										assign node1020 = (inp[7]) ? 1'b0 : node1021;
											assign node1021 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1026 = (inp[6]) ? node1066 : node1027;
							assign node1027 = (inp[5]) ? node1047 : node1028;
								assign node1028 = (inp[7]) ? node1036 : node1029;
									assign node1029 = (inp[9]) ? node1031 : 1'b1;
										assign node1031 = (inp[12]) ? node1033 : 1'b1;
											assign node1033 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1036 = (inp[12]) ? node1042 : node1037;
										assign node1037 = (inp[11]) ? node1039 : 1'b1;
											assign node1039 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1042 = (inp[9]) ? 1'b0 : node1043;
											assign node1043 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1047 = (inp[3]) ? node1059 : node1048;
									assign node1048 = (inp[12]) ? node1054 : node1049;
										assign node1049 = (inp[9]) ? node1051 : 1'b1;
											assign node1051 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1054 = (inp[10]) ? node1056 : 1'b0;
											assign node1056 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1059 = (inp[9]) ? 1'b0 : node1060;
										assign node1060 = (inp[11]) ? 1'b0 : node1061;
											assign node1061 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1066 = (inp[7]) ? node1080 : node1067;
								assign node1067 = (inp[5]) ? 1'b0 : node1068;
									assign node1068 = (inp[12]) ? node1074 : node1069;
										assign node1069 = (inp[10]) ? node1071 : 1'b1;
											assign node1071 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1074 = (inp[10]) ? 1'b0 : node1075;
											assign node1075 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1080 = (inp[10]) ? 1'b0 : node1081;
									assign node1081 = (inp[11]) ? 1'b0 : node1082;
										assign node1082 = (inp[5]) ? 1'b0 : node1083;
											assign node1083 = (inp[3]) ? 1'b0 : 1'b1;
				assign node1089 = (inp[7]) ? node1207 : node1090;
					assign node1090 = (inp[6]) ? node1146 : node1091;
						assign node1091 = (inp[11]) ? node1113 : node1092;
							assign node1092 = (inp[2]) ? node1094 : 1'b1;
								assign node1094 = (inp[9]) ? node1102 : node1095;
									assign node1095 = (inp[1]) ? node1097 : 1'b1;
										assign node1097 = (inp[10]) ? node1099 : 1'b1;
											assign node1099 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1102 = (inp[3]) ? node1108 : node1103;
										assign node1103 = (inp[10]) ? node1105 : 1'b1;
											assign node1105 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1108 = (inp[12]) ? 1'b0 : node1109;
											assign node1109 = (inp[5]) ? 1'b0 : 1'b1;
							assign node1113 = (inp[3]) ? node1133 : node1114;
								assign node1114 = (inp[12]) ? node1122 : node1115;
									assign node1115 = (inp[9]) ? node1117 : 1'b1;
										assign node1117 = (inp[1]) ? node1119 : 1'b1;
											assign node1119 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1122 = (inp[10]) ? node1128 : node1123;
										assign node1123 = (inp[5]) ? node1125 : 1'b1;
											assign node1125 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1128 = (inp[2]) ? 1'b0 : node1129;
											assign node1129 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1133 = (inp[5]) ? 1'b0 : node1134;
									assign node1134 = (inp[9]) ? node1140 : node1135;
										assign node1135 = (inp[1]) ? node1137 : 1'b1;
											assign node1137 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1140 = (inp[1]) ? 1'b0 : node1141;
											assign node1141 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1146 = (inp[9]) ? node1180 : node1147;
							assign node1147 = (inp[10]) ? node1167 : node1148;
								assign node1148 = (inp[2]) ? node1156 : node1149;
									assign node1149 = (inp[3]) ? node1151 : 1'b1;
										assign node1151 = (inp[1]) ? node1153 : 1'b1;
											assign node1153 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1156 = (inp[11]) ? node1162 : node1157;
										assign node1157 = (inp[3]) ? node1159 : 1'b1;
											assign node1159 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1162 = (inp[12]) ? 1'b0 : node1163;
											assign node1163 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1167 = (inp[1]) ? 1'b0 : node1168;
									assign node1168 = (inp[5]) ? node1174 : node1169;
										assign node1169 = (inp[3]) ? node1171 : 1'b1;
											assign node1171 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1174 = (inp[2]) ? 1'b0 : node1175;
											assign node1175 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1180 = (inp[11]) ? node1198 : node1181;
								assign node1181 = (inp[1]) ? node1193 : node1182;
									assign node1182 = (inp[12]) ? node1188 : node1183;
										assign node1183 = (inp[2]) ? node1185 : 1'b1;
											assign node1185 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1188 = (inp[2]) ? 1'b0 : node1189;
											assign node1189 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1193 = (inp[10]) ? 1'b0 : node1194;
										assign node1194 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1198 = (inp[2]) ? 1'b0 : node1199;
									assign node1199 = (inp[12]) ? 1'b0 : node1200;
										assign node1200 = (inp[3]) ? 1'b0 : node1201;
											assign node1201 = (inp[5]) ? 1'b0 : 1'b1;
					assign node1207 = (inp[3]) ? node1269 : node1208;
						assign node1208 = (inp[1]) ? node1250 : node1209;
							assign node1209 = (inp[5]) ? node1229 : node1210;
								assign node1210 = (inp[10]) ? node1218 : node1211;
									assign node1211 = (inp[12]) ? node1213 : 1'b1;
										assign node1213 = (inp[2]) ? node1215 : 1'b1;
											assign node1215 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1218 = (inp[6]) ? node1224 : node1219;
										assign node1219 = (inp[9]) ? node1221 : 1'b1;
											assign node1221 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1224 = (inp[12]) ? 1'b0 : node1225;
											assign node1225 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1229 = (inp[9]) ? node1243 : node1230;
									assign node1230 = (inp[12]) ? node1236 : node1231;
										assign node1231 = (inp[6]) ? node1233 : 1'b1;
											assign node1233 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1236 = (inp[2]) ? node1240 : node1237;
											assign node1237 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1240 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1243 = (inp[6]) ? 1'b0 : node1244;
										assign node1244 = (inp[11]) ? 1'b0 : node1245;
											assign node1245 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1250 = (inp[12]) ? node1260 : node1251;
								assign node1251 = (inp[11]) ? 1'b0 : node1252;
									assign node1252 = (inp[6]) ? node1254 : 1'b1;
										assign node1254 = (inp[5]) ? 1'b0 : node1255;
											assign node1255 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1260 = (inp[2]) ? 1'b0 : node1261;
									assign node1261 = (inp[10]) ? 1'b0 : node1262;
										assign node1262 = (inp[6]) ? 1'b0 : node1263;
											assign node1263 = (inp[9]) ? 1'b0 : 1'b1;
						assign node1269 = (inp[5]) ? node1299 : node1270;
							assign node1270 = (inp[10]) ? node1290 : node1271;
								assign node1271 = (inp[12]) ? node1283 : node1272;
									assign node1272 = (inp[1]) ? node1278 : node1273;
										assign node1273 = (inp[2]) ? node1275 : 1'b1;
											assign node1275 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1278 = (inp[11]) ? 1'b0 : node1279;
											assign node1279 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1283 = (inp[6]) ? 1'b0 : node1284;
										assign node1284 = (inp[2]) ? 1'b0 : node1285;
											assign node1285 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1290 = (inp[6]) ? 1'b0 : node1291;
									assign node1291 = (inp[9]) ? 1'b0 : node1292;
										assign node1292 = (inp[2]) ? 1'b0 : node1293;
											assign node1293 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1299 = (inp[2]) ? 1'b0 : node1300;
								assign node1300 = (inp[12]) ? 1'b0 : node1301;
									assign node1301 = (inp[11]) ? 1'b0 : node1302;
										assign node1302 = (inp[1]) ? 1'b0 : 1'b1;
			assign node1308 = (inp[1]) ? node1548 : node1309;
				assign node1309 = (inp[11]) ? node1449 : node1310;
					assign node1310 = (inp[9]) ? node1380 : node1311;
						assign node1311 = (inp[5]) ? node1341 : node1312;
							assign node1312 = (inp[2]) ? node1322 : node1313;
								assign node1313 = (inp[6]) ? node1315 : 1'b1;
									assign node1315 = (inp[7]) ? node1317 : 1'b1;
										assign node1317 = (inp[12]) ? node1319 : 1'b1;
											assign node1319 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1322 = (inp[12]) ? node1330 : node1323;
									assign node1323 = (inp[0]) ? node1325 : 1'b1;
										assign node1325 = (inp[7]) ? node1327 : 1'b1;
											assign node1327 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1330 = (inp[3]) ? node1336 : node1331;
										assign node1331 = (inp[10]) ? node1333 : 1'b1;
											assign node1333 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1336 = (inp[6]) ? 1'b0 : node1337;
											assign node1337 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1341 = (inp[3]) ? node1361 : node1342;
								assign node1342 = (inp[2]) ? node1350 : node1343;
									assign node1343 = (inp[6]) ? node1345 : 1'b1;
										assign node1345 = (inp[10]) ? node1347 : 1'b1;
											assign node1347 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1350 = (inp[0]) ? node1356 : node1351;
										assign node1351 = (inp[6]) ? node1353 : 1'b1;
											assign node1353 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1356 = (inp[10]) ? 1'b0 : node1357;
											assign node1357 = (inp[12]) ? 1'b0 : 1'b1;
								assign node1361 = (inp[10]) ? node1373 : node1362;
									assign node1362 = (inp[7]) ? node1368 : node1363;
										assign node1363 = (inp[6]) ? node1365 : 1'b1;
											assign node1365 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1368 = (inp[12]) ? 1'b0 : node1369;
											assign node1369 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1373 = (inp[0]) ? 1'b0 : node1374;
										assign node1374 = (inp[7]) ? 1'b0 : node1375;
											assign node1375 = (inp[6]) ? 1'b0 : 1'b1;
						assign node1380 = (inp[3]) ? node1420 : node1381;
							assign node1381 = (inp[12]) ? node1401 : node1382;
								assign node1382 = (inp[5]) ? node1390 : node1383;
									assign node1383 = (inp[7]) ? node1385 : 1'b1;
										assign node1385 = (inp[2]) ? node1387 : 1'b1;
											assign node1387 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1390 = (inp[0]) ? node1396 : node1391;
										assign node1391 = (inp[2]) ? node1393 : 1'b1;
											assign node1393 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1396 = (inp[2]) ? 1'b0 : node1397;
											assign node1397 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1401 = (inp[7]) ? node1413 : node1402;
									assign node1402 = (inp[2]) ? node1408 : node1403;
										assign node1403 = (inp[10]) ? node1405 : 1'b1;
											assign node1405 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1408 = (inp[10]) ? 1'b0 : node1409;
											assign node1409 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1413 = (inp[6]) ? 1'b0 : node1414;
										assign node1414 = (inp[0]) ? 1'b0 : node1415;
											assign node1415 = (inp[2]) ? 1'b0 : 1'b1;
							assign node1420 = (inp[7]) ? node1438 : node1421;
								assign node1421 = (inp[6]) ? node1433 : node1422;
									assign node1422 = (inp[12]) ? node1428 : node1423;
										assign node1423 = (inp[10]) ? node1425 : 1'b1;
											assign node1425 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1428 = (inp[0]) ? 1'b0 : node1429;
											assign node1429 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1433 = (inp[12]) ? 1'b0 : node1434;
										assign node1434 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1438 = (inp[2]) ? 1'b0 : node1439;
									assign node1439 = (inp[10]) ? node1443 : node1440;
										assign node1440 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1443 = (inp[6]) ? 1'b0 : node1444;
											assign node1444 = (inp[0]) ? 1'b0 : 1'b0;
					assign node1449 = (inp[2]) ? node1503 : node1450;
						assign node1450 = (inp[9]) ? node1480 : node1451;
							assign node1451 = (inp[12]) ? node1471 : node1452;
								assign node1452 = (inp[3]) ? node1460 : node1453;
									assign node1453 = (inp[7]) ? node1455 : 1'b1;
										assign node1455 = (inp[10]) ? node1457 : 1'b1;
											assign node1457 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1460 = (inp[7]) ? node1466 : node1461;
										assign node1461 = (inp[5]) ? node1463 : 1'b1;
											assign node1463 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1466 = (inp[6]) ? 1'b0 : node1467;
											assign node1467 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1471 = (inp[6]) ? 1'b0 : node1472;
									assign node1472 = (inp[7]) ? 1'b0 : node1473;
										assign node1473 = (inp[10]) ? node1475 : 1'b1;
											assign node1475 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1480 = (inp[10]) ? node1494 : node1481;
								assign node1481 = (inp[0]) ? 1'b0 : node1482;
									assign node1482 = (inp[7]) ? node1488 : node1483;
										assign node1483 = (inp[5]) ? node1485 : 1'b1;
											assign node1485 = (inp[12]) ? 1'b0 : 1'b0;
										assign node1488 = (inp[3]) ? 1'b0 : node1489;
											assign node1489 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1494 = (inp[3]) ? 1'b0 : node1495;
									assign node1495 = (inp[5]) ? 1'b0 : node1496;
										assign node1496 = (inp[12]) ? 1'b0 : node1497;
											assign node1497 = (inp[6]) ? 1'b0 : 1'b1;
						assign node1503 = (inp[5]) ? node1537 : node1504;
							assign node1504 = (inp[10]) ? node1526 : node1505;
								assign node1505 = (inp[9]) ? node1517 : node1506;
									assign node1506 = (inp[6]) ? node1512 : node1507;
										assign node1507 = (inp[3]) ? node1509 : 1'b1;
											assign node1509 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1512 = (inp[0]) ? 1'b0 : node1513;
											assign node1513 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1517 = (inp[0]) ? 1'b0 : node1518;
										assign node1518 = (inp[7]) ? node1522 : node1519;
											assign node1519 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1522 = (inp[6]) ? 1'b0 : 1'b0;
								assign node1526 = (inp[9]) ? 1'b0 : node1527;
									assign node1527 = (inp[0]) ? 1'b0 : node1528;
										assign node1528 = (inp[12]) ? node1532 : node1529;
											assign node1529 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1532 = (inp[7]) ? 1'b0 : 1'b0;
							assign node1537 = (inp[10]) ? 1'b0 : node1538;
								assign node1538 = (inp[0]) ? 1'b0 : node1539;
									assign node1539 = (inp[7]) ? 1'b0 : node1540;
										assign node1540 = (inp[12]) ? 1'b0 : node1541;
											assign node1541 = (inp[9]) ? 1'b0 : 1'b0;
				assign node1548 = (inp[9]) ? node1654 : node1549;
					assign node1549 = (inp[2]) ? node1613 : node1550;
						assign node1550 = (inp[12]) ? node1590 : node1551;
							assign node1551 = (inp[7]) ? node1571 : node1552;
								assign node1552 = (inp[0]) ? node1560 : node1553;
									assign node1553 = (inp[6]) ? node1555 : 1'b1;
										assign node1555 = (inp[5]) ? node1557 : 1'b1;
											assign node1557 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1560 = (inp[10]) ? node1566 : node1561;
										assign node1561 = (inp[11]) ? node1563 : 1'b1;
											assign node1563 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1566 = (inp[11]) ? 1'b0 : node1567;
											assign node1567 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1571 = (inp[5]) ? node1583 : node1572;
									assign node1572 = (inp[6]) ? node1578 : node1573;
										assign node1573 = (inp[3]) ? node1575 : 1'b1;
											assign node1575 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1578 = (inp[0]) ? 1'b0 : node1579;
											assign node1579 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1583 = (inp[3]) ? 1'b0 : node1584;
										assign node1584 = (inp[10]) ? 1'b0 : node1585;
											assign node1585 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1590 = (inp[0]) ? node1604 : node1591;
								assign node1591 = (inp[10]) ? node1599 : node1592;
									assign node1592 = (inp[3]) ? node1594 : 1'b1;
										assign node1594 = (inp[11]) ? 1'b0 : node1595;
											assign node1595 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1599 = (inp[6]) ? 1'b0 : node1600;
										assign node1600 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1604 = (inp[7]) ? 1'b0 : node1605;
									assign node1605 = (inp[3]) ? 1'b0 : node1606;
										assign node1606 = (inp[11]) ? 1'b0 : node1607;
											assign node1607 = (inp[5]) ? 1'b0 : 1'b1;
						assign node1613 = (inp[0]) ? node1643 : node1614;
							assign node1614 = (inp[6]) ? node1634 : node1615;
								assign node1615 = (inp[3]) ? node1627 : node1616;
									assign node1616 = (inp[5]) ? node1622 : node1617;
										assign node1617 = (inp[11]) ? node1619 : 1'b1;
											assign node1619 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1622 = (inp[7]) ? 1'b0 : node1623;
											assign node1623 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1627 = (inp[11]) ? 1'b0 : node1628;
										assign node1628 = (inp[5]) ? 1'b0 : node1629;
											assign node1629 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1634 = (inp[11]) ? 1'b0 : node1635;
									assign node1635 = (inp[3]) ? 1'b0 : node1636;
										assign node1636 = (inp[7]) ? 1'b0 : node1637;
											assign node1637 = (inp[12]) ? 1'b0 : 1'b1;
							assign node1643 = (inp[7]) ? 1'b0 : node1644;
								assign node1644 = (inp[6]) ? 1'b0 : node1645;
									assign node1645 = (inp[3]) ? 1'b0 : node1646;
										assign node1646 = (inp[5]) ? 1'b0 : node1647;
											assign node1647 = (inp[10]) ? 1'b0 : 1'b0;
					assign node1654 = (inp[5]) ? node1696 : node1655;
						assign node1655 = (inp[3]) ? node1685 : node1656;
							assign node1656 = (inp[2]) ? node1676 : node1657;
								assign node1657 = (inp[7]) ? node1669 : node1658;
									assign node1658 = (inp[6]) ? node1664 : node1659;
										assign node1659 = (inp[10]) ? node1661 : 1'b1;
											assign node1661 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1664 = (inp[0]) ? 1'b0 : node1665;
											assign node1665 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1669 = (inp[11]) ? 1'b0 : node1670;
										assign node1670 = (inp[10]) ? 1'b0 : node1671;
											assign node1671 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1676 = (inp[12]) ? 1'b0 : node1677;
									assign node1677 = (inp[10]) ? 1'b0 : node1678;
										assign node1678 = (inp[11]) ? 1'b0 : node1679;
											assign node1679 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1685 = (inp[10]) ? node1687 : 1'b0;
								assign node1687 = (inp[12]) ? 1'b0 : node1688;
									assign node1688 = (inp[7]) ? 1'b0 : node1689;
										assign node1689 = (inp[2]) ? 1'b0 : node1690;
											assign node1690 = (inp[6]) ? 1'b0 : 1'b0;
						assign node1696 = (inp[12]) ? 1'b0 : node1697;
							assign node1697 = (inp[0]) ? 1'b0 : node1698;
								assign node1698 = (inp[6]) ? 1'b0 : node1699;
									assign node1699 = (inp[10]) ? 1'b0 : node1700;
										assign node1700 = (inp[7]) ? 1'b0 : node1701;
											assign node1701 = (inp[2]) ? 1'b0 : 1'b1;

endmodule