module dtc_split5_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node16;
	wire [4-1:0] node19;
	wire [4-1:0] node21;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node42;
	wire [4-1:0] node45;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node80;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node91;
	wire [4-1:0] node93;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node105;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node112;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node150;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node159;
	wire [4-1:0] node161;
	wire [4-1:0] node165;
	wire [4-1:0] node166;
	wire [4-1:0] node168;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node178;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node190;
	wire [4-1:0] node192;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node211;
	wire [4-1:0] node213;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node251;
	wire [4-1:0] node253;
	wire [4-1:0] node256;
	wire [4-1:0] node258;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node270;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node279;
	wire [4-1:0] node281;
	wire [4-1:0] node284;
	wire [4-1:0] node285;
	wire [4-1:0] node286;
	wire [4-1:0] node288;
	wire [4-1:0] node290;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node309;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node320;
	wire [4-1:0] node323;
	wire [4-1:0] node325;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node336;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node349;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node377;
	wire [4-1:0] node379;
	wire [4-1:0] node382;
	wire [4-1:0] node384;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node400;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node408;
	wire [4-1:0] node410;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node417;
	wire [4-1:0] node419;
	wire [4-1:0] node422;
	wire [4-1:0] node423;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node437;
	wire [4-1:0] node439;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node445;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node457;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node489;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node499;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node506;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node512;
	wire [4-1:0] node513;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node525;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node540;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node548;
	wire [4-1:0] node549;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node563;
	wire [4-1:0] node564;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node581;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node594;
	wire [4-1:0] node596;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node605;
	wire [4-1:0] node608;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node618;
	wire [4-1:0] node620;
	wire [4-1:0] node623;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node628;
	wire [4-1:0] node631;
	wire [4-1:0] node632;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node647;
	wire [4-1:0] node649;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node660;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node666;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node673;
	wire [4-1:0] node676;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node682;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node688;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node697;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node743;
	wire [4-1:0] node745;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node801;
	wire [4-1:0] node803;
	wire [4-1:0] node805;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node813;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node824;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node846;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node854;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node867;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node940;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node950;
	wire [4-1:0] node952;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node961;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node973;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node984;
	wire [4-1:0] node985;
	wire [4-1:0] node987;
	wire [4-1:0] node991;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1008;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1053;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1083;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1106;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1118;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1122;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1141;
	wire [4-1:0] node1143;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1167;
	wire [4-1:0] node1169;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1177;
	wire [4-1:0] node1179;
	wire [4-1:0] node1181;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1190;
	wire [4-1:0] node1194;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1206;
	wire [4-1:0] node1208;
	wire [4-1:0] node1211;
	wire [4-1:0] node1213;
	wire [4-1:0] node1214;
	wire [4-1:0] node1217;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1243;
	wire [4-1:0] node1244;
	wire [4-1:0] node1247;
	wire [4-1:0] node1249;
	wire [4-1:0] node1252;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1259;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1265;
	wire [4-1:0] node1268;
	wire [4-1:0] node1269;
	wire [4-1:0] node1271;
	wire [4-1:0] node1274;
	wire [4-1:0] node1276;
	wire [4-1:0] node1277;
	wire [4-1:0] node1280;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1301;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1313;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1331;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1350;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1361;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1369;
	wire [4-1:0] node1371;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1382;
	wire [4-1:0] node1385;
	wire [4-1:0] node1387;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1394;
	wire [4-1:0] node1396;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1418;
	wire [4-1:0] node1420;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1432;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1440;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1447;
	wire [4-1:0] node1451;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1457;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1485;
	wire [4-1:0] node1488;
	wire [4-1:0] node1489;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1500;
	wire [4-1:0] node1502;
	wire [4-1:0] node1505;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1521;
	wire [4-1:0] node1523;
	wire [4-1:0] node1525;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1534;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1544;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1550;
	wire [4-1:0] node1553;
	wire [4-1:0] node1554;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1560;
	wire [4-1:0] node1563;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1569;
	wire [4-1:0] node1572;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1584;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1591;
	wire [4-1:0] node1593;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1604;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1616;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1631;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1648;
	wire [4-1:0] node1652;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1657;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1671;
	wire [4-1:0] node1674;
	wire [4-1:0] node1675;
	wire [4-1:0] node1677;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1684;
	wire [4-1:0] node1687;
	wire [4-1:0] node1689;
	wire [4-1:0] node1692;
	wire [4-1:0] node1693;
	wire [4-1:0] node1696;
	wire [4-1:0] node1698;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1708;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1732;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1740;
	wire [4-1:0] node1742;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1760;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1775;
	wire [4-1:0] node1778;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1788;
	wire [4-1:0] node1789;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1806;
	wire [4-1:0] node1808;
	wire [4-1:0] node1810;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1825;
	wire [4-1:0] node1827;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1836;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1857;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1861;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1869;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1877;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1892;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1916;
	wire [4-1:0] node1919;
	wire [4-1:0] node1922;
	wire [4-1:0] node1924;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1936;
	wire [4-1:0] node1938;
	wire [4-1:0] node1943;
	wire [4-1:0] node1945;
	wire [4-1:0] node1947;
	wire [4-1:0] node1949;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1960;
	wire [4-1:0] node1962;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1968;
	wire [4-1:0] node1971;
	wire [4-1:0] node1973;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1987;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1994;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2003;
	wire [4-1:0] node2006;
	wire [4-1:0] node2008;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2018;
	wire [4-1:0] node2021;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2029;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2035;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2042;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2051;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2062;
	wire [4-1:0] node2066;
	wire [4-1:0] node2068;
	wire [4-1:0] node2070;
	wire [4-1:0] node2072;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2084;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2112;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2150;
	wire [4-1:0] node2154;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2167;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2179;
	wire [4-1:0] node2182;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2187;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2198;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2208;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2220;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2232;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2239;
	wire [4-1:0] node2242;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2255;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2264;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2275;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2281;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2294;
	wire [4-1:0] node2298;
	wire [4-1:0] node2300;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2306;
	wire [4-1:0] node2308;
	wire [4-1:0] node2311;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2318;
	wire [4-1:0] node2321;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2328;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2332;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2339;
	wire [4-1:0] node2343;
	wire [4-1:0] node2345;
	wire [4-1:0] node2346;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2353;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2358;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2365;
	wire [4-1:0] node2368;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2374;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2384;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2390;
	wire [4-1:0] node2393;
	wire [4-1:0] node2394;
	wire [4-1:0] node2395;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2402;
	wire [4-1:0] node2405;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2416;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2422;
	wire [4-1:0] node2424;
	wire [4-1:0] node2427;
	wire [4-1:0] node2428;
	wire [4-1:0] node2429;
	wire [4-1:0] node2431;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2438;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2443;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2453;
	wire [4-1:0] node2454;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2471;
	wire [4-1:0] node2472;
	wire [4-1:0] node2473;
	wire [4-1:0] node2474;
	wire [4-1:0] node2478;
	wire [4-1:0] node2480;
	wire [4-1:0] node2483;
	wire [4-1:0] node2485;
	wire [4-1:0] node2487;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2494;
	wire [4-1:0] node2496;
	wire [4-1:0] node2499;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2505;
	wire [4-1:0] node2508;
	wire [4-1:0] node2509;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2516;
	wire [4-1:0] node2517;
	wire [4-1:0] node2518;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2526;
	wire [4-1:0] node2528;
	wire [4-1:0] node2529;
	wire [4-1:0] node2533;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2561;
	wire [4-1:0] node2564;
	wire [4-1:0] node2565;
	wire [4-1:0] node2566;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2573;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2579;
	wire [4-1:0] node2582;
	wire [4-1:0] node2585;
	wire [4-1:0] node2586;
	wire [4-1:0] node2587;
	wire [4-1:0] node2590;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2598;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2604;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2613;
	wire [4-1:0] node2617;
	wire [4-1:0] node2619;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2627;
	wire [4-1:0] node2630;
	wire [4-1:0] node2631;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2637;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2644;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2657;
	wire [4-1:0] node2661;
	wire [4-1:0] node2663;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2669;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2682;
	wire [4-1:0] node2687;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2694;
	wire [4-1:0] node2697;
	wire [4-1:0] node2699;
	wire [4-1:0] node2702;
	wire [4-1:0] node2704;
	wire [4-1:0] node2705;
	wire [4-1:0] node2707;
	wire [4-1:0] node2710;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2716;
	wire [4-1:0] node2717;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2729;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2746;
	wire [4-1:0] node2747;
	wire [4-1:0] node2753;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2759;
	wire [4-1:0] node2761;
	wire [4-1:0] node2764;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2780;
	wire [4-1:0] node2784;
	wire [4-1:0] node2786;
	wire [4-1:0] node2789;
	wire [4-1:0] node2790;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2795;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2809;
	wire [4-1:0] node2812;
	wire [4-1:0] node2814;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2820;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2826;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2832;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2840;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2846;
	wire [4-1:0] node2849;
	wire [4-1:0] node2851;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2862;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2875;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2880;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2888;
	wire [4-1:0] node2889;
	wire [4-1:0] node2890;
	wire [4-1:0] node2891;
	wire [4-1:0] node2892;
	wire [4-1:0] node2895;
	wire [4-1:0] node2898;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2909;
	wire [4-1:0] node2912;
	wire [4-1:0] node2915;
	wire [4-1:0] node2916;
	wire [4-1:0] node2920;
	wire [4-1:0] node2921;
	wire [4-1:0] node2922;
	wire [4-1:0] node2924;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2932;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2945;
	wire [4-1:0] node2949;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2966;
	wire [4-1:0] node2967;
	wire [4-1:0] node2969;
	wire [4-1:0] node2972;
	wire [4-1:0] node2974;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2981;
	wire [4-1:0] node2984;
	wire [4-1:0] node2985;
	wire [4-1:0] node2987;
	wire [4-1:0] node2991;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2996;
	wire [4-1:0] node2999;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3006;
	wire [4-1:0] node3009;
	wire [4-1:0] node3012;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3025;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3030;
	wire [4-1:0] node3032;
	wire [4-1:0] node3036;
	wire [4-1:0] node3038;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3063;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3072;
	wire [4-1:0] node3076;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3086;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3093;
	wire [4-1:0] node3096;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3104;
	wire [4-1:0] node3105;
	wire [4-1:0] node3109;
	wire [4-1:0] node3110;
	wire [4-1:0] node3113;
	wire [4-1:0] node3114;
	wire [4-1:0] node3118;
	wire [4-1:0] node3119;
	wire [4-1:0] node3120;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3125;
	wire [4-1:0] node3128;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3136;
	wire [4-1:0] node3139;
	wire [4-1:0] node3141;
	wire [4-1:0] node3144;
	wire [4-1:0] node3145;
	wire [4-1:0] node3147;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3153;
	wire [4-1:0] node3156;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3169;
	wire [4-1:0] node3172;
	wire [4-1:0] node3174;
	wire [4-1:0] node3175;
	wire [4-1:0] node3178;
	wire [4-1:0] node3180;
	wire [4-1:0] node3183;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3190;
	wire [4-1:0] node3193;
	wire [4-1:0] node3195;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3206;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3212;
	wire [4-1:0] node3216;
	wire [4-1:0] node3217;
	wire [4-1:0] node3219;
	wire [4-1:0] node3222;
	wire [4-1:0] node3224;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3240;
	wire [4-1:0] node3241;
	wire [4-1:0] node3245;
	wire [4-1:0] node3248;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3252;
	wire [4-1:0] node3255;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3263;
	wire [4-1:0] node3265;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3271;
	wire [4-1:0] node3272;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3279;
	wire [4-1:0] node3282;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3313;
	wire [4-1:0] node3314;
	wire [4-1:0] node3317;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3324;
	wire [4-1:0] node3327;
	wire [4-1:0] node3329;
	wire [4-1:0] node3331;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3340;
	wire [4-1:0] node3341;
	wire [4-1:0] node3344;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3351;
	wire [4-1:0] node3355;
	wire [4-1:0] node3358;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3364;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3371;
	wire [4-1:0] node3372;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3378;
	wire [4-1:0] node3381;
	wire [4-1:0] node3384;
	wire [4-1:0] node3385;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3393;
	wire [4-1:0] node3396;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3405;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3411;
	wire [4-1:0] node3414;
	wire [4-1:0] node3415;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3422;
	wire [4-1:0] node3423;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3431;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3437;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3448;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3455;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3462;
	wire [4-1:0] node3465;
	wire [4-1:0] node3466;
	wire [4-1:0] node3467;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3470;
	wire [4-1:0] node3473;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3478;
	wire [4-1:0] node3480;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3488;
	wire [4-1:0] node3492;
	wire [4-1:0] node3493;
	wire [4-1:0] node3495;
	wire [4-1:0] node3498;
	wire [4-1:0] node3501;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3506;
	wire [4-1:0] node3509;
	wire [4-1:0] node3512;
	wire [4-1:0] node3513;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3531;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3539;
	wire [4-1:0] node3542;
	wire [4-1:0] node3544;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3554;
	wire [4-1:0] node3558;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3577;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3587;
	wire [4-1:0] node3588;
	wire [4-1:0] node3591;
	wire [4-1:0] node3595;
	wire [4-1:0] node3596;
	wire [4-1:0] node3599;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3623;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3641;
	wire [4-1:0] node3643;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3667;
	wire [4-1:0] node3668;
	wire [4-1:0] node3671;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3680;
	wire [4-1:0] node3682;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3688;
	wire [4-1:0] node3690;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3696;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3703;
	wire [4-1:0] node3705;
	wire [4-1:0] node3707;
	wire [4-1:0] node3710;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3724;
	wire [4-1:0] node3725;
	wire [4-1:0] node3728;
	wire [4-1:0] node3729;
	wire [4-1:0] node3732;
	wire [4-1:0] node3735;
	wire [4-1:0] node3736;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3740;
	wire [4-1:0] node3745;
	wire [4-1:0] node3746;
	wire [4-1:0] node3747;
	wire [4-1:0] node3751;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3757;
	wire [4-1:0] node3760;
	wire [4-1:0] node3761;
	wire [4-1:0] node3762;
	wire [4-1:0] node3763;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3770;
	wire [4-1:0] node3774;
	wire [4-1:0] node3775;
	wire [4-1:0] node3777;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3791;
	wire [4-1:0] node3794;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3805;
	wire [4-1:0] node3806;
	wire [4-1:0] node3808;
	wire [4-1:0] node3811;
	wire [4-1:0] node3812;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3819;
	wire [4-1:0] node3821;
	wire [4-1:0] node3824;
	wire [4-1:0] node3827;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3833;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3839;
	wire [4-1:0] node3840;
	wire [4-1:0] node3841;
	wire [4-1:0] node3846;
	wire [4-1:0] node3847;
	wire [4-1:0] node3848;
	wire [4-1:0] node3850;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3861;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3868;
	wire [4-1:0] node3870;
	wire [4-1:0] node3871;
	wire [4-1:0] node3872;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3883;
	wire [4-1:0] node3884;
	wire [4-1:0] node3886;
	wire [4-1:0] node3887;
	wire [4-1:0] node3890;
	wire [4-1:0] node3893;
	wire [4-1:0] node3894;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3912;
	wire [4-1:0] node3914;
	wire [4-1:0] node3917;
	wire [4-1:0] node3918;
	wire [4-1:0] node3919;
	wire [4-1:0] node3920;
	wire [4-1:0] node3923;
	wire [4-1:0] node3927;
	wire [4-1:0] node3929;
	wire [4-1:0] node3931;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3950;
	wire [4-1:0] node3954;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3968;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3978;
	wire [4-1:0] node3981;
	wire [4-1:0] node3983;
	wire [4-1:0] node3986;
	wire [4-1:0] node3987;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3996;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4011;
	wire [4-1:0] node4013;
	wire [4-1:0] node4016;
	wire [4-1:0] node4017;
	wire [4-1:0] node4018;
	wire [4-1:0] node4022;
	wire [4-1:0] node4023;
	wire [4-1:0] node4025;
	wire [4-1:0] node4028;
	wire [4-1:0] node4031;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4037;
	wire [4-1:0] node4039;
	wire [4-1:0] node4042;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4048;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4066;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4074;
	wire [4-1:0] node4076;
	wire [4-1:0] node4079;
	wire [4-1:0] node4080;
	wire [4-1:0] node4081;
	wire [4-1:0] node4086;
	wire [4-1:0] node4088;
	wire [4-1:0] node4091;
	wire [4-1:0] node4092;
	wire [4-1:0] node4094;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4100;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4108;
	wire [4-1:0] node4109;
	wire [4-1:0] node4110;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4123;
	wire [4-1:0] node4124;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4132;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4138;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4151;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4163;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4168;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4175;
	wire [4-1:0] node4177;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4191;
	wire [4-1:0] node4194;
	wire [4-1:0] node4196;
	wire [4-1:0] node4199;
	wire [4-1:0] node4201;
	wire [4-1:0] node4204;
	wire [4-1:0] node4205;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4211;
	wire [4-1:0] node4214;
	wire [4-1:0] node4215;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4221;
	wire [4-1:0] node4222;
	wire [4-1:0] node4223;
	wire [4-1:0] node4227;
	wire [4-1:0] node4229;
	wire [4-1:0] node4232;
	wire [4-1:0] node4233;
	wire [4-1:0] node4234;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4242;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4249;
	wire [4-1:0] node4250;
	wire [4-1:0] node4253;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4260;
	wire [4-1:0] node4263;
	wire [4-1:0] node4265;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4275;
	wire [4-1:0] node4276;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4283;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4290;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4302;
	wire [4-1:0] node4303;
	wire [4-1:0] node4305;
	wire [4-1:0] node4308;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4331;
	wire [4-1:0] node4334;
	wire [4-1:0] node4336;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4344;
	wire [4-1:0] node4346;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4352;
	wire [4-1:0] node4355;
	wire [4-1:0] node4357;
	wire [4-1:0] node4358;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4369;
	wire [4-1:0] node4371;
	wire [4-1:0] node4372;
	wire [4-1:0] node4375;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4383;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4390;
	wire [4-1:0] node4391;
	wire [4-1:0] node4394;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4416;
	wire [4-1:0] node4418;
	wire [4-1:0] node4421;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4433;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4440;
	wire [4-1:0] node4443;
	wire [4-1:0] node4445;
	wire [4-1:0] node4447;
	wire [4-1:0] node4450;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4457;
	wire [4-1:0] node4458;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4467;
	wire [4-1:0] node4470;
	wire [4-1:0] node4473;
	wire [4-1:0] node4474;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4480;
	wire [4-1:0] node4482;
	wire [4-1:0] node4484;
	wire [4-1:0] node4487;
	wire [4-1:0] node4488;
	wire [4-1:0] node4490;
	wire [4-1:0] node4493;
	wire [4-1:0] node4495;
	wire [4-1:0] node4498;
	wire [4-1:0] node4499;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4503;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4518;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4527;
	wire [4-1:0] node4529;
	wire [4-1:0] node4532;
	wire [4-1:0] node4534;
	wire [4-1:0] node4535;
	wire [4-1:0] node4538;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4549;
	wire [4-1:0] node4553;
	wire [4-1:0] node4555;
	wire [4-1:0] node4557;
	wire [4-1:0] node4559;
	wire [4-1:0] node4562;
	wire [4-1:0] node4563;
	wire [4-1:0] node4564;
	wire [4-1:0] node4565;
	wire [4-1:0] node4566;
	wire [4-1:0] node4568;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4575;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4582;
	wire [4-1:0] node4584;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4592;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4599;
	wire [4-1:0] node4602;
	wire [4-1:0] node4605;
	wire [4-1:0] node4607;
	wire [4-1:0] node4608;
	wire [4-1:0] node4611;
	wire [4-1:0] node4614;
	wire [4-1:0] node4615;
	wire [4-1:0] node4616;
	wire [4-1:0] node4617;
	wire [4-1:0] node4619;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4626;
	wire [4-1:0] node4628;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4638;
	wire [4-1:0] node4639;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4648;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4656;
	wire [4-1:0] node4660;
	wire [4-1:0] node4662;
	wire [4-1:0] node4665;
	wire [4-1:0] node4666;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4675;
	wire [4-1:0] node4676;
	wire [4-1:0] node4678;
	wire [4-1:0] node4681;
	wire [4-1:0] node4683;
	wire [4-1:0] node4686;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4690;
	wire [4-1:0] node4693;
	wire [4-1:0] node4694;
	wire [4-1:0] node4697;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4711;
	wire [4-1:0] node4713;
	wire [4-1:0] node4714;
	wire [4-1:0] node4715;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4726;
	wire [4-1:0] node4728;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4734;
	wire [4-1:0] node4738;
	wire [4-1:0] node4739;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4746;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4753;
	wire [4-1:0] node4757;
	wire [4-1:0] node4758;
	wire [4-1:0] node4759;
	wire [4-1:0] node4760;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4770;
	wire [4-1:0] node4775;
	wire [4-1:0] node4778;
	wire [4-1:0] node4779;
	wire [4-1:0] node4781;
	wire [4-1:0] node4782;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4790;
	wire [4-1:0] node4792;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4800;
	wire [4-1:0] node4804;
	wire [4-1:0] node4807;
	wire [4-1:0] node4810;
	wire [4-1:0] node4811;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4819;
	wire [4-1:0] node4820;
	wire [4-1:0] node4823;
	wire [4-1:0] node4826;
	wire [4-1:0] node4828;
	wire [4-1:0] node4830;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4840;
	wire [4-1:0] node4842;
	wire [4-1:0] node4844;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4854;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4863;
	wire [4-1:0] node4864;
	wire [4-1:0] node4865;
	wire [4-1:0] node4868;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4877;
	wire [4-1:0] node4879;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4885;
	wire [4-1:0] node4888;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4894;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4901;
	wire [4-1:0] node4904;
	wire [4-1:0] node4905;
	wire [4-1:0] node4906;
	wire [4-1:0] node4907;
	wire [4-1:0] node4909;
	wire [4-1:0] node4912;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4919;
	wire [4-1:0] node4922;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4940;
	wire [4-1:0] node4942;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4949;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4954;
	wire [4-1:0] node4957;
	wire [4-1:0] node4959;
	wire [4-1:0] node4963;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4972;
	wire [4-1:0] node4975;
	wire [4-1:0] node4977;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4989;
	wire [4-1:0] node4992;
	wire [4-1:0] node4993;
	wire [4-1:0] node4997;
	wire [4-1:0] node4998;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5002;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5011;
	wire [4-1:0] node5014;
	wire [4-1:0] node5015;
	wire [4-1:0] node5016;
	wire [4-1:0] node5020;
	wire [4-1:0] node5021;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5028;
	wire [4-1:0] node5031;
	wire [4-1:0] node5032;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5038;
	wire [4-1:0] node5041;
	wire [4-1:0] node5043;
	wire [4-1:0] node5046;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5052;
	wire [4-1:0] node5056;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5061;
	wire [4-1:0] node5065;
	wire [4-1:0] node5068;
	wire [4-1:0] node5069;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5073;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5080;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5090;
	wire [4-1:0] node5091;
	wire [4-1:0] node5093;
	wire [4-1:0] node5097;
	wire [4-1:0] node5098;
	wire [4-1:0] node5099;
	wire [4-1:0] node5101;
	wire [4-1:0] node5102;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5109;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5118;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5136;
	wire [4-1:0] node5139;
	wire [4-1:0] node5140;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5148;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5153;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5160;
	wire [4-1:0] node5163;
	wire [4-1:0] node5164;
	wire [4-1:0] node5165;
	wire [4-1:0] node5168;
	wire [4-1:0] node5170;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5176;
	wire [4-1:0] node5179;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5184;
	wire [4-1:0] node5186;
	wire [4-1:0] node5189;
	wire [4-1:0] node5190;
	wire [4-1:0] node5191;
	wire [4-1:0] node5193;
	wire [4-1:0] node5197;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5209;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5214;
	wire [4-1:0] node5215;
	wire [4-1:0] node5219;
	wire [4-1:0] node5221;
	wire [4-1:0] node5222;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5229;
	wire [4-1:0] node5230;
	wire [4-1:0] node5233;
	wire [4-1:0] node5236;
	wire [4-1:0] node5237;
	wire [4-1:0] node5240;
	wire [4-1:0] node5242;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5250;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5257;
	wire [4-1:0] node5261;
	wire [4-1:0] node5263;
	wire [4-1:0] node5266;
	wire [4-1:0] node5268;
	wire [4-1:0] node5269;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5282;
	wire [4-1:0] node5285;
	wire [4-1:0] node5289;
	wire [4-1:0] node5291;
	wire [4-1:0] node5292;
	wire [4-1:0] node5295;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5300;
	wire [4-1:0] node5302;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5313;
	wire [4-1:0] node5316;
	wire [4-1:0] node5317;
	wire [4-1:0] node5319;
	wire [4-1:0] node5321;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5327;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5333;
	wire [4-1:0] node5334;
	wire [4-1:0] node5335;
	wire [4-1:0] node5338;
	wire [4-1:0] node5340;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5361;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5379;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5384;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5392;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5398;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5412;
	wire [4-1:0] node5414;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5420;
	wire [4-1:0] node5422;
	wire [4-1:0] node5425;
	wire [4-1:0] node5428;
	wire [4-1:0] node5429;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5434;
	wire [4-1:0] node5435;
	wire [4-1:0] node5438;
	wire [4-1:0] node5441;
	wire [4-1:0] node5442;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5449;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5454;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5460;
	wire [4-1:0] node5463;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5470;
	wire [4-1:0] node5471;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5488;
	wire [4-1:0] node5489;
	wire [4-1:0] node5491;
	wire [4-1:0] node5494;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5506;
	wire [4-1:0] node5509;
	wire [4-1:0] node5510;
	wire [4-1:0] node5514;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5523;
	wire [4-1:0] node5525;
	wire [4-1:0] node5528;
	wire [4-1:0] node5529;
	wire [4-1:0] node5532;
	wire [4-1:0] node5536;
	wire [4-1:0] node5537;
	wire [4-1:0] node5539;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5550;
	wire [4-1:0] node5552;
	wire [4-1:0] node5555;
	wire [4-1:0] node5556;
	wire [4-1:0] node5557;
	wire [4-1:0] node5560;
	wire [4-1:0] node5562;
	wire [4-1:0] node5565;
	wire [4-1:0] node5567;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5574;
	wire [4-1:0] node5575;
	wire [4-1:0] node5578;
	wire [4-1:0] node5581;
	wire [4-1:0] node5584;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5594;
	wire [4-1:0] node5597;
	wire [4-1:0] node5600;
	wire [4-1:0] node5603;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5611;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5619;
	wire [4-1:0] node5621;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5627;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5634;
	wire [4-1:0] node5637;
	wire [4-1:0] node5638;
	wire [4-1:0] node5639;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5645;
	wire [4-1:0] node5646;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5653;
	wire [4-1:0] node5656;
	wire [4-1:0] node5658;
	wire [4-1:0] node5661;
	wire [4-1:0] node5662;
	wire [4-1:0] node5664;
	wire [4-1:0] node5665;
	wire [4-1:0] node5668;
	wire [4-1:0] node5671;
	wire [4-1:0] node5674;
	wire [4-1:0] node5675;
	wire [4-1:0] node5676;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5683;
	wire [4-1:0] node5686;
	wire [4-1:0] node5687;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5701;
	wire [4-1:0] node5703;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5719;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5726;
	wire [4-1:0] node5728;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5734;
	wire [4-1:0] node5737;
	wire [4-1:0] node5738;
	wire [4-1:0] node5742;
	wire [4-1:0] node5743;
	wire [4-1:0] node5744;
	wire [4-1:0] node5745;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5751;
	wire [4-1:0] node5753;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5762;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5769;
	wire [4-1:0] node5771;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5777;
	wire [4-1:0] node5780;
	wire [4-1:0] node5783;
	wire [4-1:0] node5785;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5802;
	wire [4-1:0] node5804;
	wire [4-1:0] node5806;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5819;
	wire [4-1:0] node5821;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5839;
	wire [4-1:0] node5841;
	wire [4-1:0] node5845;
	wire [4-1:0] node5847;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5857;
	wire [4-1:0] node5860;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5867;
	wire [4-1:0] node5871;
	wire [4-1:0] node5872;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5878;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5885;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5893;
	wire [4-1:0] node5895;
	wire [4-1:0] node5896;
	wire [4-1:0] node5899;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5906;
	wire [4-1:0] node5908;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5916;
	wire [4-1:0] node5917;
	wire [4-1:0] node5918;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5925;
	wire [4-1:0] node5928;
	wire [4-1:0] node5930;
	wire [4-1:0] node5932;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5937;
	wire [4-1:0] node5938;
	wire [4-1:0] node5941;
	wire [4-1:0] node5944;
	wire [4-1:0] node5947;
	wire [4-1:0] node5948;
	wire [4-1:0] node5949;
	wire [4-1:0] node5951;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5962;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5968;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5977;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5983;
	wire [4-1:0] node5984;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5991;
	wire [4-1:0] node5992;
	wire [4-1:0] node5995;
	wire [4-1:0] node5998;
	wire [4-1:0] node5999;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6006;
	wire [4-1:0] node6007;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6017;
	wire [4-1:0] node6019;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6026;
	wire [4-1:0] node6027;
	wire [4-1:0] node6028;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6034;
	wire [4-1:0] node6036;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6041;
	wire [4-1:0] node6044;
	wire [4-1:0] node6047;
	wire [4-1:0] node6049;
	wire [4-1:0] node6051;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6057;
	wire [4-1:0] node6059;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6068;
	wire [4-1:0] node6069;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6075;
	wire [4-1:0] node6076;
	wire [4-1:0] node6077;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6084;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6093;
	wire [4-1:0] node6095;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6104;
	wire [4-1:0] node6107;
	wire [4-1:0] node6108;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6116;
	wire [4-1:0] node6117;
	wire [4-1:0] node6118;
	wire [4-1:0] node6121;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6127;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6136;
	wire [4-1:0] node6138;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6144;
	wire [4-1:0] node6147;
	wire [4-1:0] node6150;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6156;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6166;
	wire [4-1:0] node6167;
	wire [4-1:0] node6170;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6179;
	wire [4-1:0] node6180;
	wire [4-1:0] node6181;
	wire [4-1:0] node6184;
	wire [4-1:0] node6187;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6192;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6202;
	wire [4-1:0] node6205;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6211;
	wire [4-1:0] node6213;
	wire [4-1:0] node6216;
	wire [4-1:0] node6217;
	wire [4-1:0] node6219;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6230;
	wire [4-1:0] node6231;
	wire [4-1:0] node6235;
	wire [4-1:0] node6237;
	wire [4-1:0] node6240;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6246;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6261;
	wire [4-1:0] node6264;
	wire [4-1:0] node6267;
	wire [4-1:0] node6268;
	wire [4-1:0] node6269;
	wire [4-1:0] node6274;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6279;
	wire [4-1:0] node6282;
	wire [4-1:0] node6285;
	wire [4-1:0] node6287;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6292;
	wire [4-1:0] node6297;
	wire [4-1:0] node6298;
	wire [4-1:0] node6299;
	wire [4-1:0] node6300;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6307;
	wire [4-1:0] node6310;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6320;
	wire [4-1:0] node6321;
	wire [4-1:0] node6322;
	wire [4-1:0] node6325;
	wire [4-1:0] node6328;
	wire [4-1:0] node6329;
	wire [4-1:0] node6333;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6344;
	wire [4-1:0] node6347;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6356;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6362;
	wire [4-1:0] node6365;
	wire [4-1:0] node6368;
	wire [4-1:0] node6371;
	wire [4-1:0] node6372;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6378;
	wire [4-1:0] node6381;
	wire [4-1:0] node6383;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6389;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6399;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6402;
	wire [4-1:0] node6406;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6413;
	wire [4-1:0] node6414;
	wire [4-1:0] node6415;
	wire [4-1:0] node6417;
	wire [4-1:0] node6420;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6427;
	wire [4-1:0] node6428;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6435;
	wire [4-1:0] node6436;
	wire [4-1:0] node6438;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6445;
	wire [4-1:0] node6448;
	wire [4-1:0] node6449;
	wire [4-1:0] node6452;
	wire [4-1:0] node6453;
	wire [4-1:0] node6457;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6461;
	wire [4-1:0] node6464;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6469;
	wire [4-1:0] node6473;
	wire [4-1:0] node6475;
	wire [4-1:0] node6477;
	wire [4-1:0] node6480;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6484;
	wire [4-1:0] node6487;
	wire [4-1:0] node6488;
	wire [4-1:0] node6491;
	wire [4-1:0] node6494;
	wire [4-1:0] node6495;
	wire [4-1:0] node6497;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6513;
	wire [4-1:0] node6514;
	wire [4-1:0] node6515;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6525;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6530;
	wire [4-1:0] node6533;
	wire [4-1:0] node6536;
	wire [4-1:0] node6538;
	wire [4-1:0] node6541;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6544;
	wire [4-1:0] node6548;
	wire [4-1:0] node6549;
	wire [4-1:0] node6552;
	wire [4-1:0] node6555;
	wire [4-1:0] node6556;
	wire [4-1:0] node6557;
	wire [4-1:0] node6560;
	wire [4-1:0] node6564;
	wire [4-1:0] node6565;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6569;
	wire [4-1:0] node6572;
	wire [4-1:0] node6573;
	wire [4-1:0] node6576;
	wire [4-1:0] node6579;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6596;
	wire [4-1:0] node6599;
	wire [4-1:0] node6600;
	wire [4-1:0] node6602;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6610;
	wire [4-1:0] node6611;
	wire [4-1:0] node6612;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6628;
	wire [4-1:0] node6631;
	wire [4-1:0] node6632;
	wire [4-1:0] node6633;
	wire [4-1:0] node6634;
	wire [4-1:0] node6635;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6652;
	wire [4-1:0] node6653;
	wire [4-1:0] node6654;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6662;
	wire [4-1:0] node6663;
	wire [4-1:0] node6665;
	wire [4-1:0] node6668;
	wire [4-1:0] node6670;
	wire [4-1:0] node6673;
	wire [4-1:0] node6674;
	wire [4-1:0] node6675;
	wire [4-1:0] node6676;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6684;
	wire [4-1:0] node6687;
	wire [4-1:0] node6688;
	wire [4-1:0] node6689;
	wire [4-1:0] node6691;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6699;
	wire [4-1:0] node6700;
	wire [4-1:0] node6702;
	wire [4-1:0] node6705;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6711;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6717;
	wire [4-1:0] node6718;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6734;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6738;
	wire [4-1:0] node6743;
	wire [4-1:0] node6745;
	wire [4-1:0] node6749;
	wire [4-1:0] node6750;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6761;
	wire [4-1:0] node6764;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6770;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6775;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6782;
	wire [4-1:0] node6783;
	wire [4-1:0] node6787;
	wire [4-1:0] node6788;
	wire [4-1:0] node6792;
	wire [4-1:0] node6793;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6798;
	wire [4-1:0] node6801;
	wire [4-1:0] node6804;
	wire [4-1:0] node6805;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6816;
	wire [4-1:0] node6817;
	wire [4-1:0] node6821;
	wire [4-1:0] node6822;
	wire [4-1:0] node6825;
	wire [4-1:0] node6826;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6838;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6858;
	wire [4-1:0] node6859;
	wire [4-1:0] node6860;
	wire [4-1:0] node6862;
	wire [4-1:0] node6865;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6879;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6895;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6901;
	wire [4-1:0] node6902;
	wire [4-1:0] node6905;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6910;
	wire [4-1:0] node6914;
	wire [4-1:0] node6915;
	wire [4-1:0] node6918;
	wire [4-1:0] node6920;
	wire [4-1:0] node6923;
	wire [4-1:0] node6924;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6931;
	wire [4-1:0] node6933;
	wire [4-1:0] node6936;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6942;
	wire [4-1:0] node6945;
	wire [4-1:0] node6947;
	wire [4-1:0] node6949;
	wire [4-1:0] node6952;
	wire [4-1:0] node6953;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6957;
	wire [4-1:0] node6960;
	wire [4-1:0] node6962;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6968;
	wire [4-1:0] node6971;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6982;
	wire [4-1:0] node6985;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6994;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node6999;
	wire [4-1:0] node7003;
	wire [4-1:0] node7006;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7009;
	wire [4-1:0] node7013;
	wire [4-1:0] node7015;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7022;
	wire [4-1:0] node7023;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7031;
	wire [4-1:0] node7032;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7039;
	wire [4-1:0] node7040;
	wire [4-1:0] node7043;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7053;
	wire [4-1:0] node7054;
	wire [4-1:0] node7055;
	wire [4-1:0] node7056;
	wire [4-1:0] node7059;
	wire [4-1:0] node7062;
	wire [4-1:0] node7064;
	wire [4-1:0] node7067;
	wire [4-1:0] node7068;
	wire [4-1:0] node7069;
	wire [4-1:0] node7073;
	wire [4-1:0] node7074;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7081;
	wire [4-1:0] node7082;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7089;
	wire [4-1:0] node7092;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7096;
	wire [4-1:0] node7099;
	wire [4-1:0] node7103;
	wire [4-1:0] node7104;
	wire [4-1:0] node7107;
	wire [4-1:0] node7108;
	wire [4-1:0] node7110;
	wire [4-1:0] node7114;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7119;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7126;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7132;
	wire [4-1:0] node7135;
	wire [4-1:0] node7137;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7145;
	wire [4-1:0] node7149;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7155;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7162;
	wire [4-1:0] node7165;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7170;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7177;
	wire [4-1:0] node7180;
	wire [4-1:0] node7182;
	wire [4-1:0] node7185;
	wire [4-1:0] node7188;
	wire [4-1:0] node7190;
	wire [4-1:0] node7191;
	wire [4-1:0] node7193;
	wire [4-1:0] node7196;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7203;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7208;
	wire [4-1:0] node7212;
	wire [4-1:0] node7213;
	wire [4-1:0] node7215;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7238;
	wire [4-1:0] node7243;
	wire [4-1:0] node7244;
	wire [4-1:0] node7245;
	wire [4-1:0] node7247;
	wire [4-1:0] node7250;
	wire [4-1:0] node7253;
	wire [4-1:0] node7255;
	wire [4-1:0] node7258;
	wire [4-1:0] node7259;
	wire [4-1:0] node7260;
	wire [4-1:0] node7263;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7270;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7276;
	wire [4-1:0] node7277;
	wire [4-1:0] node7281;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7286;
	wire [4-1:0] node7292;
	wire [4-1:0] node7293;
	wire [4-1:0] node7296;
	wire [4-1:0] node7299;
	wire [4-1:0] node7300;
	wire [4-1:0] node7301;
	wire [4-1:0] node7303;
	wire [4-1:0] node7307;
	wire [4-1:0] node7309;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7328;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7337;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7346;
	wire [4-1:0] node7349;
	wire [4-1:0] node7351;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7371;
	wire [4-1:0] node7373;
	wire [4-1:0] node7376;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7382;
	wire [4-1:0] node7383;
	wire [4-1:0] node7384;
	wire [4-1:0] node7385;
	wire [4-1:0] node7386;
	wire [4-1:0] node7388;
	wire [4-1:0] node7389;
	wire [4-1:0] node7392;
	wire [4-1:0] node7395;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7401;
	wire [4-1:0] node7404;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7408;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7416;
	wire [4-1:0] node7419;
	wire [4-1:0] node7420;
	wire [4-1:0] node7424;
	wire [4-1:0] node7425;
	wire [4-1:0] node7426;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7435;
	wire [4-1:0] node7438;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7444;
	wire [4-1:0] node7445;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7456;
	wire [4-1:0] node7460;
	wire [4-1:0] node7462;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7468;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7473;
	wire [4-1:0] node7474;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7484;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7490;
	wire [4-1:0] node7493;
	wire [4-1:0] node7494;
	wire [4-1:0] node7497;
	wire [4-1:0] node7500;
	wire [4-1:0] node7501;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7504;
	wire [4-1:0] node7506;
	wire [4-1:0] node7510;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7515;
	wire [4-1:0] node7518;
	wire [4-1:0] node7519;
	wire [4-1:0] node7521;
	wire [4-1:0] node7525;
	wire [4-1:0] node7526;
	wire [4-1:0] node7527;
	wire [4-1:0] node7528;
	wire [4-1:0] node7532;
	wire [4-1:0] node7535;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7543;
	wire [4-1:0] node7546;
	wire [4-1:0] node7547;
	wire [4-1:0] node7548;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7553;
	wire [4-1:0] node7556;
	wire [4-1:0] node7558;
	wire [4-1:0] node7561;
	wire [4-1:0] node7563;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7568;
	wire [4-1:0] node7569;
	wire [4-1:0] node7572;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7579;
	wire [4-1:0] node7582;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7585;
	wire [4-1:0] node7590;
	wire [4-1:0] node7593;
	wire [4-1:0] node7594;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7600;
	wire [4-1:0] node7604;
	wire [4-1:0] node7605;
	wire [4-1:0] node7607;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7620;
	wire [4-1:0] node7621;
	wire [4-1:0] node7623;
	wire [4-1:0] node7627;
	wire [4-1:0] node7629;
	wire [4-1:0] node7632;
	wire [4-1:0] node7633;
	wire [4-1:0] node7634;
	wire [4-1:0] node7636;
	wire [4-1:0] node7638;
	wire [4-1:0] node7641;
	wire [4-1:0] node7643;
	wire [4-1:0] node7646;
	wire [4-1:0] node7647;
	wire [4-1:0] node7648;
	wire [4-1:0] node7651;
	wire [4-1:0] node7654;
	wire [4-1:0] node7655;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7663;
	wire [4-1:0] node7664;
	wire [4-1:0] node7665;
	wire [4-1:0] node7666;
	wire [4-1:0] node7667;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7674;
	wire [4-1:0] node7677;
	wire [4-1:0] node7678;
	wire [4-1:0] node7680;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7688;
	wire [4-1:0] node7689;
	wire [4-1:0] node7690;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7708;
	wire [4-1:0] node7712;
	wire [4-1:0] node7713;
	wire [4-1:0] node7716;
	wire [4-1:0] node7719;
	wire [4-1:0] node7720;
	wire [4-1:0] node7722;
	wire [4-1:0] node7725;
	wire [4-1:0] node7726;
	wire [4-1:0] node7729;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7741;
	wire [4-1:0] node7744;
	wire [4-1:0] node7745;
	wire [4-1:0] node7749;
	wire [4-1:0] node7751;
	wire [4-1:0] node7752;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7759;
	wire [4-1:0] node7760;
	wire [4-1:0] node7764;
	wire [4-1:0] node7766;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7772;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7777;
	wire [4-1:0] node7778;
	wire [4-1:0] node7781;
	wire [4-1:0] node7785;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7800;
	wire [4-1:0] node7802;
	wire [4-1:0] node7805;
	wire [4-1:0] node7807;
	wire [4-1:0] node7809;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7818;
	wire [4-1:0] node7819;
	wire [4-1:0] node7821;
	wire [4-1:0] node7824;
	wire [4-1:0] node7825;
	wire [4-1:0] node7827;
	wire [4-1:0] node7831;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7841;
	wire [4-1:0] node7844;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7849;
	wire [4-1:0] node7852;
	wire [4-1:0] node7854;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7861;
	wire [4-1:0] node7862;
	wire [4-1:0] node7864;
	wire [4-1:0] node7868;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7876;
	wire [4-1:0] node7877;
	wire [4-1:0] node7878;
	wire [4-1:0] node7881;
	wire [4-1:0] node7883;
	wire [4-1:0] node7887;
	wire [4-1:0] node7888;
	wire [4-1:0] node7889;
	wire [4-1:0] node7890;
	wire [4-1:0] node7891;
	wire [4-1:0] node7894;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7902;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7911;
	wire [4-1:0] node7913;
	wire [4-1:0] node7916;
	wire [4-1:0] node7917;
	wire [4-1:0] node7918;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7926;
	wire [4-1:0] node7928;
	wire [4-1:0] node7931;
	wire [4-1:0] node7932;
	wire [4-1:0] node7935;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7940;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7946;
	wire [4-1:0] node7949;
	wire [4-1:0] node7951;
	wire [4-1:0] node7952;
	wire [4-1:0] node7953;
	wire [4-1:0] node7956;
	wire [4-1:0] node7959;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7964;
	wire [4-1:0] node7968;
	wire [4-1:0] node7969;
	wire [4-1:0] node7972;
	wire [4-1:0] node7973;
	wire [4-1:0] node7976;
	wire [4-1:0] node7979;
	wire [4-1:0] node7980;
	wire [4-1:0] node7981;
	wire [4-1:0] node7982;
	wire [4-1:0] node7985;
	wire [4-1:0] node7987;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7992;
	wire [4-1:0] node7994;
	wire [4-1:0] node7997;
	wire [4-1:0] node8001;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8005;
	wire [4-1:0] node8009;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8015;
	wire [4-1:0] node8018;
	wire [4-1:0] node8021;
	wire [4-1:0] node8023;
	wire [4-1:0] node8026;
	wire [4-1:0] node8027;
	wire [4-1:0] node8028;
	wire [4-1:0] node8029;
	wire [4-1:0] node8031;
	wire [4-1:0] node8032;
	wire [4-1:0] node8034;
	wire [4-1:0] node8038;
	wire [4-1:0] node8039;
	wire [4-1:0] node8040;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8061;
	wire [4-1:0] node8064;
	wire [4-1:0] node8067;
	wire [4-1:0] node8068;
	wire [4-1:0] node8071;
	wire [4-1:0] node8074;
	wire [4-1:0] node8075;
	wire [4-1:0] node8076;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8086;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8096;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8104;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8108;
	wire [4-1:0] node8112;
	wire [4-1:0] node8115;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8121;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8128;
	wire [4-1:0] node8129;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8136;
	wire [4-1:0] node8139;
	wire [4-1:0] node8140;
	wire [4-1:0] node8141;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8148;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8157;
	wire [4-1:0] node8160;
	wire [4-1:0] node8161;
	wire [4-1:0] node8162;
	wire [4-1:0] node8164;
	wire [4-1:0] node8166;
	wire [4-1:0] node8169;
	wire [4-1:0] node8170;
	wire [4-1:0] node8171;
	wire [4-1:0] node8174;
	wire [4-1:0] node8177;
	wire [4-1:0] node8178;
	wire [4-1:0] node8181;
	wire [4-1:0] node8184;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8190;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8197;
	wire [4-1:0] node8200;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8205;
	wire [4-1:0] node8209;
	wire [4-1:0] node8210;
	wire [4-1:0] node8211;
	wire [4-1:0] node8212;
	wire [4-1:0] node8214;
	wire [4-1:0] node8215;
	wire [4-1:0] node8218;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8223;
	wire [4-1:0] node8226;
	wire [4-1:0] node8229;
	wire [4-1:0] node8230;
	wire [4-1:0] node8231;
	wire [4-1:0] node8235;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8242;
	wire [4-1:0] node8244;
	wire [4-1:0] node8246;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8256;
	wire [4-1:0] node8257;
	wire [4-1:0] node8260;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8268;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8275;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8282;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8289;
	wire [4-1:0] node8290;
	wire [4-1:0] node8291;
	wire [4-1:0] node8292;
	wire [4-1:0] node8293;
	wire [4-1:0] node8297;
	wire [4-1:0] node8299;
	wire [4-1:0] node8302;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8309;
	wire [4-1:0] node8310;
	wire [4-1:0] node8312;
	wire [4-1:0] node8315;
	wire [4-1:0] node8317;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8326;
	wire [4-1:0] node8327;
	wire [4-1:0] node8330;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8337;
	wire [4-1:0] node8338;
	wire [4-1:0] node8339;
	wire [4-1:0] node8344;
	wire [4-1:0] node8345;
	wire [4-1:0] node8347;
	wire [4-1:0] node8350;
	wire [4-1:0] node8351;
	wire [4-1:0] node8354;
	wire [4-1:0] node8356;
	wire [4-1:0] node8358;
	wire [4-1:0] node8361;
	wire [4-1:0] node8362;
	wire [4-1:0] node8363;
	wire [4-1:0] node8364;
	wire [4-1:0] node8366;
	wire [4-1:0] node8367;
	wire [4-1:0] node8370;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8381;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8396;
	wire [4-1:0] node8399;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8419;
	wire [4-1:0] node8421;
	wire [4-1:0] node8424;
	wire [4-1:0] node8425;
	wire [4-1:0] node8427;
	wire [4-1:0] node8430;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8435;
	wire [4-1:0] node8437;
	wire [4-1:0] node8439;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8455;
	wire [4-1:0] node8457;
	wire [4-1:0] node8458;
	wire [4-1:0] node8461;
	wire [4-1:0] node8464;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8467;
	wire [4-1:0] node8469;
	wire [4-1:0] node8472;
	wire [4-1:0] node8473;
	wire [4-1:0] node8477;
	wire [4-1:0] node8478;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8483;
	wire [4-1:0] node8487;
	wire [4-1:0] node8489;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8494;
	wire [4-1:0] node8495;
	wire [4-1:0] node8497;
	wire [4-1:0] node8501;
	wire [4-1:0] node8503;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8510;
	wire [4-1:0] node8512;
	wire [4-1:0] node8515;
	wire [4-1:0] node8516;
	wire [4-1:0] node8517;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8524;
	wire [4-1:0] node8525;
	wire [4-1:0] node8528;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8540;
	wire [4-1:0] node8543;
	wire [4-1:0] node8545;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8552;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8559;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8565;
	wire [4-1:0] node8567;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8575;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8588;
	wire [4-1:0] node8590;
	wire [4-1:0] node8594;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8603;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8629;
	wire [4-1:0] node8632;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8640;
	wire [4-1:0] node8642;
	wire [4-1:0] node8645;
	wire [4-1:0] node8647;
	wire [4-1:0] node8650;
	wire [4-1:0] node8651;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8657;
	wire [4-1:0] node8658;
	wire [4-1:0] node8661;
	wire [4-1:0] node8664;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8672;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8683;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8689;
	wire [4-1:0] node8690;
	wire [4-1:0] node8694;
	wire [4-1:0] node8695;
	wire [4-1:0] node8700;
	wire [4-1:0] node8701;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8710;
	wire [4-1:0] node8712;
	wire [4-1:0] node8715;
	wire [4-1:0] node8716;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8720;
	wire [4-1:0] node8721;
	wire [4-1:0] node8725;
	wire [4-1:0] node8726;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8742;
	wire [4-1:0] node8743;
	wire [4-1:0] node8746;
	wire [4-1:0] node8747;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8755;
	wire [4-1:0] node8756;
	wire [4-1:0] node8760;
	wire [4-1:0] node8761;
	wire [4-1:0] node8762;
	wire [4-1:0] node8763;
	wire [4-1:0] node8765;
	wire [4-1:0] node8768;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8777;
	wire [4-1:0] node8781;
	wire [4-1:0] node8783;
	wire [4-1:0] node8786;
	wire [4-1:0] node8787;
	wire [4-1:0] node8789;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8797;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8802;
	wire [4-1:0] node8804;
	wire [4-1:0] node8807;
	wire [4-1:0] node8810;
	wire [4-1:0] node8811;
	wire [4-1:0] node8813;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8824;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8834;
	wire [4-1:0] node8837;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8844;
	wire [4-1:0] node8848;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8859;
	wire [4-1:0] node8860;
	wire [4-1:0] node8864;
	wire [4-1:0] node8865;
	wire [4-1:0] node8868;
	wire [4-1:0] node8871;
	wire [4-1:0] node8872;
	wire [4-1:0] node8873;
	wire [4-1:0] node8876;
	wire [4-1:0] node8878;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8885;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8891;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8898;
	wire [4-1:0] node8899;
	wire [4-1:0] node8900;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8905;
	wire [4-1:0] node8908;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8916;
	wire [4-1:0] node8919;
	wire [4-1:0] node8920;
	wire [4-1:0] node8921;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8933;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8940;
	wire [4-1:0] node8943;
	wire [4-1:0] node8944;
	wire [4-1:0] node8946;
	wire [4-1:0] node8949;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8958;
	wire [4-1:0] node8959;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8972;
	wire [4-1:0] node8974;
	wire [4-1:0] node8977;
	wire [4-1:0] node8978;
	wire [4-1:0] node8981;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8993;
	wire [4-1:0] node8996;
	wire [4-1:0] node8997;
	wire [4-1:0] node9001;
	wire [4-1:0] node9002;
	wire [4-1:0] node9005;
	wire [4-1:0] node9006;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9013;
	wire [4-1:0] node9014;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9020;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9026;
	wire [4-1:0] node9027;
	wire [4-1:0] node9031;
	wire [4-1:0] node9034;
	wire [4-1:0] node9035;
	wire [4-1:0] node9036;
	wire [4-1:0] node9039;
	wire [4-1:0] node9043;
	wire [4-1:0] node9044;
	wire [4-1:0] node9046;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9061;
	wire [4-1:0] node9064;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9073;
	wire [4-1:0] node9075;
	wire [4-1:0] node9078;
	wire [4-1:0] node9080;
	wire [4-1:0] node9083;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9090;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9093;
	wire [4-1:0] node9094;
	wire [4-1:0] node9099;
	wire [4-1:0] node9101;
	wire [4-1:0] node9104;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9109;
	wire [4-1:0] node9112;
	wire [4-1:0] node9113;
	wire [4-1:0] node9115;
	wire [4-1:0] node9118;
	wire [4-1:0] node9119;
	wire [4-1:0] node9123;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9134;
	wire [4-1:0] node9137;
	wire [4-1:0] node9138;
	wire [4-1:0] node9141;
	wire [4-1:0] node9143;
	wire [4-1:0] node9146;
	wire [4-1:0] node9147;
	wire [4-1:0] node9148;
	wire [4-1:0] node9149;
	wire [4-1:0] node9154;
	wire [4-1:0] node9155;
	wire [4-1:0] node9157;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9167;
	wire [4-1:0] node9170;
	wire [4-1:0] node9172;
	wire [4-1:0] node9175;
	wire [4-1:0] node9176;
	wire [4-1:0] node9177;
	wire [4-1:0] node9181;
	wire [4-1:0] node9184;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9187;
	wire [4-1:0] node9190;
	wire [4-1:0] node9191;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9197;
	wire [4-1:0] node9200;
	wire [4-1:0] node9203;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9209;
	wire [4-1:0] node9213;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9219;
	wire [4-1:0] node9222;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9228;
	wire [4-1:0] node9229;
	wire [4-1:0] node9230;
	wire [4-1:0] node9233;
	wire [4-1:0] node9234;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9242;
	wire [4-1:0] node9245;
	wire [4-1:0] node9246;
	wire [4-1:0] node9247;
	wire [4-1:0] node9250;
	wire [4-1:0] node9254;
	wire [4-1:0] node9255;
	wire [4-1:0] node9256;
	wire [4-1:0] node9259;
	wire [4-1:0] node9262;
	wire [4-1:0] node9263;
	wire [4-1:0] node9266;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9271;
	wire [4-1:0] node9272;
	wire [4-1:0] node9274;
	wire [4-1:0] node9277;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9285;
	wire [4-1:0] node9288;
	wire [4-1:0] node9291;
	wire [4-1:0] node9292;
	wire [4-1:0] node9293;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9300;
	wire [4-1:0] node9303;
	wire [4-1:0] node9305;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9316;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9322;
	wire [4-1:0] node9325;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9331;
	wire [4-1:0] node9333;
	wire [4-1:0] node9336;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9343;
	wire [4-1:0] node9344;
	wire [4-1:0] node9346;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9356;
	wire [4-1:0] node9357;
	wire [4-1:0] node9361;
	wire [4-1:0] node9363;
	wire [4-1:0] node9364;
	wire [4-1:0] node9367;
	wire [4-1:0] node9370;
	wire [4-1:0] node9371;
	wire [4-1:0] node9373;
	wire [4-1:0] node9375;
	wire [4-1:0] node9378;
	wire [4-1:0] node9379;
	wire [4-1:0] node9380;
	wire [4-1:0] node9382;
	wire [4-1:0] node9385;
	wire [4-1:0] node9388;
	wire [4-1:0] node9389;
	wire [4-1:0] node9391;
	wire [4-1:0] node9395;
	wire [4-1:0] node9396;
	wire [4-1:0] node9397;
	wire [4-1:0] node9398;
	wire [4-1:0] node9399;
	wire [4-1:0] node9402;
	wire [4-1:0] node9405;
	wire [4-1:0] node9406;
	wire [4-1:0] node9407;
	wire [4-1:0] node9408;
	wire [4-1:0] node9412;
	wire [4-1:0] node9414;
	wire [4-1:0] node9417;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9424;
	wire [4-1:0] node9427;
	wire [4-1:0] node9429;
	wire [4-1:0] node9431;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9436;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9445;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9449;
	wire [4-1:0] node9450;
	wire [4-1:0] node9454;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9460;
	wire [4-1:0] node9461;
	wire [4-1:0] node9464;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9469;
	wire [4-1:0] node9471;
	wire [4-1:0] node9474;
	wire [4-1:0] node9477;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9480;
	wire [4-1:0] node9484;
	wire [4-1:0] node9487;
	wire [4-1:0] node9490;
	wire [4-1:0] node9491;
	wire [4-1:0] node9492;
	wire [4-1:0] node9493;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9496;
	wire [4-1:0] node9499;
	wire [4-1:0] node9502;
	wire [4-1:0] node9504;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9510;
	wire [4-1:0] node9512;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9526;
	wire [4-1:0] node9528;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9544;
	wire [4-1:0] node9548;
	wire [4-1:0] node9551;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9555;
	wire [4-1:0] node9556;
	wire [4-1:0] node9559;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9565;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9572;
	wire [4-1:0] node9574;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9580;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9588;
	wire [4-1:0] node9592;
	wire [4-1:0] node9593;
	wire [4-1:0] node9594;
	wire [4-1:0] node9595;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9601;
	wire [4-1:0] node9602;
	wire [4-1:0] node9605;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9615;
	wire [4-1:0] node9618;
	wire [4-1:0] node9620;
	wire [4-1:0] node9622;
	wire [4-1:0] node9625;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9629;
	wire [4-1:0] node9632;
	wire [4-1:0] node9633;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9639;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9648;
	wire [4-1:0] node9651;
	wire [4-1:0] node9653;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9665;
	wire [4-1:0] node9668;
	wire [4-1:0] node9671;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9676;
	wire [4-1:0] node9679;
	wire [4-1:0] node9681;
	wire [4-1:0] node9684;
	wire [4-1:0] node9685;
	wire [4-1:0] node9686;
	wire [4-1:0] node9689;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9701;
	wire [4-1:0] node9702;
	wire [4-1:0] node9703;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9709;
	wire [4-1:0] node9713;
	wire [4-1:0] node9714;
	wire [4-1:0] node9715;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9723;
	wire [4-1:0] node9726;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9731;
	wire [4-1:0] node9732;
	wire [4-1:0] node9737;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9741;
	wire [4-1:0] node9744;
	wire [4-1:0] node9745;
	wire [4-1:0] node9748;
	wire [4-1:0] node9750;
	wire [4-1:0] node9753;
	wire [4-1:0] node9754;
	wire [4-1:0] node9755;
	wire [4-1:0] node9759;
	wire [4-1:0] node9761;
	wire [4-1:0] node9763;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9769;
	wire [4-1:0] node9770;
	wire [4-1:0] node9774;
	wire [4-1:0] node9776;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9786;
	wire [4-1:0] node9787;
	wire [4-1:0] node9788;
	wire [4-1:0] node9789;
	wire [4-1:0] node9790;
	wire [4-1:0] node9796;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9805;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9813;
	wire [4-1:0] node9814;
	wire [4-1:0] node9815;
	wire [4-1:0] node9816;
	wire [4-1:0] node9817;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9824;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9830;
	wire [4-1:0] node9833;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9859;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9864;
	wire [4-1:0] node9867;
	wire [4-1:0] node9868;
	wire [4-1:0] node9869;
	wire [4-1:0] node9872;
	wire [4-1:0] node9876;
	wire [4-1:0] node9877;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9886;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9894;
	wire [4-1:0] node9897;
	wire [4-1:0] node9898;
	wire [4-1:0] node9899;
	wire [4-1:0] node9901;
	wire [4-1:0] node9904;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9910;
	wire [4-1:0] node9914;
	wire [4-1:0] node9915;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9918;
	wire [4-1:0] node9919;
	wire [4-1:0] node9921;
	wire [4-1:0] node9923;
	wire [4-1:0] node9926;
	wire [4-1:0] node9927;
	wire [4-1:0] node9931;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9936;
	wire [4-1:0] node9938;
	wire [4-1:0] node9941;
	wire [4-1:0] node9942;
	wire [4-1:0] node9945;
	wire [4-1:0] node9947;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9954;
	wire [4-1:0] node9957;
	wire [4-1:0] node9958;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9968;
	wire [4-1:0] node9970;
	wire [4-1:0] node9973;
	wire [4-1:0] node9974;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9978;
	wire [4-1:0] node9981;
	wire [4-1:0] node9982;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9992;
	wire [4-1:0] node9994;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10001;
	wire [4-1:0] node10004;
	wire [4-1:0] node10006;
	wire [4-1:0] node10008;
	wire [4-1:0] node10011;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10017;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10025;
	wire [4-1:0] node10026;
	wire [4-1:0] node10028;
	wire [4-1:0] node10031;
	wire [4-1:0] node10034;
	wire [4-1:0] node10035;
	wire [4-1:0] node10036;
	wire [4-1:0] node10037;
	wire [4-1:0] node10043;
	wire [4-1:0] node10044;
	wire [4-1:0] node10045;
	wire [4-1:0] node10047;
	wire [4-1:0] node10050;
	wire [4-1:0] node10051;
	wire [4-1:0] node10052;
	wire [4-1:0] node10056;
	wire [4-1:0] node10059;
	wire [4-1:0] node10060;
	wire [4-1:0] node10062;
	wire [4-1:0] node10065;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10072;
	wire [4-1:0] node10073;
	wire [4-1:0] node10074;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10080;
	wire [4-1:0] node10084;
	wire [4-1:0] node10085;
	wire [4-1:0] node10086;
	wire [4-1:0] node10089;
	wire [4-1:0] node10093;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10097;
	wire [4-1:0] node10100;
	wire [4-1:0] node10103;
	wire [4-1:0] node10104;
	wire [4-1:0] node10107;
	wire [4-1:0] node10109;
	wire [4-1:0] node10112;
	wire [4-1:0] node10113;
	wire [4-1:0] node10114;
	wire [4-1:0] node10115;
	wire [4-1:0] node10119;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10125;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10132;
	wire [4-1:0] node10133;
	wire [4-1:0] node10134;
	wire [4-1:0] node10135;
	wire [4-1:0] node10136;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10145;
	wire [4-1:0] node10148;
	wire [4-1:0] node10151;
	wire [4-1:0] node10153;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10161;
	wire [4-1:0] node10162;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10169;
	wire [4-1:0] node10172;
	wire [4-1:0] node10173;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10185;
	wire [4-1:0] node10186;
	wire [4-1:0] node10187;
	wire [4-1:0] node10190;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10203;
	wire [4-1:0] node10206;
	wire [4-1:0] node10209;
	wire [4-1:0] node10210;
	wire [4-1:0] node10213;
	wire [4-1:0] node10215;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10223;
	wire [4-1:0] node10227;
	wire [4-1:0] node10228;
	wire [4-1:0] node10231;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10242;
	wire [4-1:0] node10243;
	wire [4-1:0] node10245;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10251;
	wire [4-1:0] node10252;
	wire [4-1:0] node10255;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10262;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10267;
	wire [4-1:0] node10270;
	wire [4-1:0] node10273;
	wire [4-1:0] node10275;
	wire [4-1:0] node10277;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10288;
	wire [4-1:0] node10291;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10296;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10303;
	wire [4-1:0] node10306;
	wire [4-1:0] node10307;
	wire [4-1:0] node10309;
	wire [4-1:0] node10312;
	wire [4-1:0] node10314;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10325;
	wire [4-1:0] node10327;
	wire [4-1:0] node10328;
	wire [4-1:0] node10332;
	wire [4-1:0] node10333;
	wire [4-1:0] node10336;
	wire [4-1:0] node10337;
	wire [4-1:0] node10341;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10348;
	wire [4-1:0] node10349;
	wire [4-1:0] node10351;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10360;
	wire [4-1:0] node10363;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10369;
	wire [4-1:0] node10370;
	wire [4-1:0] node10374;
	wire [4-1:0] node10378;
	wire [4-1:0] node10380;
	wire [4-1:0] node10381;
	wire [4-1:0] node10382;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10389;
	wire [4-1:0] node10390;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10396;
	wire [4-1:0] node10397;
	wire [4-1:0] node10400;
	wire [4-1:0] node10402;
	wire [4-1:0] node10405;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10418;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10434;
	wire [4-1:0] node10438;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10443;
	wire [4-1:0] node10446;
	wire [4-1:0] node10449;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10454;
	wire [4-1:0] node10457;
	wire [4-1:0] node10459;
	wire [4-1:0] node10460;
	wire [4-1:0] node10463;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10468;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10472;
	wire [4-1:0] node10473;
	wire [4-1:0] node10474;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10480;
	wire [4-1:0] node10483;
	wire [4-1:0] node10484;
	wire [4-1:0] node10487;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10496;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10502;
	wire [4-1:0] node10506;
	wire [4-1:0] node10509;
	wire [4-1:0] node10510;
	wire [4-1:0] node10512;
	wire [4-1:0] node10515;
	wire [4-1:0] node10516;
	wire [4-1:0] node10520;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10526;
	wire [4-1:0] node10528;
	wire [4-1:0] node10530;
	wire [4-1:0] node10533;
	wire [4-1:0] node10534;
	wire [4-1:0] node10537;
	wire [4-1:0] node10539;
	wire [4-1:0] node10540;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10546;
	wire [4-1:0] node10547;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10554;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10563;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10572;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10577;
	wire [4-1:0] node10578;
	wire [4-1:0] node10579;
	wire [4-1:0] node10582;
	wire [4-1:0] node10584;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10590;
	wire [4-1:0] node10592;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10599;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10605;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10616;
	wire [4-1:0] node10618;
	wire [4-1:0] node10619;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10625;
	wire [4-1:0] node10626;
	wire [4-1:0] node10627;
	wire [4-1:0] node10630;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10637;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10645;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10657;
	wire [4-1:0] node10660;
	wire [4-1:0] node10663;
	wire [4-1:0] node10666;
	wire [4-1:0] node10667;
	wire [4-1:0] node10668;
	wire [4-1:0] node10669;
	wire [4-1:0] node10670;
	wire [4-1:0] node10671;
	wire [4-1:0] node10672;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10682;
	wire [4-1:0] node10684;
	wire [4-1:0] node10687;
	wire [4-1:0] node10688;
	wire [4-1:0] node10689;
	wire [4-1:0] node10691;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10702;
	wire [4-1:0] node10703;
	wire [4-1:0] node10704;
	wire [4-1:0] node10707;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10713;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10724;
	wire [4-1:0] node10728;
	wire [4-1:0] node10729;
	wire [4-1:0] node10732;
	wire [4-1:0] node10735;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10738;
	wire [4-1:0] node10739;
	wire [4-1:0] node10740;
	wire [4-1:0] node10743;
	wire [4-1:0] node10746;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10753;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10763;
	wire [4-1:0] node10764;
	wire [4-1:0] node10766;
	wire [4-1:0] node10769;
	wire [4-1:0] node10770;
	wire [4-1:0] node10773;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10786;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10793;
	wire [4-1:0] node10797;
	wire [4-1:0] node10800;
	wire [4-1:0] node10802;
	wire [4-1:0] node10803;
	wire [4-1:0] node10804;
	wire [4-1:0] node10808;
	wire [4-1:0] node10811;
	wire [4-1:0] node10812;
	wire [4-1:0] node10813;
	wire [4-1:0] node10815;
	wire [4-1:0] node10816;
	wire [4-1:0] node10820;
	wire [4-1:0] node10823;
	wire [4-1:0] node10824;
	wire [4-1:0] node10825;
	wire [4-1:0] node10828;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10834;
	wire [4-1:0] node10837;
	wire [4-1:0] node10840;
	wire [4-1:0] node10841;
	wire [4-1:0] node10842;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10847;
	wire [4-1:0] node10850;
	wire [4-1:0] node10853;
	wire [4-1:0] node10854;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10860;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10867;
	wire [4-1:0] node10868;
	wire [4-1:0] node10872;
	wire [4-1:0] node10873;
	wire [4-1:0] node10874;
	wire [4-1:0] node10877;
	wire [4-1:0] node10878;
	wire [4-1:0] node10881;
	wire [4-1:0] node10884;
	wire [4-1:0] node10885;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10891;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10898;
	wire [4-1:0] node10900;
	wire [4-1:0] node10903;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10907;
	wire [4-1:0] node10908;
	wire [4-1:0] node10909;
	wire [4-1:0] node10911;
	wire [4-1:0] node10912;
	wire [4-1:0] node10916;
	wire [4-1:0] node10917;
	wire [4-1:0] node10918;
	wire [4-1:0] node10922;
	wire [4-1:0] node10925;
	wire [4-1:0] node10926;
	wire [4-1:0] node10927;
	wire [4-1:0] node10931;
	wire [4-1:0] node10933;
	wire [4-1:0] node10936;
	wire [4-1:0] node10937;
	wire [4-1:0] node10938;
	wire [4-1:0] node10939;
	wire [4-1:0] node10942;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10949;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10954;
	wire [4-1:0] node10957;
	wire [4-1:0] node10960;
	wire [4-1:0] node10962;
	wire [4-1:0] node10963;
	wire [4-1:0] node10967;
	wire [4-1:0] node10968;
	wire [4-1:0] node10969;
	wire [4-1:0] node10970;
	wire [4-1:0] node10971;
	wire [4-1:0] node10973;
	wire [4-1:0] node10977;
	wire [4-1:0] node10979;
	wire [4-1:0] node10982;
	wire [4-1:0] node10983;
	wire [4-1:0] node10985;
	wire [4-1:0] node10987;
	wire [4-1:0] node10990;
	wire [4-1:0] node10991;
	wire [4-1:0] node10992;
	wire [4-1:0] node10995;
	wire [4-1:0] node10998;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11003;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11010;
	wire [4-1:0] node11012;
	wire [4-1:0] node11013;
	wire [4-1:0] node11017;
	wire [4-1:0] node11018;
	wire [4-1:0] node11021;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11027;
	wire [4-1:0] node11028;
	wire [4-1:0] node11031;
	wire [4-1:0] node11032;
	wire [4-1:0] node11033;
	wire [4-1:0] node11036;
	wire [4-1:0] node11040;
	wire [4-1:0] node11041;
	wire [4-1:0] node11043;
	wire [4-1:0] node11044;
	wire [4-1:0] node11048;
	wire [4-1:0] node11049;
	wire [4-1:0] node11051;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11057;
	wire [4-1:0] node11058;
	wire [4-1:0] node11059;
	wire [4-1:0] node11063;
	wire [4-1:0] node11065;
	wire [4-1:0] node11068;
	wire [4-1:0] node11071;
	wire [4-1:0] node11073;
	wire [4-1:0] node11076;
	wire [4-1:0] node11077;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11080;
	wire [4-1:0] node11084;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11094;
	wire [4-1:0] node11095;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11103;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11108;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11113;
	wire [4-1:0] node11118;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11122;
	wire [4-1:0] node11125;
	wire [4-1:0] node11128;
	wire [4-1:0] node11130;
	wire [4-1:0] node11132;
	wire [4-1:0] node11135;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11139;
	wire [4-1:0] node11141;
	wire [4-1:0] node11142;
	wire [4-1:0] node11145;
	wire [4-1:0] node11148;
	wire [4-1:0] node11149;
	wire [4-1:0] node11150;
	wire [4-1:0] node11153;
	wire [4-1:0] node11156;
	wire [4-1:0] node11158;
	wire [4-1:0] node11160;
	wire [4-1:0] node11163;
	wire [4-1:0] node11164;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11170;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11176;
	wire [4-1:0] node11179;
	wire [4-1:0] node11180;
	wire [4-1:0] node11182;
	wire [4-1:0] node11185;
	wire [4-1:0] node11188;
	wire [4-1:0] node11189;
	wire [4-1:0] node11190;
	wire [4-1:0] node11191;
	wire [4-1:0] node11192;
	wire [4-1:0] node11195;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11203;
	wire [4-1:0] node11205;
	wire [4-1:0] node11208;
	wire [4-1:0] node11209;
	wire [4-1:0] node11210;
	wire [4-1:0] node11212;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11218;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11225;
	wire [4-1:0] node11226;
	wire [4-1:0] node11227;
	wire [4-1:0] node11230;
	wire [4-1:0] node11232;
	wire [4-1:0] node11235;
	wire [4-1:0] node11236;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11246;
	wire [4-1:0] node11247;
	wire [4-1:0] node11248;
	wire [4-1:0] node11253;
	wire [4-1:0] node11254;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11262;
	wire [4-1:0] node11263;
	wire [4-1:0] node11266;
	wire [4-1:0] node11268;
	wire [4-1:0] node11271;
	wire [4-1:0] node11272;
	wire [4-1:0] node11274;
	wire [4-1:0] node11275;
	wire [4-1:0] node11279;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11284;
	wire [4-1:0] node11285;
	wire [4-1:0] node11286;
	wire [4-1:0] node11287;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11294;
	wire [4-1:0] node11295;
	wire [4-1:0] node11298;
	wire [4-1:0] node11300;
	wire [4-1:0] node11303;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11309;
	wire [4-1:0] node11312;
	wire [4-1:0] node11313;
	wire [4-1:0] node11317;
	wire [4-1:0] node11318;
	wire [4-1:0] node11320;
	wire [4-1:0] node11323;
	wire [4-1:0] node11326;
	wire [4-1:0] node11327;
	wire [4-1:0] node11328;
	wire [4-1:0] node11329;
	wire [4-1:0] node11333;
	wire [4-1:0] node11335;
	wire [4-1:0] node11337;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11346;
	wire [4-1:0] node11349;
	wire [4-1:0] node11352;
	wire [4-1:0] node11354;
	wire [4-1:0] node11357;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11361;
	wire [4-1:0] node11364;
	wire [4-1:0] node11367;
	wire [4-1:0] node11368;
	wire [4-1:0] node11372;
	wire [4-1:0] node11373;
	wire [4-1:0] node11376;
	wire [4-1:0] node11377;
	wire [4-1:0] node11380;
	wire [4-1:0] node11383;
	wire [4-1:0] node11384;
	wire [4-1:0] node11385;
	wire [4-1:0] node11388;
	wire [4-1:0] node11391;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11394;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11403;
	wire [4-1:0] node11406;
	wire [4-1:0] node11407;
	wire [4-1:0] node11408;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11411;
	wire [4-1:0] node11413;
	wire [4-1:0] node11416;
	wire [4-1:0] node11419;
	wire [4-1:0] node11420;
	wire [4-1:0] node11421;
	wire [4-1:0] node11425;
	wire [4-1:0] node11426;
	wire [4-1:0] node11429;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11438;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11448;
	wire [4-1:0] node11451;
	wire [4-1:0] node11452;
	wire [4-1:0] node11455;
	wire [4-1:0] node11458;
	wire [4-1:0] node11461;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11469;
	wire [4-1:0] node11472;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11479;
	wire [4-1:0] node11482;
	wire [4-1:0] node11483;
	wire [4-1:0] node11484;
	wire [4-1:0] node11485;
	wire [4-1:0] node11486;
	wire [4-1:0] node11488;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11496;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11501;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11509;
	wire [4-1:0] node11511;
	wire [4-1:0] node11514;
	wire [4-1:0] node11515;
	wire [4-1:0] node11516;
	wire [4-1:0] node11517;
	wire [4-1:0] node11518;
	wire [4-1:0] node11523;
	wire [4-1:0] node11526;
	wire [4-1:0] node11527;
	wire [4-1:0] node11530;
	wire [4-1:0] node11531;
	wire [4-1:0] node11534;
	wire [4-1:0] node11536;
	wire [4-1:0] node11539;
	wire [4-1:0] node11540;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11545;
	wire [4-1:0] node11549;
	wire [4-1:0] node11550;
	wire [4-1:0] node11553;
	wire [4-1:0] node11556;
	wire [4-1:0] node11557;
	wire [4-1:0] node11558;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11566;
	wire [4-1:0] node11567;
	wire [4-1:0] node11569;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11577;
	wire [4-1:0] node11578;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11583;
	wire [4-1:0] node11587;
	wire [4-1:0] node11588;
	wire [4-1:0] node11590;
	wire [4-1:0] node11591;
	wire [4-1:0] node11595;
	wire [4-1:0] node11596;
	wire [4-1:0] node11599;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11608;
	wire [4-1:0] node11609;
	wire [4-1:0] node11610;
	wire [4-1:0] node11615;
	wire [4-1:0] node11617;
	wire [4-1:0] node11620;
	wire [4-1:0] node11621;
	wire [4-1:0] node11622;
	wire [4-1:0] node11623;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11630;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11639;
	wire [4-1:0] node11640;
	wire [4-1:0] node11644;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11651;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11657;
	wire [4-1:0] node11658;
	wire [4-1:0] node11661;
	wire [4-1:0] node11665;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11671;
	wire [4-1:0] node11672;
	wire [4-1:0] node11675;
	wire [4-1:0] node11678;
	wire [4-1:0] node11679;
	wire [4-1:0] node11680;
	wire [4-1:0] node11681;
	wire [4-1:0] node11683;
	wire [4-1:0] node11686;
	wire [4-1:0] node11689;
	wire [4-1:0] node11691;
	wire [4-1:0] node11694;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11700;
	wire [4-1:0] node11701;
	wire [4-1:0] node11703;
	wire [4-1:0] node11706;
	wire [4-1:0] node11709;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11714;
	wire [4-1:0] node11720;
	wire [4-1:0] node11721;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11728;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11734;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11740;
	wire [4-1:0] node11743;
	wire [4-1:0] node11747;
	wire [4-1:0] node11748;
	wire [4-1:0] node11749;
	wire [4-1:0] node11754;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11759;
	wire [4-1:0] node11760;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11767;
	wire [4-1:0] node11770;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11776;
	wire [4-1:0] node11778;
	wire [4-1:0] node11781;
	wire [4-1:0] node11782;
	wire [4-1:0] node11783;
	wire [4-1:0] node11784;
	wire [4-1:0] node11787;
	wire [4-1:0] node11790;
	wire [4-1:0] node11792;
	wire [4-1:0] node11795;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11800;
	wire [4-1:0] node11803;
	wire [4-1:0] node11805;
	wire [4-1:0] node11808;
	wire [4-1:0] node11809;
	wire [4-1:0] node11810;
	wire [4-1:0] node11811;
	wire [4-1:0] node11812;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11820;
	wire [4-1:0] node11822;
	wire [4-1:0] node11825;
	wire [4-1:0] node11827;
	wire [4-1:0] node11828;
	wire [4-1:0] node11832;
	wire [4-1:0] node11833;
	wire [4-1:0] node11834;
	wire [4-1:0] node11836;
	wire [4-1:0] node11839;
	wire [4-1:0] node11842;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11846;
	wire [4-1:0] node11850;
	wire [4-1:0] node11853;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11858;
	wire [4-1:0] node11862;
	wire [4-1:0] node11864;
	wire [4-1:0] node11867;
	wire [4-1:0] node11868;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11874;
	wire [4-1:0] node11877;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11885;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11890;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11899;
	wire [4-1:0] node11900;
	wire [4-1:0] node11902;
	wire [4-1:0] node11904;
	wire [4-1:0] node11905;
	wire [4-1:0] node11906;
	wire [4-1:0] node11910;
	wire [4-1:0] node11913;
	wire [4-1:0] node11914;
	wire [4-1:0] node11915;
	wire [4-1:0] node11917;
	wire [4-1:0] node11920;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11927;
	wire [4-1:0] node11928;
	wire [4-1:0] node11931;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11936;
	wire [4-1:0] node11937;
	wire [4-1:0] node11938;
	wire [4-1:0] node11939;
	wire [4-1:0] node11943;
	wire [4-1:0] node11945;
	wire [4-1:0] node11946;
	wire [4-1:0] node11950;
	wire [4-1:0] node11951;
	wire [4-1:0] node11952;
	wire [4-1:0] node11953;
	wire [4-1:0] node11955;
	wire [4-1:0] node11959;
	wire [4-1:0] node11961;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11976;
	wire [4-1:0] node11979;
	wire [4-1:0] node11981;
	wire [4-1:0] node11984;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11988;
	wire [4-1:0] node11991;
	wire [4-1:0] node11994;
	wire [4-1:0] node11996;
	wire [4-1:0] node11999;
	wire [4-1:0] node12000;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12012;
	wire [4-1:0] node12015;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12020;
	wire [4-1:0] node12024;
	wire [4-1:0] node12025;
	wire [4-1:0] node12026;
	wire [4-1:0] node12027;
	wire [4-1:0] node12029;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12034;
	wire [4-1:0] node12037;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12043;
	wire [4-1:0] node12046;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12055;
	wire [4-1:0] node12058;
	wire [4-1:0] node12059;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12065;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12070;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12078;
	wire [4-1:0] node12080;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12091;
	wire [4-1:0] node12092;
	wire [4-1:0] node12093;
	wire [4-1:0] node12094;
	wire [4-1:0] node12095;
	wire [4-1:0] node12098;
	wire [4-1:0] node12099;
	wire [4-1:0] node12103;
	wire [4-1:0] node12106;
	wire [4-1:0] node12107;
	wire [4-1:0] node12108;
	wire [4-1:0] node12111;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12117;
	wire [4-1:0] node12119;
	wire [4-1:0] node12122;
	wire [4-1:0] node12124;
	wire [4-1:0] node12127;
	wire [4-1:0] node12128;
	wire [4-1:0] node12129;
	wire [4-1:0] node12133;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12142;
	wire [4-1:0] node12143;
	wire [4-1:0] node12146;
	wire [4-1:0] node12149;
	wire [4-1:0] node12150;
	wire [4-1:0] node12151;
	wire [4-1:0] node12155;
	wire [4-1:0] node12156;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12163;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12169;
	wire [4-1:0] node12170;
	wire [4-1:0] node12173;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12179;
	wire [4-1:0] node12183;
	wire [4-1:0] node12184;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12187;
	wire [4-1:0] node12190;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12202;
	wire [4-1:0] node12204;
	wire [4-1:0] node12207;
	wire [4-1:0] node12209;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12215;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12228;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12232;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12239;
	wire [4-1:0] node12240;
	wire [4-1:0] node12243;
	wire [4-1:0] node12247;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12253;
	wire [4-1:0] node12255;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12261;
	wire [4-1:0] node12262;
	wire [4-1:0] node12264;
	wire [4-1:0] node12267;
	wire [4-1:0] node12269;
	wire [4-1:0] node12270;
	wire [4-1:0] node12272;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12279;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12285;
	wire [4-1:0] node12286;
	wire [4-1:0] node12290;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12297;
	wire [4-1:0] node12301;
	wire [4-1:0] node12302;
	wire [4-1:0] node12303;
	wire [4-1:0] node12304;
	wire [4-1:0] node12307;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12319;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12325;
	wire [4-1:0] node12326;
	wire [4-1:0] node12330;
	wire [4-1:0] node12331;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12335;
	wire [4-1:0] node12338;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12349;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12356;
	wire [4-1:0] node12359;
	wire [4-1:0] node12360;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12376;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12388;
	wire [4-1:0] node12390;
	wire [4-1:0] node12391;
	wire [4-1:0] node12394;
	wire [4-1:0] node12397;
	wire [4-1:0] node12398;
	wire [4-1:0] node12399;
	wire [4-1:0] node12400;
	wire [4-1:0] node12401;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12406;
	wire [4-1:0] node12409;
	wire [4-1:0] node12411;
	wire [4-1:0] node12414;
	wire [4-1:0] node12417;
	wire [4-1:0] node12419;
	wire [4-1:0] node12422;
	wire [4-1:0] node12423;
	wire [4-1:0] node12424;
	wire [4-1:0] node12426;
	wire [4-1:0] node12429;
	wire [4-1:0] node12432;
	wire [4-1:0] node12433;
	wire [4-1:0] node12434;
	wire [4-1:0] node12436;
	wire [4-1:0] node12439;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12444;
	wire [4-1:0] node12449;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12454;
	wire [4-1:0] node12456;
	wire [4-1:0] node12457;
	wire [4-1:0] node12460;
	wire [4-1:0] node12463;
	wire [4-1:0] node12464;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12473;
	wire [4-1:0] node12476;
	wire [4-1:0] node12478;
	wire [4-1:0] node12481;
	wire [4-1:0] node12483;
	wire [4-1:0] node12484;
	wire [4-1:0] node12487;
	wire [4-1:0] node12489;
	wire [4-1:0] node12492;
	wire [4-1:0] node12493;
	wire [4-1:0] node12494;
	wire [4-1:0] node12495;
	wire [4-1:0] node12496;
	wire [4-1:0] node12498;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12506;
	wire [4-1:0] node12509;
	wire [4-1:0] node12510;
	wire [4-1:0] node12511;
	wire [4-1:0] node12515;
	wire [4-1:0] node12516;
	wire [4-1:0] node12517;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12526;
	wire [4-1:0] node12527;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12532;
	wire [4-1:0] node12535;
	wire [4-1:0] node12536;
	wire [4-1:0] node12540;
	wire [4-1:0] node12542;
	wire [4-1:0] node12545;
	wire [4-1:0] node12546;
	wire [4-1:0] node12547;
	wire [4-1:0] node12550;
	wire [4-1:0] node12553;
	wire [4-1:0] node12554;
	wire [4-1:0] node12557;
	wire [4-1:0] node12560;
	wire [4-1:0] node12561;
	wire [4-1:0] node12563;
	wire [4-1:0] node12566;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12573;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12578;
	wire [4-1:0] node12581;
	wire [4-1:0] node12583;
	wire [4-1:0] node12586;
	wire [4-1:0] node12587;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12594;
	wire [4-1:0] node12597;
	wire [4-1:0] node12599;
	wire [4-1:0] node12600;
	wire [4-1:0] node12604;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12608;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12615;
	wire [4-1:0] node12619;
	wire [4-1:0] node12620;
	wire [4-1:0] node12622;
	wire [4-1:0] node12626;
	wire [4-1:0] node12627;
	wire [4-1:0] node12628;
	wire [4-1:0] node12629;
	wire [4-1:0] node12633;
	wire [4-1:0] node12635;
	wire [4-1:0] node12638;
	wire [4-1:0] node12639;
	wire [4-1:0] node12640;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12649;
	wire [4-1:0] node12650;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12654;
	wire [4-1:0] node12656;
	wire [4-1:0] node12659;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12669;
	wire [4-1:0] node12672;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12676;
	wire [4-1:0] node12679;
	wire [4-1:0] node12681;
	wire [4-1:0] node12684;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12689;
	wire [4-1:0] node12691;
	wire [4-1:0] node12693;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12700;
	wire [4-1:0] node12703;
	wire [4-1:0] node12704;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12716;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12722;
	wire [4-1:0] node12723;
	wire [4-1:0] node12724;
	wire [4-1:0] node12725;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12729;
	wire [4-1:0] node12733;
	wire [4-1:0] node12735;
	wire [4-1:0] node12736;
	wire [4-1:0] node12737;
	wire [4-1:0] node12741;
	wire [4-1:0] node12743;
	wire [4-1:0] node12746;
	wire [4-1:0] node12747;
	wire [4-1:0] node12749;
	wire [4-1:0] node12752;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12758;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12764;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12779;
	wire [4-1:0] node12780;
	wire [4-1:0] node12781;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12790;
	wire [4-1:0] node12791;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12804;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12810;
	wire [4-1:0] node12811;
	wire [4-1:0] node12812;
	wire [4-1:0] node12815;
	wire [4-1:0] node12819;
	wire [4-1:0] node12821;
	wire [4-1:0] node12822;
	wire [4-1:0] node12824;
	wire [4-1:0] node12827;
	wire [4-1:0] node12828;
	wire [4-1:0] node12832;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12836;
	wire [4-1:0] node12839;
	wire [4-1:0] node12842;
	wire [4-1:0] node12844;
	wire [4-1:0] node12847;
	wire [4-1:0] node12849;
	wire [4-1:0] node12851;
	wire [4-1:0] node12853;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12858;
	wire [4-1:0] node12859;
	wire [4-1:0] node12864;
	wire [4-1:0] node12865;
	wire [4-1:0] node12868;
	wire [4-1:0] node12869;
	wire [4-1:0] node12873;
	wire [4-1:0] node12874;
	wire [4-1:0] node12875;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12881;
	wire [4-1:0] node12884;
	wire [4-1:0] node12885;
	wire [4-1:0] node12889;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12900;
	wire [4-1:0] node12901;
	wire [4-1:0] node12904;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12909;
	wire [4-1:0] node12913;
	wire [4-1:0] node12914;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12922;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12925;
	wire [4-1:0] node12929;
	wire [4-1:0] node12931;
	wire [4-1:0] node12934;
	wire [4-1:0] node12935;
	wire [4-1:0] node12939;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12945;
	wire [4-1:0] node12948;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12951;
	wire [4-1:0] node12955;
	wire [4-1:0] node12956;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12964;
	wire [4-1:0] node12965;
	wire [4-1:0] node12969;
	wire [4-1:0] node12970;
	wire [4-1:0] node12971;
	wire [4-1:0] node12972;
	wire [4-1:0] node12974;
	wire [4-1:0] node12976;
	wire [4-1:0] node12979;
	wire [4-1:0] node12980;
	wire [4-1:0] node12983;
	wire [4-1:0] node12986;
	wire [4-1:0] node12987;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13001;
	wire [4-1:0] node13004;
	wire [4-1:0] node13005;
	wire [4-1:0] node13006;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13013;
	wire [4-1:0] node13016;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13031;
	wire [4-1:0] node13032;
	wire [4-1:0] node13035;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13047;
	wire [4-1:0] node13048;
	wire [4-1:0] node13052;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13055;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13058;
	wire [4-1:0] node13060;
	wire [4-1:0] node13063;
	wire [4-1:0] node13065;
	wire [4-1:0] node13066;
	wire [4-1:0] node13069;
	wire [4-1:0] node13072;
	wire [4-1:0] node13073;
	wire [4-1:0] node13074;
	wire [4-1:0] node13076;
	wire [4-1:0] node13080;
	wire [4-1:0] node13082;
	wire [4-1:0] node13084;
	wire [4-1:0] node13087;
	wire [4-1:0] node13088;
	wire [4-1:0] node13089;
	wire [4-1:0] node13090;
	wire [4-1:0] node13092;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13102;
	wire [4-1:0] node13105;
	wire [4-1:0] node13106;
	wire [4-1:0] node13108;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13116;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13119;
	wire [4-1:0] node13120;
	wire [4-1:0] node13123;
	wire [4-1:0] node13127;
	wire [4-1:0] node13129;
	wire [4-1:0] node13130;
	wire [4-1:0] node13131;
	wire [4-1:0] node13134;
	wire [4-1:0] node13138;
	wire [4-1:0] node13139;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13147;
	wire [4-1:0] node13150;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13156;
	wire [4-1:0] node13157;
	wire [4-1:0] node13158;
	wire [4-1:0] node13160;
	wire [4-1:0] node13162;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13173;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13178;
	wire [4-1:0] node13179;
	wire [4-1:0] node13182;
	wire [4-1:0] node13185;
	wire [4-1:0] node13187;
	wire [4-1:0] node13190;
	wire [4-1:0] node13191;
	wire [4-1:0] node13192;
	wire [4-1:0] node13194;
	wire [4-1:0] node13197;
	wire [4-1:0] node13198;
	wire [4-1:0] node13201;
	wire [4-1:0] node13204;
	wire [4-1:0] node13206;
	wire [4-1:0] node13209;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13213;
	wire [4-1:0] node13214;
	wire [4-1:0] node13218;
	wire [4-1:0] node13220;
	wire [4-1:0] node13221;
	wire [4-1:0] node13225;
	wire [4-1:0] node13226;
	wire [4-1:0] node13227;
	wire [4-1:0] node13229;
	wire [4-1:0] node13231;
	wire [4-1:0] node13235;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13240;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13247;
	wire [4-1:0] node13248;
	wire [4-1:0] node13249;
	wire [4-1:0] node13250;
	wire [4-1:0] node13253;
	wire [4-1:0] node13257;
	wire [4-1:0] node13258;
	wire [4-1:0] node13259;
	wire [4-1:0] node13261;
	wire [4-1:0] node13264;
	wire [4-1:0] node13266;
	wire [4-1:0] node13269;
	wire [4-1:0] node13271;
	wire [4-1:0] node13274;
	wire [4-1:0] node13275;
	wire [4-1:0] node13277;
	wire [4-1:0] node13279;
	wire [4-1:0] node13281;
	wire [4-1:0] node13284;
	wire [4-1:0] node13287;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13291;
	wire [4-1:0] node13294;
	wire [4-1:0] node13296;
	wire [4-1:0] node13297;
	wire [4-1:0] node13301;
	wire [4-1:0] node13302;
	wire [4-1:0] node13304;
	wire [4-1:0] node13306;
	wire [4-1:0] node13309;
	wire [4-1:0] node13312;
	wire [4-1:0] node13313;
	wire [4-1:0] node13314;
	wire [4-1:0] node13315;
	wire [4-1:0] node13316;
	wire [4-1:0] node13318;
	wire [4-1:0] node13321;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13327;
	wire [4-1:0] node13329;
	wire [4-1:0] node13330;
	wire [4-1:0] node13333;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13340;
	wire [4-1:0] node13344;
	wire [4-1:0] node13347;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13353;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13358;
	wire [4-1:0] node13359;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13365;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13371;
	wire [4-1:0] node13376;
	wire [4-1:0] node13377;
	wire [4-1:0] node13380;
	wire [4-1:0] node13381;
	wire [4-1:0] node13385;
	wire [4-1:0] node13386;
	wire [4-1:0] node13387;
	wire [4-1:0] node13388;
	wire [4-1:0] node13389;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13394;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13405;
	wire [4-1:0] node13407;
	wire [4-1:0] node13410;
	wire [4-1:0] node13411;
	wire [4-1:0] node13416;
	wire [4-1:0] node13418;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13425;
	wire [4-1:0] node13426;
	wire [4-1:0] node13429;
	wire [4-1:0] node13432;
	wire [4-1:0] node13434;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13440;
	wire [4-1:0] node13441;
	wire [4-1:0] node13444;
	wire [4-1:0] node13447;
	wire [4-1:0] node13449;
	wire [4-1:0] node13450;
	wire [4-1:0] node13454;
	wire [4-1:0] node13455;
	wire [4-1:0] node13456;
	wire [4-1:0] node13457;
	wire [4-1:0] node13458;
	wire [4-1:0] node13461;
	wire [4-1:0] node13464;
	wire [4-1:0] node13465;
	wire [4-1:0] node13469;
	wire [4-1:0] node13470;
	wire [4-1:0] node13471;
	wire [4-1:0] node13472;
	wire [4-1:0] node13474;
	wire [4-1:0] node13477;
	wire [4-1:0] node13481;
	wire [4-1:0] node13483;
	wire [4-1:0] node13485;
	wire [4-1:0] node13486;
	wire [4-1:0] node13490;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13494;
	wire [4-1:0] node13496;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13502;
	wire [4-1:0] node13505;
	wire [4-1:0] node13506;
	wire [4-1:0] node13510;
	wire [4-1:0] node13511;
	wire [4-1:0] node13514;
	wire [4-1:0] node13516;
	wire [4-1:0] node13519;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13524;
	wire [4-1:0] node13525;
	wire [4-1:0] node13527;
	wire [4-1:0] node13530;
	wire [4-1:0] node13532;
	wire [4-1:0] node13533;
	wire [4-1:0] node13537;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13545;
	wire [4-1:0] node13546;
	wire [4-1:0] node13547;
	wire [4-1:0] node13552;
	wire [4-1:0] node13553;
	wire [4-1:0] node13554;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13564;
	wire [4-1:0] node13568;
	wire [4-1:0] node13569;
	wire [4-1:0] node13571;
	wire [4-1:0] node13572;
	wire [4-1:0] node13573;
	wire [4-1:0] node13576;
	wire [4-1:0] node13579;
	wire [4-1:0] node13580;
	wire [4-1:0] node13584;
	wire [4-1:0] node13585;
	wire [4-1:0] node13587;
	wire [4-1:0] node13590;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13598;
	wire [4-1:0] node13600;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13609;
	wire [4-1:0] node13610;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13616;
	wire [4-1:0] node13619;
	wire [4-1:0] node13622;
	wire [4-1:0] node13623;
	wire [4-1:0] node13627;
	wire [4-1:0] node13628;
	wire [4-1:0] node13629;
	wire [4-1:0] node13631;
	wire [4-1:0] node13632;
	wire [4-1:0] node13633;
	wire [4-1:0] node13637;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13644;
	wire [4-1:0] node13647;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13652;
	wire [4-1:0] node13656;
	wire [4-1:0] node13657;
	wire [4-1:0] node13658;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13661;
	wire [4-1:0] node13663;
	wire [4-1:0] node13665;
	wire [4-1:0] node13667;
	wire [4-1:0] node13670;
	wire [4-1:0] node13671;
	wire [4-1:0] node13675;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13682;
	wire [4-1:0] node13683;
	wire [4-1:0] node13687;
	wire [4-1:0] node13689;
	wire [4-1:0] node13692;
	wire [4-1:0] node13693;
	wire [4-1:0] node13694;
	wire [4-1:0] node13695;
	wire [4-1:0] node13696;
	wire [4-1:0] node13697;
	wire [4-1:0] node13700;
	wire [4-1:0] node13705;
	wire [4-1:0] node13706;
	wire [4-1:0] node13708;
	wire [4-1:0] node13710;
	wire [4-1:0] node13713;
	wire [4-1:0] node13716;
	wire [4-1:0] node13717;
	wire [4-1:0] node13719;
	wire [4-1:0] node13720;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13726;
	wire [4-1:0] node13728;
	wire [4-1:0] node13731;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13737;
	wire [4-1:0] node13738;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13748;
	wire [4-1:0] node13750;
	wire [4-1:0] node13753;
	wire [4-1:0] node13755;
	wire [4-1:0] node13758;
	wire [4-1:0] node13760;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13766;
	wire [4-1:0] node13767;
	wire [4-1:0] node13768;
	wire [4-1:0] node13773;
	wire [4-1:0] node13774;
	wire [4-1:0] node13775;
	wire [4-1:0] node13779;
	wire [4-1:0] node13780;
	wire [4-1:0] node13782;
	wire [4-1:0] node13785;
	wire [4-1:0] node13786;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13797;
	wire [4-1:0] node13799;
	wire [4-1:0] node13802;
	wire [4-1:0] node13805;
	wire [4-1:0] node13807;
	wire [4-1:0] node13808;
	wire [4-1:0] node13812;
	wire [4-1:0] node13813;
	wire [4-1:0] node13814;
	wire [4-1:0] node13815;
	wire [4-1:0] node13819;
	wire [4-1:0] node13822;
	wire [4-1:0] node13823;
	wire [4-1:0] node13824;
	wire [4-1:0] node13828;
	wire [4-1:0] node13831;
	wire [4-1:0] node13832;
	wire [4-1:0] node13833;
	wire [4-1:0] node13834;
	wire [4-1:0] node13836;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13844;
	wire [4-1:0] node13846;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13856;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13863;
	wire [4-1:0] node13864;
	wire [4-1:0] node13865;
	wire [4-1:0] node13867;
	wire [4-1:0] node13870;
	wire [4-1:0] node13874;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13878;
	wire [4-1:0] node13880;
	wire [4-1:0] node13883;
	wire [4-1:0] node13884;
	wire [4-1:0] node13885;
	wire [4-1:0] node13888;
	wire [4-1:0] node13892;
	wire [4-1:0] node13894;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13899;
	wire [4-1:0] node13901;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13907;
	wire [4-1:0] node13910;
	wire [4-1:0] node13914;
	wire [4-1:0] node13915;
	wire [4-1:0] node13916;
	wire [4-1:0] node13917;
	wire [4-1:0] node13919;
	wire [4-1:0] node13923;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13934;
	wire [4-1:0] node13935;
	wire [4-1:0] node13936;
	wire [4-1:0] node13939;
	wire [4-1:0] node13943;
	wire [4-1:0] node13944;
	wire [4-1:0] node13947;
	wire [4-1:0] node13950;
	wire [4-1:0] node13951;
	wire [4-1:0] node13952;
	wire [4-1:0] node13955;
	wire [4-1:0] node13958;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13965;
	wire [4-1:0] node13966;
	wire [4-1:0] node13967;
	wire [4-1:0] node13968;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13971;
	wire [4-1:0] node13972;
	wire [4-1:0] node13973;
	wire [4-1:0] node13974;
	wire [4-1:0] node13978;
	wire [4-1:0] node13980;
	wire [4-1:0] node13984;
	wire [4-1:0] node13985;
	wire [4-1:0] node13987;
	wire [4-1:0] node13989;
	wire [4-1:0] node13992;
	wire [4-1:0] node13994;
	wire [4-1:0] node13995;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14004;
	wire [4-1:0] node14008;
	wire [4-1:0] node14009;
	wire [4-1:0] node14010;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14014;
	wire [4-1:0] node14018;
	wire [4-1:0] node14021;
	wire [4-1:0] node14022;
	wire [4-1:0] node14023;
	wire [4-1:0] node14027;
	wire [4-1:0] node14028;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14037;
	wire [4-1:0] node14040;
	wire [4-1:0] node14042;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14047;
	wire [4-1:0] node14048;
	wire [4-1:0] node14049;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14055;
	wire [4-1:0] node14058;
	wire [4-1:0] node14060;
	wire [4-1:0] node14064;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14069;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14075;
	wire [4-1:0] node14076;
	wire [4-1:0] node14077;
	wire [4-1:0] node14080;
	wire [4-1:0] node14083;
	wire [4-1:0] node14084;
	wire [4-1:0] node14089;
	wire [4-1:0] node14090;
	wire [4-1:0] node14091;
	wire [4-1:0] node14094;
	wire [4-1:0] node14098;
	wire [4-1:0] node14099;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14102;
	wire [4-1:0] node14103;
	wire [4-1:0] node14106;
	wire [4-1:0] node14108;
	wire [4-1:0] node14111;
	wire [4-1:0] node14113;
	wire [4-1:0] node14115;
	wire [4-1:0] node14118;
	wire [4-1:0] node14119;
	wire [4-1:0] node14120;
	wire [4-1:0] node14121;
	wire [4-1:0] node14122;
	wire [4-1:0] node14127;
	wire [4-1:0] node14129;
	wire [4-1:0] node14131;
	wire [4-1:0] node14134;
	wire [4-1:0] node14136;
	wire [4-1:0] node14139;
	wire [4-1:0] node14140;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14145;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14150;
	wire [4-1:0] node14154;
	wire [4-1:0] node14155;
	wire [4-1:0] node14158;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14169;
	wire [4-1:0] node14170;
	wire [4-1:0] node14171;
	wire [4-1:0] node14172;
	wire [4-1:0] node14175;
	wire [4-1:0] node14179;
	wire [4-1:0] node14180;
	wire [4-1:0] node14183;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14188;
	wire [4-1:0] node14189;
	wire [4-1:0] node14191;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14202;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14212;
	wire [4-1:0] node14213;
	wire [4-1:0] node14217;
	wire [4-1:0] node14218;
	wire [4-1:0] node14222;
	wire [4-1:0] node14223;
	wire [4-1:0] node14224;
	wire [4-1:0] node14227;
	wire [4-1:0] node14228;
	wire [4-1:0] node14231;
	wire [4-1:0] node14234;
	wire [4-1:0] node14235;
	wire [4-1:0] node14236;
	wire [4-1:0] node14239;
	wire [4-1:0] node14242;
	wire [4-1:0] node14243;
	wire [4-1:0] node14245;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14251;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14255;
	wire [4-1:0] node14258;
	wire [4-1:0] node14259;
	wire [4-1:0] node14262;
	wire [4-1:0] node14265;
	wire [4-1:0] node14267;
	wire [4-1:0] node14269;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14274;
	wire [4-1:0] node14277;
	wire [4-1:0] node14280;
	wire [4-1:0] node14281;
	wire [4-1:0] node14283;
	wire [4-1:0] node14286;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14292;
	wire [4-1:0] node14293;
	wire [4-1:0] node14296;
	wire [4-1:0] node14298;
	wire [4-1:0] node14301;
	wire [4-1:0] node14302;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14310;
	wire [4-1:0] node14312;
	wire [4-1:0] node14313;
	wire [4-1:0] node14316;
	wire [4-1:0] node14318;
	wire [4-1:0] node14321;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14326;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14332;
	wire [4-1:0] node14335;
	wire [4-1:0] node14337;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14343;
	wire [4-1:0] node14344;
	wire [4-1:0] node14345;
	wire [4-1:0] node14346;
	wire [4-1:0] node14350;
	wire [4-1:0] node14352;
	wire [4-1:0] node14356;
	wire [4-1:0] node14357;
	wire [4-1:0] node14359;
	wire [4-1:0] node14363;
	wire [4-1:0] node14364;
	wire [4-1:0] node14366;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14372;
	wire [4-1:0] node14374;
	wire [4-1:0] node14377;
	wire [4-1:0] node14379;
	wire [4-1:0] node14382;
	wire [4-1:0] node14383;
	wire [4-1:0] node14384;
	wire [4-1:0] node14385;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14395;
	wire [4-1:0] node14400;
	wire [4-1:0] node14401;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14407;
	wire [4-1:0] node14410;
	wire [4-1:0] node14411;
	wire [4-1:0] node14412;
	wire [4-1:0] node14415;
	wire [4-1:0] node14418;
	wire [4-1:0] node14420;
	wire [4-1:0] node14421;
	wire [4-1:0] node14424;
	wire [4-1:0] node14427;
	wire [4-1:0] node14428;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14432;
	wire [4-1:0] node14433;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14440;
	wire [4-1:0] node14444;
	wire [4-1:0] node14445;
	wire [4-1:0] node14449;
	wire [4-1:0] node14450;
	wire [4-1:0] node14451;
	wire [4-1:0] node14452;
	wire [4-1:0] node14453;
	wire [4-1:0] node14458;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14466;
	wire [4-1:0] node14467;
	wire [4-1:0] node14468;
	wire [4-1:0] node14469;
	wire [4-1:0] node14470;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14484;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14489;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14496;
	wire [4-1:0] node14499;
	wire [4-1:0] node14501;
	wire [4-1:0] node14504;
	wire [4-1:0] node14505;
	wire [4-1:0] node14506;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14514;
	wire [4-1:0] node14517;
	wire [4-1:0] node14518;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14522;
	wire [4-1:0] node14525;
	wire [4-1:0] node14526;
	wire [4-1:0] node14527;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14534;
	wire [4-1:0] node14537;
	wire [4-1:0] node14540;
	wire [4-1:0] node14541;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14546;
	wire [4-1:0] node14550;
	wire [4-1:0] node14552;
	wire [4-1:0] node14554;
	wire [4-1:0] node14557;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14573;
	wire [4-1:0] node14576;
	wire [4-1:0] node14577;
	wire [4-1:0] node14581;
	wire [4-1:0] node14582;
	wire [4-1:0] node14583;
	wire [4-1:0] node14584;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14595;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14604;
	wire [4-1:0] node14605;
	wire [4-1:0] node14606;
	wire [4-1:0] node14607;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14614;
	wire [4-1:0] node14617;
	wire [4-1:0] node14619;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14630;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14636;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14644;
	wire [4-1:0] node14645;
	wire [4-1:0] node14647;
	wire [4-1:0] node14650;
	wire [4-1:0] node14652;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14659;
	wire [4-1:0] node14662;
	wire [4-1:0] node14665;
	wire [4-1:0] node14666;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14670;
	wire [4-1:0] node14673;
	wire [4-1:0] node14675;
	wire [4-1:0] node14678;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14683;
	wire [4-1:0] node14684;
	wire [4-1:0] node14688;
	wire [4-1:0] node14689;
	wire [4-1:0] node14693;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14700;
	wire [4-1:0] node14701;
	wire [4-1:0] node14702;
	wire [4-1:0] node14703;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14710;
	wire [4-1:0] node14713;
	wire [4-1:0] node14716;
	wire [4-1:0] node14719;
	wire [4-1:0] node14720;
	wire [4-1:0] node14721;
	wire [4-1:0] node14722;
	wire [4-1:0] node14726;
	wire [4-1:0] node14727;
	wire [4-1:0] node14730;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14737;
	wire [4-1:0] node14740;
	wire [4-1:0] node14741;
	wire [4-1:0] node14742;
	wire [4-1:0] node14743;
	wire [4-1:0] node14746;
	wire [4-1:0] node14749;
	wire [4-1:0] node14750;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14757;
	wire [4-1:0] node14760;
	wire [4-1:0] node14762;
	wire [4-1:0] node14765;
	wire [4-1:0] node14766;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14770;
	wire [4-1:0] node14771;
	wire [4-1:0] node14775;
	wire [4-1:0] node14776;
	wire [4-1:0] node14778;
	wire [4-1:0] node14782;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14787;
	wire [4-1:0] node14788;
	wire [4-1:0] node14792;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14800;
	wire [4-1:0] node14802;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14808;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14814;
	wire [4-1:0] node14818;
	wire [4-1:0] node14821;
	wire [4-1:0] node14823;
	wire [4-1:0] node14824;
	wire [4-1:0] node14827;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14832;
	wire [4-1:0] node14833;
	wire [4-1:0] node14834;
	wire [4-1:0] node14836;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14843;
	wire [4-1:0] node14846;
	wire [4-1:0] node14847;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14853;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14862;
	wire [4-1:0] node14865;
	wire [4-1:0] node14866;
	wire [4-1:0] node14867;
	wire [4-1:0] node14872;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14877;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14884;
	wire [4-1:0] node14889;
	wire [4-1:0] node14890;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14896;
	wire [4-1:0] node14898;
	wire [4-1:0] node14902;
	wire [4-1:0] node14903;
	wire [4-1:0] node14906;
	wire [4-1:0] node14909;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14912;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14918;
	wire [4-1:0] node14921;
	wire [4-1:0] node14923;
	wire [4-1:0] node14926;
	wire [4-1:0] node14928;
	wire [4-1:0] node14930;
	wire [4-1:0] node14933;
	wire [4-1:0] node14934;
	wire [4-1:0] node14935;
	wire [4-1:0] node14936;
	wire [4-1:0] node14939;
	wire [4-1:0] node14942;
	wire [4-1:0] node14944;
	wire [4-1:0] node14947;
	wire [4-1:0] node14948;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14953;
	wire [4-1:0] node14958;
	wire [4-1:0] node14959;
	wire [4-1:0] node14960;
	wire [4-1:0] node14962;
	wire [4-1:0] node14965;
	wire [4-1:0] node14967;
	wire [4-1:0] node14970;
	wire [4-1:0] node14972;
	wire [4-1:0] node14974;
	wire [4-1:0] node14977;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14980;
	wire [4-1:0] node14981;
	wire [4-1:0] node14984;
	wire [4-1:0] node14987;
	wire [4-1:0] node14988;
	wire [4-1:0] node14991;
	wire [4-1:0] node14994;
	wire [4-1:0] node14995;
	wire [4-1:0] node14998;
	wire [4-1:0] node15001;
	wire [4-1:0] node15002;
	wire [4-1:0] node15003;
	wire [4-1:0] node15005;
	wire [4-1:0] node15008;
	wire [4-1:0] node15009;
	wire [4-1:0] node15012;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15019;
	wire [4-1:0] node15022;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15025;
	wire [4-1:0] node15029;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15033;
	wire [4-1:0] node15036;
	wire [4-1:0] node15040;
	wire [4-1:0] node15041;
	wire [4-1:0] node15042;
	wire [4-1:0] node15046;
	wire [4-1:0] node15047;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15056;
	wire [4-1:0] node15059;
	wire [4-1:0] node15061;
	wire [4-1:0] node15064;
	wire [4-1:0] node15065;
	wire [4-1:0] node15068;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15072;
	wire [4-1:0] node15075;
	wire [4-1:0] node15076;
	wire [4-1:0] node15079;
	wire [4-1:0] node15082;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15088;
	wire [4-1:0] node15091;
	wire [4-1:0] node15092;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15095;
	wire [4-1:0] node15096;
	wire [4-1:0] node15097;
	wire [4-1:0] node15098;
	wire [4-1:0] node15099;
	wire [4-1:0] node15102;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15111;
	wire [4-1:0] node15112;
	wire [4-1:0] node15113;
	wire [4-1:0] node15116;
	wire [4-1:0] node15119;
	wire [4-1:0] node15121;
	wire [4-1:0] node15124;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15130;
	wire [4-1:0] node15131;
	wire [4-1:0] node15132;
	wire [4-1:0] node15133;
	wire [4-1:0] node15137;
	wire [4-1:0] node15138;
	wire [4-1:0] node15142;
	wire [4-1:0] node15143;
	wire [4-1:0] node15146;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15151;
	wire [4-1:0] node15152;
	wire [4-1:0] node15153;
	wire [4-1:0] node15154;
	wire [4-1:0] node15158;
	wire [4-1:0] node15159;
	wire [4-1:0] node15163;
	wire [4-1:0] node15166;
	wire [4-1:0] node15167;
	wire [4-1:0] node15170;
	wire [4-1:0] node15173;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15177;
	wire [4-1:0] node15181;
	wire [4-1:0] node15184;
	wire [4-1:0] node15185;
	wire [4-1:0] node15186;
	wire [4-1:0] node15187;
	wire [4-1:0] node15189;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15196;
	wire [4-1:0] node15199;
	wire [4-1:0] node15200;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15212;
	wire [4-1:0] node15214;
	wire [4-1:0] node15217;
	wire [4-1:0] node15219;
	wire [4-1:0] node15220;
	wire [4-1:0] node15221;
	wire [4-1:0] node15224;
	wire [4-1:0] node15228;
	wire [4-1:0] node15229;
	wire [4-1:0] node15230;
	wire [4-1:0] node15231;
	wire [4-1:0] node15235;
	wire [4-1:0] node15236;
	wire [4-1:0] node15237;
	wire [4-1:0] node15241;
	wire [4-1:0] node15243;
	wire [4-1:0] node15244;
	wire [4-1:0] node15247;
	wire [4-1:0] node15250;
	wire [4-1:0] node15251;
	wire [4-1:0] node15252;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15260;
	wire [4-1:0] node15263;
	wire [4-1:0] node15264;
	wire [4-1:0] node15265;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15268;
	wire [4-1:0] node15271;
	wire [4-1:0] node15274;
	wire [4-1:0] node15276;
	wire [4-1:0] node15278;
	wire [4-1:0] node15281;
	wire [4-1:0] node15282;
	wire [4-1:0] node15283;
	wire [4-1:0] node15286;
	wire [4-1:0] node15289;
	wire [4-1:0] node15290;
	wire [4-1:0] node15291;
	wire [4-1:0] node15295;
	wire [4-1:0] node15297;
	wire [4-1:0] node15298;
	wire [4-1:0] node15301;
	wire [4-1:0] node15304;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15309;
	wire [4-1:0] node15312;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15326;
	wire [4-1:0] node15328;
	wire [4-1:0] node15331;
	wire [4-1:0] node15332;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15339;
	wire [4-1:0] node15342;
	wire [4-1:0] node15345;
	wire [4-1:0] node15346;
	wire [4-1:0] node15350;
	wire [4-1:0] node15351;
	wire [4-1:0] node15354;
	wire [4-1:0] node15357;
	wire [4-1:0] node15358;
	wire [4-1:0] node15361;
	wire [4-1:0] node15364;
	wire [4-1:0] node15365;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15368;
	wire [4-1:0] node15369;
	wire [4-1:0] node15370;
	wire [4-1:0] node15371;
	wire [4-1:0] node15373;
	wire [4-1:0] node15376;
	wire [4-1:0] node15378;
	wire [4-1:0] node15381;
	wire [4-1:0] node15382;
	wire [4-1:0] node15384;
	wire [4-1:0] node15388;
	wire [4-1:0] node15389;
	wire [4-1:0] node15391;
	wire [4-1:0] node15392;
	wire [4-1:0] node15393;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15400;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15407;
	wire [4-1:0] node15408;
	wire [4-1:0] node15412;
	wire [4-1:0] node15414;
	wire [4-1:0] node15415;
	wire [4-1:0] node15417;
	wire [4-1:0] node15420;
	wire [4-1:0] node15422;
	wire [4-1:0] node15425;
	wire [4-1:0] node15426;
	wire [4-1:0] node15427;
	wire [4-1:0] node15428;
	wire [4-1:0] node15429;
	wire [4-1:0] node15433;
	wire [4-1:0] node15434;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15444;
	wire [4-1:0] node15445;
	wire [4-1:0] node15449;
	wire [4-1:0] node15450;
	wire [4-1:0] node15451;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15458;
	wire [4-1:0] node15461;
	wire [4-1:0] node15462;
	wire [4-1:0] node15464;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15471;
	wire [4-1:0] node15472;
	wire [4-1:0] node15473;
	wire [4-1:0] node15476;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15483;
	wire [4-1:0] node15486;
	wire [4-1:0] node15487;
	wire [4-1:0] node15490;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15495;
	wire [4-1:0] node15496;
	wire [4-1:0] node15498;
	wire [4-1:0] node15499;
	wire [4-1:0] node15503;
	wire [4-1:0] node15505;
	wire [4-1:0] node15508;
	wire [4-1:0] node15510;
	wire [4-1:0] node15511;
	wire [4-1:0] node15514;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15525;
	wire [4-1:0] node15526;
	wire [4-1:0] node15528;
	wire [4-1:0] node15529;
	wire [4-1:0] node15532;
	wire [4-1:0] node15535;
	wire [4-1:0] node15537;
	wire [4-1:0] node15540;
	wire [4-1:0] node15541;
	wire [4-1:0] node15542;
	wire [4-1:0] node15543;
	wire [4-1:0] node15544;
	wire [4-1:0] node15548;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15555;
	wire [4-1:0] node15556;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15561;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15575;
	wire [4-1:0] node15578;
	wire [4-1:0] node15579;
	wire [4-1:0] node15580;
	wire [4-1:0] node15582;
	wire [4-1:0] node15585;
	wire [4-1:0] node15587;
	wire [4-1:0] node15588;
	wire [4-1:0] node15589;
	wire [4-1:0] node15594;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15598;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15604;
	wire [4-1:0] node15607;
	wire [4-1:0] node15609;
	wire [4-1:0] node15612;
	wire [4-1:0] node15613;
	wire [4-1:0] node15616;
	wire [4-1:0] node15617;
	wire [4-1:0] node15620;
	wire [4-1:0] node15623;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15626;
	wire [4-1:0] node15629;
	wire [4-1:0] node15632;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15637;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15646;
	wire [4-1:0] node15647;
	wire [4-1:0] node15650;
	wire [4-1:0] node15653;
	wire [4-1:0] node15654;
	wire [4-1:0] node15655;
	wire [4-1:0] node15656;
	wire [4-1:0] node15658;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15665;
	wire [4-1:0] node15668;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15675;
	wire [4-1:0] node15678;
	wire [4-1:0] node15679;
	wire [4-1:0] node15680;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15686;
	wire [4-1:0] node15689;
	wire [4-1:0] node15690;
	wire [4-1:0] node15691;
	wire [4-1:0] node15694;
	wire [4-1:0] node15697;
	wire [4-1:0] node15699;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15705;
	wire [4-1:0] node15708;
	wire [4-1:0] node15712;
	wire [4-1:0] node15713;
	wire [4-1:0] node15715;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15722;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15727;
	wire [4-1:0] node15728;
	wire [4-1:0] node15729;
	wire [4-1:0] node15732;
	wire [4-1:0] node15733;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15738;
	wire [4-1:0] node15743;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15757;
	wire [4-1:0] node15760;
	wire [4-1:0] node15761;
	wire [4-1:0] node15762;
	wire [4-1:0] node15764;
	wire [4-1:0] node15767;
	wire [4-1:0] node15768;
	wire [4-1:0] node15772;
	wire [4-1:0] node15773;
	wire [4-1:0] node15775;
	wire [4-1:0] node15779;
	wire [4-1:0] node15782;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15785;
	wire [4-1:0] node15786;
	wire [4-1:0] node15787;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15793;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15800;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15806;
	wire [4-1:0] node15809;
	wire [4-1:0] node15811;
	wire [4-1:0] node15812;
	wire [4-1:0] node15816;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15822;
	wire [4-1:0] node15823;
	wire [4-1:0] node15826;
	wire [4-1:0] node15829;
	wire [4-1:0] node15830;
	wire [4-1:0] node15831;
	wire [4-1:0] node15832;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15841;
	wire [4-1:0] node15842;
	wire [4-1:0] node15843;
	wire [4-1:0] node15847;
	wire [4-1:0] node15848;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15854;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15860;
	wire [4-1:0] node15862;
	wire [4-1:0] node15865;
	wire [4-1:0] node15866;
	wire [4-1:0] node15867;
	wire [4-1:0] node15868;
	wire [4-1:0] node15872;
	wire [4-1:0] node15875;
	wire [4-1:0] node15876;
	wire [4-1:0] node15879;
	wire [4-1:0] node15882;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15888;
	wire [4-1:0] node15892;
	wire [4-1:0] node15894;
	wire [4-1:0] node15897;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15900;
	wire [4-1:0] node15901;
	wire [4-1:0] node15902;
	wire [4-1:0] node15905;
	wire [4-1:0] node15908;
	wire [4-1:0] node15909;
	wire [4-1:0] node15911;
	wire [4-1:0] node15915;
	wire [4-1:0] node15916;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15924;
	wire [4-1:0] node15927;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15932;
	wire [4-1:0] node15934;
	wire [4-1:0] node15935;
	wire [4-1:0] node15939;
	wire [4-1:0] node15941;
	wire [4-1:0] node15942;
	wire [4-1:0] node15945;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15952;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15958;
	wire [4-1:0] node15959;
	wire [4-1:0] node15960;
	wire [4-1:0] node15963;
	wire [4-1:0] node15966;
	wire [4-1:0] node15968;
	wire [4-1:0] node15971;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15976;
	wire [4-1:0] node15979;
	wire [4-1:0] node15980;
	wire [4-1:0] node15982;
	wire [4-1:0] node15985;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15990;
	wire [4-1:0] node15993;
	wire [4-1:0] node15996;
	wire [4-1:0] node15997;
	wire [4-1:0] node15998;
	wire [4-1:0] node16001;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16011;
	wire [4-1:0] node16014;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16020;
	wire [4-1:0] node16023;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16028;
	wire [4-1:0] node16031;
	wire [4-1:0] node16032;
	wire [4-1:0] node16035;
	wire [4-1:0] node16038;
	wire [4-1:0] node16039;
	wire [4-1:0] node16040;
	wire [4-1:0] node16041;
	wire [4-1:0] node16042;
	wire [4-1:0] node16043;
	wire [4-1:0] node16045;
	wire [4-1:0] node16048;
	wire [4-1:0] node16050;
	wire [4-1:0] node16053;
	wire [4-1:0] node16054;
	wire [4-1:0] node16056;
	wire [4-1:0] node16059;
	wire [4-1:0] node16062;
	wire [4-1:0] node16063;
	wire [4-1:0] node16064;
	wire [4-1:0] node16066;
	wire [4-1:0] node16067;
	wire [4-1:0] node16070;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16079;
	wire [4-1:0] node16081;
	wire [4-1:0] node16084;
	wire [4-1:0] node16085;
	wire [4-1:0] node16086;
	wire [4-1:0] node16089;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16095;
	wire [4-1:0] node16096;
	wire [4-1:0] node16100;
	wire [4-1:0] node16101;
	wire [4-1:0] node16104;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16112;
	wire [4-1:0] node16113;
	wire [4-1:0] node16115;
	wire [4-1:0] node16118;
	wire [4-1:0] node16121;
	wire [4-1:0] node16122;
	wire [4-1:0] node16123;
	wire [4-1:0] node16125;
	wire [4-1:0] node16129;
	wire [4-1:0] node16131;
	wire [4-1:0] node16134;
	wire [4-1:0] node16135;
	wire [4-1:0] node16136;
	wire [4-1:0] node16137;
	wire [4-1:0] node16141;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16151;
	wire [4-1:0] node16152;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16155;
	wire [4-1:0] node16159;
	wire [4-1:0] node16161;
	wire [4-1:0] node16164;
	wire [4-1:0] node16165;
	wire [4-1:0] node16167;
	wire [4-1:0] node16170;
	wire [4-1:0] node16173;
	wire [4-1:0] node16174;
	wire [4-1:0] node16177;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16182;
	wire [4-1:0] node16183;
	wire [4-1:0] node16185;
	wire [4-1:0] node16188;
	wire [4-1:0] node16190;
	wire [4-1:0] node16193;
	wire [4-1:0] node16194;
	wire [4-1:0] node16195;
	wire [4-1:0] node16199;
	wire [4-1:0] node16200;
	wire [4-1:0] node16204;
	wire [4-1:0] node16205;
	wire [4-1:0] node16208;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16214;
	wire [4-1:0] node16215;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16219;
	wire [4-1:0] node16221;
	wire [4-1:0] node16224;
	wire [4-1:0] node16226;
	wire [4-1:0] node16229;
	wire [4-1:0] node16230;
	wire [4-1:0] node16233;
	wire [4-1:0] node16235;
	wire [4-1:0] node16238;
	wire [4-1:0] node16239;
	wire [4-1:0] node16240;
	wire [4-1:0] node16241;
	wire [4-1:0] node16242;
	wire [4-1:0] node16244;
	wire [4-1:0] node16245;
	wire [4-1:0] node16248;
	wire [4-1:0] node16252;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16261;
	wire [4-1:0] node16263;
	wire [4-1:0] node16266;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16275;
	wire [4-1:0] node16279;
	wire [4-1:0] node16280;
	wire [4-1:0] node16282;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16289;
	wire [4-1:0] node16291;
	wire [4-1:0] node16294;
	wire [4-1:0] node16295;
	wire [4-1:0] node16296;
	wire [4-1:0] node16299;
	wire [4-1:0] node16302;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16307;
	wire [4-1:0] node16308;
	wire [4-1:0] node16309;
	wire [4-1:0] node16312;
	wire [4-1:0] node16315;
	wire [4-1:0] node16316;
	wire [4-1:0] node16319;
	wire [4-1:0] node16322;
	wire [4-1:0] node16323;
	wire [4-1:0] node16324;
	wire [4-1:0] node16325;
	wire [4-1:0] node16328;
	wire [4-1:0] node16331;
	wire [4-1:0] node16333;
	wire [4-1:0] node16334;
	wire [4-1:0] node16335;
	wire [4-1:0] node16339;
	wire [4-1:0] node16341;
	wire [4-1:0] node16344;
	wire [4-1:0] node16345;
	wire [4-1:0] node16346;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16352;
	wire [4-1:0] node16356;
	wire [4-1:0] node16357;
	wire [4-1:0] node16361;
	wire [4-1:0] node16362;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16365;
	wire [4-1:0] node16369;
	wire [4-1:0] node16370;
	wire [4-1:0] node16373;
	wire [4-1:0] node16376;
	wire [4-1:0] node16377;
	wire [4-1:0] node16378;
	wire [4-1:0] node16381;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16388;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16397;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16403;
	wire [4-1:0] node16407;
	wire [4-1:0] node16408;
	wire [4-1:0] node16411;
	wire [4-1:0] node16414;
	wire [4-1:0] node16415;
	wire [4-1:0] node16416;
	wire [4-1:0] node16417;
	wire [4-1:0] node16418;
	wire [4-1:0] node16421;
	wire [4-1:0] node16422;
	wire [4-1:0] node16425;
	wire [4-1:0] node16427;
	wire [4-1:0] node16428;
	wire [4-1:0] node16429;
	wire [4-1:0] node16433;
	wire [4-1:0] node16435;
	wire [4-1:0] node16438;
	wire [4-1:0] node16439;
	wire [4-1:0] node16440;
	wire [4-1:0] node16441;
	wire [4-1:0] node16444;
	wire [4-1:0] node16447;
	wire [4-1:0] node16448;
	wire [4-1:0] node16452;
	wire [4-1:0] node16453;
	wire [4-1:0] node16454;
	wire [4-1:0] node16457;
	wire [4-1:0] node16460;
	wire [4-1:0] node16463;
	wire [4-1:0] node16464;
	wire [4-1:0] node16465;
	wire [4-1:0] node16466;
	wire [4-1:0] node16467;
	wire [4-1:0] node16470;
	wire [4-1:0] node16473;
	wire [4-1:0] node16474;
	wire [4-1:0] node16475;
	wire [4-1:0] node16478;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16484;
	wire [4-1:0] node16487;
	wire [4-1:0] node16490;
	wire [4-1:0] node16491;
	wire [4-1:0] node16492;
	wire [4-1:0] node16494;
	wire [4-1:0] node16499;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16503;
	wire [4-1:0] node16505;
	wire [4-1:0] node16510;
	wire [4-1:0] node16511;
	wire [4-1:0] node16512;
	wire [4-1:0] node16513;
	wire [4-1:0] node16517;
	wire [4-1:0] node16518;
	wire [4-1:0] node16521;
	wire [4-1:0] node16525;
	wire [4-1:0] node16526;
	wire [4-1:0] node16527;
	wire [4-1:0] node16530;
	wire [4-1:0] node16533;
	wire [4-1:0] node16535;
	wire [4-1:0] node16538;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16541;
	wire [4-1:0] node16542;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16548;
	wire [4-1:0] node16549;
	wire [4-1:0] node16553;
	wire [4-1:0] node16554;
	wire [4-1:0] node16555;
	wire [4-1:0] node16559;
	wire [4-1:0] node16561;
	wire [4-1:0] node16562;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16571;
	wire [4-1:0] node16573;
	wire [4-1:0] node16576;
	wire [4-1:0] node16577;
	wire [4-1:0] node16579;
	wire [4-1:0] node16582;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16589;
	wire [4-1:0] node16590;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16596;
	wire [4-1:0] node16599;
	wire [4-1:0] node16600;
	wire [4-1:0] node16602;
	wire [4-1:0] node16605;
	wire [4-1:0] node16606;
	wire [4-1:0] node16609;
	wire [4-1:0] node16612;
	wire [4-1:0] node16613;
	wire [4-1:0] node16614;
	wire [4-1:0] node16615;
	wire [4-1:0] node16617;
	wire [4-1:0] node16620;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16634;
	wire [4-1:0] node16635;
	wire [4-1:0] node16638;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16645;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16651;
	wire [4-1:0] node16654;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16661;
	wire [4-1:0] node16662;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16668;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16674;
	wire [4-1:0] node16678;
	wire [4-1:0] node16679;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16685;
	wire [4-1:0] node16687;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16695;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16700;
	wire [4-1:0] node16703;
	wire [4-1:0] node16706;
	wire [4-1:0] node16707;
	wire [4-1:0] node16708;
	wire [4-1:0] node16712;
	wire [4-1:0] node16715;
	wire [4-1:0] node16716;
	wire [4-1:0] node16717;
	wire [4-1:0] node16719;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16730;
	wire [4-1:0] node16733;
	wire [4-1:0] node16735;
	wire [4-1:0] node16738;
	wire [4-1:0] node16739;
	wire [4-1:0] node16740;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16745;
	wire [4-1:0] node16747;
	wire [4-1:0] node16750;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16755;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16762;
	wire [4-1:0] node16765;
	wire [4-1:0] node16766;
	wire [4-1:0] node16767;
	wire [4-1:0] node16770;
	wire [4-1:0] node16773;
	wire [4-1:0] node16776;
	wire [4-1:0] node16777;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16784;
	wire [4-1:0] node16785;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16792;
	wire [4-1:0] node16795;
	wire [4-1:0] node16796;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16802;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16807;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16817;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16822;
	wire [4-1:0] node16826;
	wire [4-1:0] node16827;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16837;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16845;
	wire [4-1:0] node16846;
	wire [4-1:0] node16847;
	wire [4-1:0] node16848;
	wire [4-1:0] node16849;
	wire [4-1:0] node16851;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16858;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16865;
	wire [4-1:0] node16866;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16878;
	wire [4-1:0] node16879;
	wire [4-1:0] node16880;
	wire [4-1:0] node16881;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16892;
	wire [4-1:0] node16895;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16901;
	wire [4-1:0] node16902;
	wire [4-1:0] node16906;
	wire [4-1:0] node16907;
	wire [4-1:0] node16908;
	wire [4-1:0] node16910;
	wire [4-1:0] node16913;
	wire [4-1:0] node16914;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16923;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16936;
	wire [4-1:0] node16939;
	wire [4-1:0] node16940;
	wire [4-1:0] node16942;
	wire [4-1:0] node16945;
	wire [4-1:0] node16947;
	wire [4-1:0] node16950;
	wire [4-1:0] node16951;
	wire [4-1:0] node16953;
	wire [4-1:0] node16954;
	wire [4-1:0] node16958;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16964;
	wire [4-1:0] node16966;
	wire [4-1:0] node16969;
	wire [4-1:0] node16970;
	wire [4-1:0] node16971;
	wire [4-1:0] node16972;
	wire [4-1:0] node16973;
	wire [4-1:0] node16977;
	wire [4-1:0] node16978;
	wire [4-1:0] node16982;
	wire [4-1:0] node16983;
	wire [4-1:0] node16984;
	wire [4-1:0] node16988;
	wire [4-1:0] node16991;
	wire [4-1:0] node16992;
	wire [4-1:0] node16993;
	wire [4-1:0] node16995;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17003;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17009;
	wire [4-1:0] node17012;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17015;
	wire [4-1:0] node17016;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17020;
	wire [4-1:0] node17021;
	wire [4-1:0] node17025;
	wire [4-1:0] node17027;
	wire [4-1:0] node17029;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17036;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17043;
	wire [4-1:0] node17046;
	wire [4-1:0] node17047;
	wire [4-1:0] node17048;
	wire [4-1:0] node17052;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17057;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17063;
	wire [4-1:0] node17065;
	wire [4-1:0] node17066;
	wire [4-1:0] node17070;
	wire [4-1:0] node17071;
	wire [4-1:0] node17073;
	wire [4-1:0] node17077;
	wire [4-1:0] node17078;
	wire [4-1:0] node17079;
	wire [4-1:0] node17081;
	wire [4-1:0] node17084;
	wire [4-1:0] node17086;
	wire [4-1:0] node17089;
	wire [4-1:0] node17090;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17097;
	wire [4-1:0] node17100;
	wire [4-1:0] node17101;
	wire [4-1:0] node17102;
	wire [4-1:0] node17103;
	wire [4-1:0] node17106;
	wire [4-1:0] node17107;
	wire [4-1:0] node17109;
	wire [4-1:0] node17112;
	wire [4-1:0] node17113;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17119;
	wire [4-1:0] node17121;
	wire [4-1:0] node17124;
	wire [4-1:0] node17125;
	wire [4-1:0] node17126;
	wire [4-1:0] node17130;
	wire [4-1:0] node17132;
	wire [4-1:0] node17135;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17140;
	wire [4-1:0] node17143;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17148;
	wire [4-1:0] node17150;
	wire [4-1:0] node17152;
	wire [4-1:0] node17154;
	wire [4-1:0] node17157;
	wire [4-1:0] node17159;
	wire [4-1:0] node17161;
	wire [4-1:0] node17164;
	wire [4-1:0] node17165;
	wire [4-1:0] node17166;
	wire [4-1:0] node17168;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17176;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17187;
	wire [4-1:0] node17189;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17196;
	wire [4-1:0] node17199;
	wire [4-1:0] node17200;
	wire [4-1:0] node17201;
	wire [4-1:0] node17202;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17208;
	wire [4-1:0] node17210;
	wire [4-1:0] node17213;
	wire [4-1:0] node17214;
	wire [4-1:0] node17216;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17222;
	wire [4-1:0] node17223;
	wire [4-1:0] node17226;
	wire [4-1:0] node17229;
	wire [4-1:0] node17230;
	wire [4-1:0] node17234;
	wire [4-1:0] node17235;
	wire [4-1:0] node17239;
	wire [4-1:0] node17240;
	wire [4-1:0] node17241;
	wire [4-1:0] node17243;
	wire [4-1:0] node17244;
	wire [4-1:0] node17250;
	wire [4-1:0] node17251;
	wire [4-1:0] node17252;
	wire [4-1:0] node17253;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17259;
	wire [4-1:0] node17263;
	wire [4-1:0] node17264;
	wire [4-1:0] node17265;
	wire [4-1:0] node17268;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17276;
	wire [4-1:0] node17278;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17288;
	wire [4-1:0] node17289;
	wire [4-1:0] node17293;
	wire [4-1:0] node17295;
	wire [4-1:0] node17296;
	wire [4-1:0] node17297;
	wire [4-1:0] node17302;
	wire [4-1:0] node17303;
	wire [4-1:0] node17304;
	wire [4-1:0] node17305;
	wire [4-1:0] node17307;
	wire [4-1:0] node17311;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17318;
	wire [4-1:0] node17319;
	wire [4-1:0] node17322;
	wire [4-1:0] node17325;
	wire [4-1:0] node17326;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17332;
	wire [4-1:0] node17335;
	wire [4-1:0] node17337;
	wire [4-1:0] node17340;
	wire [4-1:0] node17341;
	wire [4-1:0] node17342;
	wire [4-1:0] node17344;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17353;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17357;
	wire [4-1:0] node17359;
	wire [4-1:0] node17362;
	wire [4-1:0] node17365;
	wire [4-1:0] node17366;
	wire [4-1:0] node17368;
	wire [4-1:0] node17371;
	wire [4-1:0] node17374;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17378;
	wire [4-1:0] node17381;
	wire [4-1:0] node17382;
	wire [4-1:0] node17386;
	wire [4-1:0] node17389;
	wire [4-1:0] node17390;
	wire [4-1:0] node17391;
	wire [4-1:0] node17392;
	wire [4-1:0] node17393;
	wire [4-1:0] node17394;
	wire [4-1:0] node17398;
	wire [4-1:0] node17399;
	wire [4-1:0] node17402;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17415;
	wire [4-1:0] node17418;
	wire [4-1:0] node17420;
	wire [4-1:0] node17423;
	wire [4-1:0] node17424;
	wire [4-1:0] node17425;
	wire [4-1:0] node17427;
	wire [4-1:0] node17430;
	wire [4-1:0] node17431;
	wire [4-1:0] node17435;
	wire [4-1:0] node17438;
	wire [4-1:0] node17439;
	wire [4-1:0] node17440;
	wire [4-1:0] node17441;
	wire [4-1:0] node17442;
	wire [4-1:0] node17443;
	wire [4-1:0] node17444;
	wire [4-1:0] node17447;
	wire [4-1:0] node17450;
	wire [4-1:0] node17451;
	wire [4-1:0] node17452;
	wire [4-1:0] node17455;
	wire [4-1:0] node17458;
	wire [4-1:0] node17459;
	wire [4-1:0] node17463;
	wire [4-1:0] node17464;
	wire [4-1:0] node17465;
	wire [4-1:0] node17466;
	wire [4-1:0] node17469;
	wire [4-1:0] node17473;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17476;
	wire [4-1:0] node17479;
	wire [4-1:0] node17482;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17489;
	wire [4-1:0] node17490;
	wire [4-1:0] node17493;
	wire [4-1:0] node17496;
	wire [4-1:0] node17497;
	wire [4-1:0] node17498;
	wire [4-1:0] node17499;
	wire [4-1:0] node17501;
	wire [4-1:0] node17503;
	wire [4-1:0] node17506;
	wire [4-1:0] node17507;
	wire [4-1:0] node17508;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17517;
	wire [4-1:0] node17518;
	wire [4-1:0] node17521;
	wire [4-1:0] node17522;
	wire [4-1:0] node17526;
	wire [4-1:0] node17527;
	wire [4-1:0] node17531;
	wire [4-1:0] node17532;
	wire [4-1:0] node17534;
	wire [4-1:0] node17536;
	wire [4-1:0] node17539;
	wire [4-1:0] node17541;
	wire [4-1:0] node17542;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17548;
	wire [4-1:0] node17549;
	wire [4-1:0] node17550;
	wire [4-1:0] node17554;
	wire [4-1:0] node17555;
	wire [4-1:0] node17556;
	wire [4-1:0] node17559;
	wire [4-1:0] node17563;
	wire [4-1:0] node17564;
	wire [4-1:0] node17567;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17574;
	wire [4-1:0] node17575;
	wire [4-1:0] node17576;
	wire [4-1:0] node17577;
	wire [4-1:0] node17580;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17589;
	wire [4-1:0] node17590;
	wire [4-1:0] node17591;
	wire [4-1:0] node17592;
	wire [4-1:0] node17594;
	wire [4-1:0] node17595;
	wire [4-1:0] node17597;
	wire [4-1:0] node17600;
	wire [4-1:0] node17603;
	wire [4-1:0] node17605;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17611;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17617;
	wire [4-1:0] node17618;
	wire [4-1:0] node17619;
	wire [4-1:0] node17623;
	wire [4-1:0] node17626;
	wire [4-1:0] node17628;
	wire [4-1:0] node17629;
	wire [4-1:0] node17633;
	wire [4-1:0] node17634;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17637;
	wire [4-1:0] node17638;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17647;
	wire [4-1:0] node17648;
	wire [4-1:0] node17652;
	wire [4-1:0] node17653;
	wire [4-1:0] node17655;
	wire [4-1:0] node17657;
	wire [4-1:0] node17660;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17671;
	wire [4-1:0] node17672;
	wire [4-1:0] node17673;
	wire [4-1:0] node17675;
	wire [4-1:0] node17676;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17685;
	wire [4-1:0] node17686;
	wire [4-1:0] node17687;
	wire [4-1:0] node17689;
	wire [4-1:0] node17693;
	wire [4-1:0] node17694;
	wire [4-1:0] node17696;
	wire [4-1:0] node17700;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17704;
	wire [4-1:0] node17705;
	wire [4-1:0] node17708;
	wire [4-1:0] node17711;
	wire [4-1:0] node17712;
	wire [4-1:0] node17715;
	wire [4-1:0] node17718;
	wire [4-1:0] node17719;
	wire [4-1:0] node17720;
	wire [4-1:0] node17724;
	wire [4-1:0] node17726;
	wire [4-1:0] node17728;
	wire [4-1:0] node17731;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17739;
	wire [4-1:0] node17743;
	wire [4-1:0] node17744;
	wire [4-1:0] node17745;
	wire [4-1:0] node17748;
	wire [4-1:0] node17751;
	wire [4-1:0] node17754;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17759;
	wire [4-1:0] node17762;
	wire [4-1:0] node17766;
	wire [4-1:0] node17768;
	wire [4-1:0] node17771;
	wire [4-1:0] node17772;
	wire [4-1:0] node17773;
	wire [4-1:0] node17775;
	wire [4-1:0] node17776;
	wire [4-1:0] node17778;
	wire [4-1:0] node17781;
	wire [4-1:0] node17783;
	wire [4-1:0] node17786;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17790;
	wire [4-1:0] node17793;
	wire [4-1:0] node17795;
	wire [4-1:0] node17798;
	wire [4-1:0] node17799;
	wire [4-1:0] node17803;
	wire [4-1:0] node17804;
	wire [4-1:0] node17806;
	wire [4-1:0] node17809;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17812;
	wire [4-1:0] node17815;
	wire [4-1:0] node17819;
	wire [4-1:0] node17820;
	wire [4-1:0] node17823;
	wire [4-1:0] node17826;
	wire [4-1:0] node17827;
	wire [4-1:0] node17828;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17832;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17841;
	wire [4-1:0] node17842;
	wire [4-1:0] node17843;
	wire [4-1:0] node17844;
	wire [4-1:0] node17847;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17857;
	wire [4-1:0] node17860;
	wire [4-1:0] node17861;
	wire [4-1:0] node17866;
	wire [4-1:0] node17867;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17870;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17875;
	wire [4-1:0] node17880;
	wire [4-1:0] node17881;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17887;
	wire [4-1:0] node17888;
	wire [4-1:0] node17893;
	wire [4-1:0] node17894;
	wire [4-1:0] node17895;
	wire [4-1:0] node17898;
	wire [4-1:0] node17902;
	wire [4-1:0] node17903;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17907;
	wire [4-1:0] node17911;
	wire [4-1:0] node17912;
	wire [4-1:0] node17914;
	wire [4-1:0] node17918;
	wire [4-1:0] node17920;
	wire [4-1:0] node17922;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17927;
	wire [4-1:0] node17928;
	wire [4-1:0] node17929;
	wire [4-1:0] node17930;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17934;
	wire [4-1:0] node17936;
	wire [4-1:0] node17939;
	wire [4-1:0] node17941;
	wire [4-1:0] node17944;
	wire [4-1:0] node17946;
	wire [4-1:0] node17947;
	wire [4-1:0] node17949;
	wire [4-1:0] node17952;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17957;
	wire [4-1:0] node17959;
	wire [4-1:0] node17962;
	wire [4-1:0] node17965;
	wire [4-1:0] node17967;
	wire [4-1:0] node17969;
	wire [4-1:0] node17970;
	wire [4-1:0] node17974;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17980;
	wire [4-1:0] node17981;
	wire [4-1:0] node17985;
	wire [4-1:0] node17986;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17994;
	wire [4-1:0] node17995;
	wire [4-1:0] node17996;
	wire [4-1:0] node17998;
	wire [4-1:0] node18002;
	wire [4-1:0] node18003;
	wire [4-1:0] node18006;
	wire [4-1:0] node18009;
	wire [4-1:0] node18010;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18015;
	wire [4-1:0] node18018;
	wire [4-1:0] node18021;
	wire [4-1:0] node18022;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18030;
	wire [4-1:0] node18031;
	wire [4-1:0] node18033;
	wire [4-1:0] node18034;
	wire [4-1:0] node18037;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18042;
	wire [4-1:0] node18045;
	wire [4-1:0] node18049;
	wire [4-1:0] node18050;
	wire [4-1:0] node18051;
	wire [4-1:0] node18052;
	wire [4-1:0] node18055;
	wire [4-1:0] node18058;
	wire [4-1:0] node18059;
	wire [4-1:0] node18060;
	wire [4-1:0] node18063;
	wire [4-1:0] node18067;
	wire [4-1:0] node18068;
	wire [4-1:0] node18071;
	wire [4-1:0] node18074;
	wire [4-1:0] node18075;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18078;
	wire [4-1:0] node18079;
	wire [4-1:0] node18080;
	wire [4-1:0] node18084;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18091;
	wire [4-1:0] node18093;
	wire [4-1:0] node18094;
	wire [4-1:0] node18097;
	wire [4-1:0] node18100;
	wire [4-1:0] node18101;
	wire [4-1:0] node18102;
	wire [4-1:0] node18104;
	wire [4-1:0] node18105;
	wire [4-1:0] node18108;
	wire [4-1:0] node18111;
	wire [4-1:0] node18113;
	wire [4-1:0] node18114;
	wire [4-1:0] node18117;
	wire [4-1:0] node18120;
	wire [4-1:0] node18122;
	wire [4-1:0] node18124;
	wire [4-1:0] node18127;
	wire [4-1:0] node18128;
	wire [4-1:0] node18129;
	wire [4-1:0] node18130;
	wire [4-1:0] node18131;
	wire [4-1:0] node18134;
	wire [4-1:0] node18138;
	wire [4-1:0] node18139;
	wire [4-1:0] node18140;
	wire [4-1:0] node18141;
	wire [4-1:0] node18144;
	wire [4-1:0] node18148;
	wire [4-1:0] node18149;
	wire [4-1:0] node18151;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18158;
	wire [4-1:0] node18161;
	wire [4-1:0] node18162;
	wire [4-1:0] node18163;
	wire [4-1:0] node18164;
	wire [4-1:0] node18169;
	wire [4-1:0] node18170;
	wire [4-1:0] node18171;
	wire [4-1:0] node18173;
	wire [4-1:0] node18177;
	wire [4-1:0] node18180;
	wire [4-1:0] node18181;
	wire [4-1:0] node18182;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18187;
	wire [4-1:0] node18188;
	wire [4-1:0] node18190;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18200;
	wire [4-1:0] node18201;
	wire [4-1:0] node18205;
	wire [4-1:0] node18206;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18212;
	wire [4-1:0] node18214;
	wire [4-1:0] node18215;
	wire [4-1:0] node18216;
	wire [4-1:0] node18221;
	wire [4-1:0] node18223;
	wire [4-1:0] node18225;
	wire [4-1:0] node18228;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18234;
	wire [4-1:0] node18236;
	wire [4-1:0] node18239;
	wire [4-1:0] node18240;
	wire [4-1:0] node18241;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18244;
	wire [4-1:0] node18245;
	wire [4-1:0] node18248;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18257;
	wire [4-1:0] node18258;
	wire [4-1:0] node18260;
	wire [4-1:0] node18261;
	wire [4-1:0] node18264;
	wire [4-1:0] node18267;
	wire [4-1:0] node18268;
	wire [4-1:0] node18269;
	wire [4-1:0] node18274;
	wire [4-1:0] node18275;
	wire [4-1:0] node18276;
	wire [4-1:0] node18279;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18285;
	wire [4-1:0] node18288;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18295;
	wire [4-1:0] node18300;
	wire [4-1:0] node18302;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18307;
	wire [4-1:0] node18310;
	wire [4-1:0] node18313;
	wire [4-1:0] node18314;
	wire [4-1:0] node18315;
	wire [4-1:0] node18319;
	wire [4-1:0] node18320;
	wire [4-1:0] node18323;
	wire [4-1:0] node18326;
	wire [4-1:0] node18327;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18337;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18345;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18355;
	wire [4-1:0] node18356;
	wire [4-1:0] node18359;
	wire [4-1:0] node18362;
	wire [4-1:0] node18363;
	wire [4-1:0] node18364;
	wire [4-1:0] node18365;
	wire [4-1:0] node18368;
	wire [4-1:0] node18371;
	wire [4-1:0] node18373;
	wire [4-1:0] node18374;
	wire [4-1:0] node18375;
	wire [4-1:0] node18378;
	wire [4-1:0] node18382;
	wire [4-1:0] node18383;
	wire [4-1:0] node18384;
	wire [4-1:0] node18386;
	wire [4-1:0] node18387;
	wire [4-1:0] node18391;
	wire [4-1:0] node18392;
	wire [4-1:0] node18395;
	wire [4-1:0] node18398;
	wire [4-1:0] node18399;
	wire [4-1:0] node18400;
	wire [4-1:0] node18403;
	wire [4-1:0] node18406;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18411;
	wire [4-1:0] node18412;
	wire [4-1:0] node18413;
	wire [4-1:0] node18414;
	wire [4-1:0] node18415;
	wire [4-1:0] node18418;
	wire [4-1:0] node18421;
	wire [4-1:0] node18422;
	wire [4-1:0] node18425;
	wire [4-1:0] node18428;
	wire [4-1:0] node18429;
	wire [4-1:0] node18430;
	wire [4-1:0] node18433;
	wire [4-1:0] node18436;
	wire [4-1:0] node18439;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18444;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18450;
	wire [4-1:0] node18451;
	wire [4-1:0] node18455;
	wire [4-1:0] node18456;
	wire [4-1:0] node18459;
	wire [4-1:0] node18462;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18465;
	wire [4-1:0] node18466;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18473;
	wire [4-1:0] node18476;
	wire [4-1:0] node18478;
	wire [4-1:0] node18481;
	wire [4-1:0] node18483;
	wire [4-1:0] node18486;
	wire [4-1:0] node18487;
	wire [4-1:0] node18489;
	wire [4-1:0] node18492;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18498;
	wire [4-1:0] node18501;
	wire [4-1:0] node18502;
	wire [4-1:0] node18503;
	wire [4-1:0] node18504;
	wire [4-1:0] node18505;
	wire [4-1:0] node18509;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18514;
	wire [4-1:0] node18518;
	wire [4-1:0] node18519;
	wire [4-1:0] node18521;
	wire [4-1:0] node18524;
	wire [4-1:0] node18525;
	wire [4-1:0] node18528;
	wire [4-1:0] node18531;
	wire [4-1:0] node18532;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18535;
	wire [4-1:0] node18537;
	wire [4-1:0] node18540;
	wire [4-1:0] node18542;
	wire [4-1:0] node18546;
	wire [4-1:0] node18547;
	wire [4-1:0] node18548;
	wire [4-1:0] node18551;
	wire [4-1:0] node18553;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18560;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18567;
	wire [4-1:0] node18568;
	wire [4-1:0] node18572;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18575;
	wire [4-1:0] node18576;
	wire [4-1:0] node18577;
	wire [4-1:0] node18578;
	wire [4-1:0] node18579;
	wire [4-1:0] node18583;
	wire [4-1:0] node18584;
	wire [4-1:0] node18585;
	wire [4-1:0] node18589;
	wire [4-1:0] node18590;
	wire [4-1:0] node18594;
	wire [4-1:0] node18595;
	wire [4-1:0] node18598;
	wire [4-1:0] node18599;
	wire [4-1:0] node18601;
	wire [4-1:0] node18604;
	wire [4-1:0] node18607;
	wire [4-1:0] node18608;
	wire [4-1:0] node18609;
	wire [4-1:0] node18611;
	wire [4-1:0] node18613;
	wire [4-1:0] node18614;
	wire [4-1:0] node18618;
	wire [4-1:0] node18619;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18625;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18631;
	wire [4-1:0] node18636;
	wire [4-1:0] node18637;
	wire [4-1:0] node18638;
	wire [4-1:0] node18639;
	wire [4-1:0] node18640;
	wire [4-1:0] node18642;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18650;
	wire [4-1:0] node18654;
	wire [4-1:0] node18657;
	wire [4-1:0] node18659;
	wire [4-1:0] node18662;
	wire [4-1:0] node18663;
	wire [4-1:0] node18664;
	wire [4-1:0] node18665;
	wire [4-1:0] node18666;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18675;
	wire [4-1:0] node18677;
	wire [4-1:0] node18680;
	wire [4-1:0] node18681;
	wire [4-1:0] node18682;
	wire [4-1:0] node18683;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18692;
	wire [4-1:0] node18693;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18703;
	wire [4-1:0] node18704;
	wire [4-1:0] node18705;
	wire [4-1:0] node18706;
	wire [4-1:0] node18710;
	wire [4-1:0] node18711;
	wire [4-1:0] node18712;
	wire [4-1:0] node18717;
	wire [4-1:0] node18718;
	wire [4-1:0] node18719;
	wire [4-1:0] node18722;
	wire [4-1:0] node18723;
	wire [4-1:0] node18725;
	wire [4-1:0] node18728;
	wire [4-1:0] node18729;
	wire [4-1:0] node18733;
	wire [4-1:0] node18734;
	wire [4-1:0] node18735;
	wire [4-1:0] node18736;
	wire [4-1:0] node18741;
	wire [4-1:0] node18743;
	wire [4-1:0] node18746;
	wire [4-1:0] node18747;
	wire [4-1:0] node18748;
	wire [4-1:0] node18749;
	wire [4-1:0] node18752;
	wire [4-1:0] node18753;
	wire [4-1:0] node18757;
	wire [4-1:0] node18758;
	wire [4-1:0] node18759;
	wire [4-1:0] node18763;
	wire [4-1:0] node18764;
	wire [4-1:0] node18768;
	wire [4-1:0] node18769;
	wire [4-1:0] node18770;
	wire [4-1:0] node18771;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18781;
	wire [4-1:0] node18782;
	wire [4-1:0] node18783;
	wire [4-1:0] node18784;
	wire [4-1:0] node18785;
	wire [4-1:0] node18787;
	wire [4-1:0] node18790;
	wire [4-1:0] node18792;
	wire [4-1:0] node18795;
	wire [4-1:0] node18796;
	wire [4-1:0] node18797;
	wire [4-1:0] node18799;
	wire [4-1:0] node18802;
	wire [4-1:0] node18805;
	wire [4-1:0] node18806;
	wire [4-1:0] node18809;
	wire [4-1:0] node18811;
	wire [4-1:0] node18814;
	wire [4-1:0] node18815;
	wire [4-1:0] node18817;
	wire [4-1:0] node18820;
	wire [4-1:0] node18822;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18827;
	wire [4-1:0] node18829;
	wire [4-1:0] node18830;
	wire [4-1:0] node18833;
	wire [4-1:0] node18836;
	wire [4-1:0] node18837;
	wire [4-1:0] node18838;
	wire [4-1:0] node18841;
	wire [4-1:0] node18844;
	wire [4-1:0] node18846;
	wire [4-1:0] node18848;
	wire [4-1:0] node18851;
	wire [4-1:0] node18852;
	wire [4-1:0] node18853;
	wire [4-1:0] node18857;
	wire [4-1:0] node18858;
	wire [4-1:0] node18861;
	wire [4-1:0] node18864;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18873;
	wire [4-1:0] node18877;
	wire [4-1:0] node18878;
	wire [4-1:0] node18879;
	wire [4-1:0] node18880;
	wire [4-1:0] node18882;
	wire [4-1:0] node18885;
	wire [4-1:0] node18887;
	wire [4-1:0] node18891;
	wire [4-1:0] node18892;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18899;
	wire [4-1:0] node18900;
	wire [4-1:0] node18904;
	wire [4-1:0] node18905;
	wire [4-1:0] node18906;
	wire [4-1:0] node18907;
	wire [4-1:0] node18908;
	wire [4-1:0] node18910;
	wire [4-1:0] node18913;
	wire [4-1:0] node18917;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18923;
	wire [4-1:0] node18925;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18931;
	wire [4-1:0] node18934;
	wire [4-1:0] node18935;
	wire [4-1:0] node18937;
	wire [4-1:0] node18940;
	wire [4-1:0] node18942;
	wire [4-1:0] node18945;
	wire [4-1:0] node18946;
	wire [4-1:0] node18947;
	wire [4-1:0] node18948;
	wire [4-1:0] node18949;
	wire [4-1:0] node18950;
	wire [4-1:0] node18952;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18959;
	wire [4-1:0] node18962;
	wire [4-1:0] node18963;
	wire [4-1:0] node18967;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18970;
	wire [4-1:0] node18973;
	wire [4-1:0] node18977;
	wire [4-1:0] node18978;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18986;
	wire [4-1:0] node18988;
	wire [4-1:0] node18991;
	wire [4-1:0] node18992;
	wire [4-1:0] node18993;
	wire [4-1:0] node18994;
	wire [4-1:0] node18998;
	wire [4-1:0] node18999;
	wire [4-1:0] node19003;
	wire [4-1:0] node19004;
	wire [4-1:0] node19005;
	wire [4-1:0] node19007;
	wire [4-1:0] node19008;
	wire [4-1:0] node19013;
	wire [4-1:0] node19014;
	wire [4-1:0] node19015;
	wire [4-1:0] node19020;
	wire [4-1:0] node19021;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19026;
	wire [4-1:0] node19029;
	wire [4-1:0] node19030;
	wire [4-1:0] node19031;
	wire [4-1:0] node19032;
	wire [4-1:0] node19036;
	wire [4-1:0] node19037;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19046;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19050;
	wire [4-1:0] node19054;
	wire [4-1:0] node19055;
	wire [4-1:0] node19057;
	wire [4-1:0] node19060;
	wire [4-1:0] node19061;
	wire [4-1:0] node19062;
	wire [4-1:0] node19065;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19076;
	wire [4-1:0] node19080;
	wire [4-1:0] node19081;
	wire [4-1:0] node19082;
	wire [4-1:0] node19086;
	wire [4-1:0] node19087;
	wire [4-1:0] node19091;
	wire [4-1:0] node19093;
	wire [4-1:0] node19094;
	wire [4-1:0] node19095;
	wire [4-1:0] node19096;
	wire [4-1:0] node19099;
	wire [4-1:0] node19103;
	wire [4-1:0] node19104;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19114;
	wire [4-1:0] node19117;
	wire [4-1:0] node19119;
	wire [4-1:0] node19122;
	wire [4-1:0] node19124;
	wire [4-1:0] node19125;
	wire [4-1:0] node19127;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19135;
	wire [4-1:0] node19136;
	wire [4-1:0] node19137;
	wire [4-1:0] node19139;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19147;
	wire [4-1:0] node19150;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19153;
	wire [4-1:0] node19154;
	wire [4-1:0] node19159;
	wire [4-1:0] node19160;
	wire [4-1:0] node19161;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19171;
	wire [4-1:0] node19174;
	wire [4-1:0] node19175;
	wire [4-1:0] node19176;
	wire [4-1:0] node19181;
	wire [4-1:0] node19182;
	wire [4-1:0] node19183;
	wire [4-1:0] node19184;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19187;
	wire [4-1:0] node19188;
	wire [4-1:0] node19189;
	wire [4-1:0] node19190;
	wire [4-1:0] node19193;
	wire [4-1:0] node19196;
	wire [4-1:0] node19197;
	wire [4-1:0] node19201;
	wire [4-1:0] node19202;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19208;
	wire [4-1:0] node19209;
	wire [4-1:0] node19212;
	wire [4-1:0] node19215;
	wire [4-1:0] node19217;
	wire [4-1:0] node19220;
	wire [4-1:0] node19221;
	wire [4-1:0] node19223;
	wire [4-1:0] node19225;
	wire [4-1:0] node19229;
	wire [4-1:0] node19230;
	wire [4-1:0] node19231;
	wire [4-1:0] node19232;
	wire [4-1:0] node19235;
	wire [4-1:0] node19239;
	wire [4-1:0] node19240;
	wire [4-1:0] node19241;
	wire [4-1:0] node19243;
	wire [4-1:0] node19245;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19250;
	wire [4-1:0] node19255;
	wire [4-1:0] node19256;
	wire [4-1:0] node19257;
	wire [4-1:0] node19261;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19271;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19279;
	wire [4-1:0] node19282;
	wire [4-1:0] node19284;
	wire [4-1:0] node19287;
	wire [4-1:0] node19288;
	wire [4-1:0] node19290;
	wire [4-1:0] node19293;
	wire [4-1:0] node19295;
	wire [4-1:0] node19298;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19303;
	wire [4-1:0] node19306;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19309;
	wire [4-1:0] node19313;
	wire [4-1:0] node19314;
	wire [4-1:0] node19317;
	wire [4-1:0] node19320;
	wire [4-1:0] node19321;
	wire [4-1:0] node19324;
	wire [4-1:0] node19327;
	wire [4-1:0] node19328;
	wire [4-1:0] node19331;
	wire [4-1:0] node19334;
	wire [4-1:0] node19335;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19338;
	wire [4-1:0] node19339;
	wire [4-1:0] node19341;
	wire [4-1:0] node19344;
	wire [4-1:0] node19346;
	wire [4-1:0] node19349;
	wire [4-1:0] node19350;
	wire [4-1:0] node19352;
	wire [4-1:0] node19355;
	wire [4-1:0] node19356;
	wire [4-1:0] node19360;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19365;
	wire [4-1:0] node19367;
	wire [4-1:0] node19370;
	wire [4-1:0] node19371;
	wire [4-1:0] node19375;
	wire [4-1:0] node19376;
	wire [4-1:0] node19377;
	wire [4-1:0] node19381;
	wire [4-1:0] node19383;
	wire [4-1:0] node19386;
	wire [4-1:0] node19387;
	wire [4-1:0] node19389;
	wire [4-1:0] node19390;
	wire [4-1:0] node19394;
	wire [4-1:0] node19395;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19401;
	wire [4-1:0] node19402;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19410;
	wire [4-1:0] node19411;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19418;
	wire [4-1:0] node19419;
	wire [4-1:0] node19423;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19431;
	wire [4-1:0] node19433;
	wire [4-1:0] node19436;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19447;
	wire [4-1:0] node19448;
	wire [4-1:0] node19450;
	wire [4-1:0] node19453;
	wire [4-1:0] node19455;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19461;
	wire [4-1:0] node19462;
	wire [4-1:0] node19464;
	wire [4-1:0] node19465;
	wire [4-1:0] node19468;
	wire [4-1:0] node19472;
	wire [4-1:0] node19473;
	wire [4-1:0] node19475;
	wire [4-1:0] node19478;
	wire [4-1:0] node19479;
	wire [4-1:0] node19480;
	wire [4-1:0] node19484;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19489;
	wire [4-1:0] node19491;
	wire [4-1:0] node19494;
	wire [4-1:0] node19495;
	wire [4-1:0] node19497;
	wire [4-1:0] node19500;
	wire [4-1:0] node19502;
	wire [4-1:0] node19505;
	wire [4-1:0] node19506;
	wire [4-1:0] node19508;
	wire [4-1:0] node19511;
	wire [4-1:0] node19512;
	wire [4-1:0] node19514;
	wire [4-1:0] node19517;
	wire [4-1:0] node19520;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19524;
	wire [4-1:0] node19525;
	wire [4-1:0] node19526;
	wire [4-1:0] node19529;
	wire [4-1:0] node19534;
	wire [4-1:0] node19536;
	wire [4-1:0] node19537;
	wire [4-1:0] node19540;
	wire [4-1:0] node19543;
	wire [4-1:0] node19544;
	wire [4-1:0] node19545;
	wire [4-1:0] node19546;
	wire [4-1:0] node19549;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19556;
	wire [4-1:0] node19559;
	wire [4-1:0] node19561;
	wire [4-1:0] node19562;
	wire [4-1:0] node19563;
	wire [4-1:0] node19567;
	wire [4-1:0] node19569;
	wire [4-1:0] node19572;
	wire [4-1:0] node19573;
	wire [4-1:0] node19574;
	wire [4-1:0] node19575;
	wire [4-1:0] node19578;
	wire [4-1:0] node19581;
	wire [4-1:0] node19582;
	wire [4-1:0] node19584;
	wire [4-1:0] node19586;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19594;
	wire [4-1:0] node19595;
	wire [4-1:0] node19597;
	wire [4-1:0] node19598;
	wire [4-1:0] node19601;
	wire [4-1:0] node19604;
	wire [4-1:0] node19605;
	wire [4-1:0] node19608;
	wire [4-1:0] node19611;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19621;
	wire [4-1:0] node19624;
	wire [4-1:0] node19626;
	wire [4-1:0] node19629;
	wire [4-1:0] node19630;
	wire [4-1:0] node19633;
	wire [4-1:0] node19636;
	wire [4-1:0] node19637;
	wire [4-1:0] node19640;
	wire [4-1:0] node19643;
	wire [4-1:0] node19644;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19654;
	wire [4-1:0] node19655;
	wire [4-1:0] node19659;
	wire [4-1:0] node19660;
	wire [4-1:0] node19662;
	wire [4-1:0] node19664;
	wire [4-1:0] node19667;
	wire [4-1:0] node19668;
	wire [4-1:0] node19671;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19681;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19688;
	wire [4-1:0] node19691;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19695;
	wire [4-1:0] node19696;
	wire [4-1:0] node19700;
	wire [4-1:0] node19702;
	wire [4-1:0] node19705;
	wire [4-1:0] node19706;
	wire [4-1:0] node19709;
	wire [4-1:0] node19712;
	wire [4-1:0] node19714;
	wire [4-1:0] node19717;
	wire [4-1:0] node19719;
	wire [4-1:0] node19720;
	wire [4-1:0] node19721;
	wire [4-1:0] node19724;
	wire [4-1:0] node19727;
	wire [4-1:0] node19728;
	wire [4-1:0] node19731;
	wire [4-1:0] node19734;
	wire [4-1:0] node19735;
	wire [4-1:0] node19736;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19739;
	wire [4-1:0] node19740;
	wire [4-1:0] node19743;
	wire [4-1:0] node19747;
	wire [4-1:0] node19748;
	wire [4-1:0] node19750;
	wire [4-1:0] node19753;
	wire [4-1:0] node19754;
	wire [4-1:0] node19758;
	wire [4-1:0] node19759;
	wire [4-1:0] node19761;
	wire [4-1:0] node19764;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19771;
	wire [4-1:0] node19774;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19778;
	wire [4-1:0] node19781;
	wire [4-1:0] node19782;
	wire [4-1:0] node19785;
	wire [4-1:0] node19788;
	wire [4-1:0] node19789;
	wire [4-1:0] node19790;
	wire [4-1:0] node19791;
	wire [4-1:0] node19795;
	wire [4-1:0] node19796;
	wire [4-1:0] node19799;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19806;
	wire [4-1:0] node19809;
	wire [4-1:0] node19810;
	wire [4-1:0] node19811;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19814;
	wire [4-1:0] node19818;
	wire [4-1:0] node19819;
	wire [4-1:0] node19823;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19829;
	wire [4-1:0] node19830;
	wire [4-1:0] node19835;
	wire [4-1:0] node19836;
	wire [4-1:0] node19837;
	wire [4-1:0] node19838;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19848;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19851;
	wire [4-1:0] node19852;
	wire [4-1:0] node19853;
	wire [4-1:0] node19854;
	wire [4-1:0] node19855;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19859;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19865;
	wire [4-1:0] node19867;
	wire [4-1:0] node19870;
	wire [4-1:0] node19871;
	wire [4-1:0] node19872;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19881;
	wire [4-1:0] node19884;
	wire [4-1:0] node19885;
	wire [4-1:0] node19888;
	wire [4-1:0] node19891;
	wire [4-1:0] node19892;
	wire [4-1:0] node19894;
	wire [4-1:0] node19895;
	wire [4-1:0] node19897;
	wire [4-1:0] node19900;
	wire [4-1:0] node19903;
	wire [4-1:0] node19904;
	wire [4-1:0] node19905;
	wire [4-1:0] node19908;
	wire [4-1:0] node19911;
	wire [4-1:0] node19912;
	wire [4-1:0] node19914;
	wire [4-1:0] node19918;
	wire [4-1:0] node19919;
	wire [4-1:0] node19920;
	wire [4-1:0] node19922;
	wire [4-1:0] node19924;
	wire [4-1:0] node19927;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19934;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19941;
	wire [4-1:0] node19942;
	wire [4-1:0] node19943;
	wire [4-1:0] node19948;
	wire [4-1:0] node19949;
	wire [4-1:0] node19951;
	wire [4-1:0] node19954;
	wire [4-1:0] node19957;
	wire [4-1:0] node19958;
	wire [4-1:0] node19959;
	wire [4-1:0] node19960;
	wire [4-1:0] node19962;
	wire [4-1:0] node19964;
	wire [4-1:0] node19966;
	wire [4-1:0] node19969;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19976;
	wire [4-1:0] node19977;
	wire [4-1:0] node19979;
	wire [4-1:0] node19981;
	wire [4-1:0] node19983;
	wire [4-1:0] node19986;
	wire [4-1:0] node19987;
	wire [4-1:0] node19988;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19999;
	wire [4-1:0] node20003;
	wire [4-1:0] node20004;
	wire [4-1:0] node20005;
	wire [4-1:0] node20007;
	wire [4-1:0] node20008;
	wire [4-1:0] node20009;
	wire [4-1:0] node20012;
	wire [4-1:0] node20016;
	wire [4-1:0] node20018;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20024;
	wire [4-1:0] node20027;
	wire [4-1:0] node20028;
	wire [4-1:0] node20030;
	wire [4-1:0] node20031;
	wire [4-1:0] node20033;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20041;
	wire [4-1:0] node20042;
	wire [4-1:0] node20043;
	wire [4-1:0] node20047;
	wire [4-1:0] node20049;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20056;
	wire [4-1:0] node20057;
	wire [4-1:0] node20060;
	wire [4-1:0] node20061;
	wire [4-1:0] node20062;
	wire [4-1:0] node20067;
	wire [4-1:0] node20068;
	wire [4-1:0] node20071;
	wire [4-1:0] node20073;
	wire [4-1:0] node20076;
	wire [4-1:0] node20077;
	wire [4-1:0] node20079;
	wire [4-1:0] node20080;
	wire [4-1:0] node20083;
	wire [4-1:0] node20086;
	wire [4-1:0] node20087;
	wire [4-1:0] node20088;
	wire [4-1:0] node20091;
	wire [4-1:0] node20094;
	wire [4-1:0] node20095;
	wire [4-1:0] node20096;
	wire [4-1:0] node20101;
	wire [4-1:0] node20102;
	wire [4-1:0] node20103;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20115;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20122;
	wire [4-1:0] node20126;
	wire [4-1:0] node20129;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20133;
	wire [4-1:0] node20136;
	wire [4-1:0] node20138;
	wire [4-1:0] node20141;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20146;
	wire [4-1:0] node20149;
	wire [4-1:0] node20150;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20158;
	wire [4-1:0] node20160;
	wire [4-1:0] node20164;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20170;
	wire [4-1:0] node20171;
	wire [4-1:0] node20175;
	wire [4-1:0] node20176;
	wire [4-1:0] node20177;
	wire [4-1:0] node20178;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20187;
	wire [4-1:0] node20189;
	wire [4-1:0] node20190;
	wire [4-1:0] node20192;
	wire [4-1:0] node20196;
	wire [4-1:0] node20197;
	wire [4-1:0] node20198;
	wire [4-1:0] node20200;
	wire [4-1:0] node20202;
	wire [4-1:0] node20205;
	wire [4-1:0] node20206;
	wire [4-1:0] node20207;
	wire [4-1:0] node20212;
	wire [4-1:0] node20213;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20219;
	wire [4-1:0] node20220;
	wire [4-1:0] node20224;
	wire [4-1:0] node20226;
	wire [4-1:0] node20228;
	wire [4-1:0] node20231;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20234;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20238;
	wire [4-1:0] node20240;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20245;
	wire [4-1:0] node20248;
	wire [4-1:0] node20251;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20257;
	wire [4-1:0] node20258;
	wire [4-1:0] node20260;
	wire [4-1:0] node20263;
	wire [4-1:0] node20264;
	wire [4-1:0] node20267;
	wire [4-1:0] node20269;
	wire [4-1:0] node20272;
	wire [4-1:0] node20273;
	wire [4-1:0] node20275;
	wire [4-1:0] node20278;
	wire [4-1:0] node20279;
	wire [4-1:0] node20283;
	wire [4-1:0] node20284;
	wire [4-1:0] node20285;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20289;
	wire [4-1:0] node20294;
	wire [4-1:0] node20295;
	wire [4-1:0] node20296;
	wire [4-1:0] node20299;
	wire [4-1:0] node20302;
	wire [4-1:0] node20303;
	wire [4-1:0] node20307;
	wire [4-1:0] node20308;
	wire [4-1:0] node20309;
	wire [4-1:0] node20311;
	wire [4-1:0] node20312;
	wire [4-1:0] node20315;
	wire [4-1:0] node20318;
	wire [4-1:0] node20320;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20325;
	wire [4-1:0] node20328;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20336;
	wire [4-1:0] node20337;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20340;
	wire [4-1:0] node20342;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20347;
	wire [4-1:0] node20350;
	wire [4-1:0] node20354;
	wire [4-1:0] node20355;
	wire [4-1:0] node20356;
	wire [4-1:0] node20359;
	wire [4-1:0] node20363;
	wire [4-1:0] node20364;
	wire [4-1:0] node20366;
	wire [4-1:0] node20367;
	wire [4-1:0] node20370;
	wire [4-1:0] node20373;
	wire [4-1:0] node20375;
	wire [4-1:0] node20377;
	wire [4-1:0] node20378;
	wire [4-1:0] node20381;
	wire [4-1:0] node20384;
	wire [4-1:0] node20385;
	wire [4-1:0] node20386;
	wire [4-1:0] node20387;
	wire [4-1:0] node20389;
	wire [4-1:0] node20390;
	wire [4-1:0] node20393;
	wire [4-1:0] node20396;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20402;
	wire [4-1:0] node20405;
	wire [4-1:0] node20407;
	wire [4-1:0] node20408;
	wire [4-1:0] node20412;
	wire [4-1:0] node20413;
	wire [4-1:0] node20414;
	wire [4-1:0] node20417;
	wire [4-1:0] node20420;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20425;
	wire [4-1:0] node20428;
	wire [4-1:0] node20431;
	wire [4-1:0] node20432;
	wire [4-1:0] node20433;
	wire [4-1:0] node20434;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20439;
	wire [4-1:0] node20443;
	wire [4-1:0] node20444;
	wire [4-1:0] node20447;
	wire [4-1:0] node20450;
	wire [4-1:0] node20451;
	wire [4-1:0] node20452;
	wire [4-1:0] node20454;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20461;
	wire [4-1:0] node20462;
	wire [4-1:0] node20465;
	wire [4-1:0] node20469;
	wire [4-1:0] node20470;
	wire [4-1:0] node20471;
	wire [4-1:0] node20475;
	wire [4-1:0] node20476;
	wire [4-1:0] node20480;
	wire [4-1:0] node20481;
	wire [4-1:0] node20482;
	wire [4-1:0] node20483;
	wire [4-1:0] node20486;
	wire [4-1:0] node20489;
	wire [4-1:0] node20491;
	wire [4-1:0] node20493;
	wire [4-1:0] node20496;
	wire [4-1:0] node20497;
	wire [4-1:0] node20499;
	wire [4-1:0] node20502;
	wire [4-1:0] node20503;
	wire [4-1:0] node20505;
	wire [4-1:0] node20506;
	wire [4-1:0] node20511;
	wire [4-1:0] node20512;
	wire [4-1:0] node20513;
	wire [4-1:0] node20514;
	wire [4-1:0] node20516;
	wire [4-1:0] node20519;
	wire [4-1:0] node20520;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20530;
	wire [4-1:0] node20531;
	wire [4-1:0] node20535;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20542;
	wire [4-1:0] node20543;
	wire [4-1:0] node20544;
	wire [4-1:0] node20545;
	wire [4-1:0] node20548;
	wire [4-1:0] node20552;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20562;
	wire [4-1:0] node20563;
	wire [4-1:0] node20566;
	wire [4-1:0] node20569;
	wire [4-1:0] node20570;
	wire [4-1:0] node20571;
	wire [4-1:0] node20576;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20581;
	wire [4-1:0] node20582;
	wire [4-1:0] node20583;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20589;
	wire [4-1:0] node20590;
	wire [4-1:0] node20596;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20600;
	wire [4-1:0] node20603;
	wire [4-1:0] node20604;
	wire [4-1:0] node20605;
	wire [4-1:0] node20608;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20616;
	wire [4-1:0] node20617;
	wire [4-1:0] node20620;
	wire [4-1:0] node20621;
	wire [4-1:0] node20624;
	wire [4-1:0] node20627;
	wire [4-1:0] node20628;
	wire [4-1:0] node20629;
	wire [4-1:0] node20630;
	wire [4-1:0] node20631;
	wire [4-1:0] node20635;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20642;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20648;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20654;
	wire [4-1:0] node20657;
	wire [4-1:0] node20658;
	wire [4-1:0] node20660;
	wire [4-1:0] node20661;
	wire [4-1:0] node20664;
	wire [4-1:0] node20667;
	wire [4-1:0] node20669;
	wire [4-1:0] node20670;
	wire [4-1:0] node20672;
	wire [4-1:0] node20675;
	wire [4-1:0] node20676;
	wire [4-1:0] node20680;
	wire [4-1:0] node20681;
	wire [4-1:0] node20682;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20687;
	wire [4-1:0] node20689;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20694;
	wire [4-1:0] node20698;
	wire [4-1:0] node20700;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20705;
	wire [4-1:0] node20707;
	wire [4-1:0] node20711;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20716;
	wire [4-1:0] node20720;
	wire [4-1:0] node20721;
	wire [4-1:0] node20722;
	wire [4-1:0] node20723;
	wire [4-1:0] node20724;
	wire [4-1:0] node20727;
	wire [4-1:0] node20730;
	wire [4-1:0] node20731;
	wire [4-1:0] node20735;
	wire [4-1:0] node20736;
	wire [4-1:0] node20737;
	wire [4-1:0] node20739;
	wire [4-1:0] node20742;
	wire [4-1:0] node20744;
	wire [4-1:0] node20748;
	wire [4-1:0] node20749;
	wire [4-1:0] node20750;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20758;
	wire [4-1:0] node20759;
	wire [4-1:0] node20760;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20771;
	wire [4-1:0] node20772;
	wire [4-1:0] node20773;
	wire [4-1:0] node20774;
	wire [4-1:0] node20775;
	wire [4-1:0] node20776;
	wire [4-1:0] node20777;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20785;
	wire [4-1:0] node20788;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20791;
	wire [4-1:0] node20794;
	wire [4-1:0] node20798;
	wire [4-1:0] node20801;
	wire [4-1:0] node20802;
	wire [4-1:0] node20804;
	wire [4-1:0] node20806;
	wire [4-1:0] node20809;
	wire [4-1:0] node20810;
	wire [4-1:0] node20812;
	wire [4-1:0] node20815;
	wire [4-1:0] node20816;
	wire [4-1:0] node20817;
	wire [4-1:0] node20820;
	wire [4-1:0] node20824;
	wire [4-1:0] node20825;
	wire [4-1:0] node20826;
	wire [4-1:0] node20827;
	wire [4-1:0] node20828;
	wire [4-1:0] node20833;
	wire [4-1:0] node20834;
	wire [4-1:0] node20837;
	wire [4-1:0] node20839;
	wire [4-1:0] node20840;
	wire [4-1:0] node20844;
	wire [4-1:0] node20845;
	wire [4-1:0] node20846;
	wire [4-1:0] node20847;
	wire [4-1:0] node20848;
	wire [4-1:0] node20851;
	wire [4-1:0] node20855;
	wire [4-1:0] node20856;
	wire [4-1:0] node20859;
	wire [4-1:0] node20862;
	wire [4-1:0] node20863;
	wire [4-1:0] node20864;
	wire [4-1:0] node20867;
	wire [4-1:0] node20869;
	wire [4-1:0] node20872;
	wire [4-1:0] node20873;
	wire [4-1:0] node20876;
	wire [4-1:0] node20879;
	wire [4-1:0] node20880;
	wire [4-1:0] node20881;
	wire [4-1:0] node20882;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20889;
	wire [4-1:0] node20890;
	wire [4-1:0] node20891;
	wire [4-1:0] node20892;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20902;
	wire [4-1:0] node20903;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20907;
	wire [4-1:0] node20911;
	wire [4-1:0] node20913;
	wire [4-1:0] node20916;
	wire [4-1:0] node20918;
	wire [4-1:0] node20919;
	wire [4-1:0] node20922;
	wire [4-1:0] node20925;
	wire [4-1:0] node20926;
	wire [4-1:0] node20927;
	wire [4-1:0] node20928;
	wire [4-1:0] node20929;
	wire [4-1:0] node20934;
	wire [4-1:0] node20935;
	wire [4-1:0] node20937;
	wire [4-1:0] node20940;
	wire [4-1:0] node20941;
	wire [4-1:0] node20943;
	wire [4-1:0] node20946;
	wire [4-1:0] node20947;
	wire [4-1:0] node20951;
	wire [4-1:0] node20952;
	wire [4-1:0] node20953;
	wire [4-1:0] node20954;
	wire [4-1:0] node20955;
	wire [4-1:0] node20961;
	wire [4-1:0] node20962;
	wire [4-1:0] node20963;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20977;
	wire [4-1:0] node20978;
	wire [4-1:0] node20979;
	wire [4-1:0] node20980;
	wire [4-1:0] node20981;
	wire [4-1:0] node20982;
	wire [4-1:0] node20983;
	wire [4-1:0] node20987;
	wire [4-1:0] node20989;
	wire [4-1:0] node20991;
	wire [4-1:0] node20994;
	wire [4-1:0] node20995;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21001;
	wire [4-1:0] node21002;
	wire [4-1:0] node21006;
	wire [4-1:0] node21009;
	wire [4-1:0] node21010;
	wire [4-1:0] node21012;
	wire [4-1:0] node21013;
	wire [4-1:0] node21016;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21024;
	wire [4-1:0] node21025;
	wire [4-1:0] node21026;
	wire [4-1:0] node21028;
	wire [4-1:0] node21029;
	wire [4-1:0] node21032;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21038;
	wire [4-1:0] node21042;
	wire [4-1:0] node21043;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21049;
	wire [4-1:0] node21052;
	wire [4-1:0] node21053;
	wire [4-1:0] node21055;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21061;
	wire [4-1:0] node21064;
	wire [4-1:0] node21066;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21073;
	wire [4-1:0] node21074;
	wire [4-1:0] node21075;
	wire [4-1:0] node21078;
	wire [4-1:0] node21083;
	wire [4-1:0] node21084;
	wire [4-1:0] node21085;
	wire [4-1:0] node21089;
	wire [4-1:0] node21090;
	wire [4-1:0] node21091;
	wire [4-1:0] node21095;
	wire [4-1:0] node21097;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21107;
	wire [4-1:0] node21109;
	wire [4-1:0] node21112;
	wire [4-1:0] node21113;
	wire [4-1:0] node21116;
	wire [4-1:0] node21119;
	wire [4-1:0] node21120;
	wire [4-1:0] node21121;
	wire [4-1:0] node21123;
	wire [4-1:0] node21124;
	wire [4-1:0] node21128;
	wire [4-1:0] node21129;
	wire [4-1:0] node21131;
	wire [4-1:0] node21134;
	wire [4-1:0] node21136;
	wire [4-1:0] node21138;
	wire [4-1:0] node21141;
	wire [4-1:0] node21142;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21145;
	wire [4-1:0] node21150;
	wire [4-1:0] node21151;
	wire [4-1:0] node21152;
	wire [4-1:0] node21155;
	wire [4-1:0] node21159;
	wire [4-1:0] node21160;
	wire [4-1:0] node21163;
	wire [4-1:0] node21165;
	wire [4-1:0] node21166;
	wire [4-1:0] node21170;
	wire [4-1:0] node21171;
	wire [4-1:0] node21172;
	wire [4-1:0] node21173;
	wire [4-1:0] node21174;
	wire [4-1:0] node21175;
	wire [4-1:0] node21177;
	wire [4-1:0] node21178;
	wire [4-1:0] node21181;
	wire [4-1:0] node21185;
	wire [4-1:0] node21186;
	wire [4-1:0] node21187;
	wire [4-1:0] node21189;
	wire [4-1:0] node21192;
	wire [4-1:0] node21193;
	wire [4-1:0] node21196;
	wire [4-1:0] node21199;
	wire [4-1:0] node21202;
	wire [4-1:0] node21203;
	wire [4-1:0] node21204;
	wire [4-1:0] node21206;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21214;
	wire [4-1:0] node21215;
	wire [4-1:0] node21218;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21224;
	wire [4-1:0] node21225;
	wire [4-1:0] node21228;
	wire [4-1:0] node21231;
	wire [4-1:0] node21232;
	wire [4-1:0] node21235;
	wire [4-1:0] node21238;
	wire [4-1:0] node21239;
	wire [4-1:0] node21241;
	wire [4-1:0] node21245;
	wire [4-1:0] node21246;
	wire [4-1:0] node21248;
	wire [4-1:0] node21250;
	wire [4-1:0] node21253;
	wire [4-1:0] node21254;
	wire [4-1:0] node21255;
	wire [4-1:0] node21259;
	wire [4-1:0] node21260;
	wire [4-1:0] node21262;
	wire [4-1:0] node21266;
	wire [4-1:0] node21267;
	wire [4-1:0] node21268;
	wire [4-1:0] node21269;
	wire [4-1:0] node21270;
	wire [4-1:0] node21274;
	wire [4-1:0] node21275;
	wire [4-1:0] node21278;
	wire [4-1:0] node21281;
	wire [4-1:0] node21282;
	wire [4-1:0] node21283;
	wire [4-1:0] node21286;
	wire [4-1:0] node21290;
	wire [4-1:0] node21291;
	wire [4-1:0] node21292;
	wire [4-1:0] node21293;
	wire [4-1:0] node21295;
	wire [4-1:0] node21299;
	wire [4-1:0] node21301;
	wire [4-1:0] node21304;
	wire [4-1:0] node21305;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21310;
	wire [4-1:0] node21313;
	wire [4-1:0] node21316;
	wire [4-1:0] node21317;
	wire [4-1:0] node21318;
	wire [4-1:0] node21322;
	wire [4-1:0] node21323;
	wire [4-1:0] node21327;
	wire [4-1:0] node21328;
	wire [4-1:0] node21329;
	wire [4-1:0] node21330;
	wire [4-1:0] node21331;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21336;
	wire [4-1:0] node21339;
	wire [4-1:0] node21341;
	wire [4-1:0] node21343;
	wire [4-1:0] node21344;
	wire [4-1:0] node21347;
	wire [4-1:0] node21350;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21353;
	wire [4-1:0] node21354;
	wire [4-1:0] node21359;
	wire [4-1:0] node21361;
	wire [4-1:0] node21364;
	wire [4-1:0] node21366;
	wire [4-1:0] node21367;
	wire [4-1:0] node21369;
	wire [4-1:0] node21373;
	wire [4-1:0] node21374;
	wire [4-1:0] node21375;
	wire [4-1:0] node21377;
	wire [4-1:0] node21379;
	wire [4-1:0] node21382;
	wire [4-1:0] node21383;
	wire [4-1:0] node21384;
	wire [4-1:0] node21388;
	wire [4-1:0] node21390;
	wire [4-1:0] node21392;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21399;
	wire [4-1:0] node21400;
	wire [4-1:0] node21402;
	wire [4-1:0] node21404;
	wire [4-1:0] node21408;
	wire [4-1:0] node21409;
	wire [4-1:0] node21410;
	wire [4-1:0] node21411;
	wire [4-1:0] node21412;
	wire [4-1:0] node21413;
	wire [4-1:0] node21416;
	wire [4-1:0] node21420;
	wire [4-1:0] node21421;
	wire [4-1:0] node21422;
	wire [4-1:0] node21426;
	wire [4-1:0] node21429;
	wire [4-1:0] node21430;
	wire [4-1:0] node21432;
	wire [4-1:0] node21433;
	wire [4-1:0] node21437;
	wire [4-1:0] node21439;
	wire [4-1:0] node21442;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21445;
	wire [4-1:0] node21448;
	wire [4-1:0] node21449;
	wire [4-1:0] node21453;
	wire [4-1:0] node21455;
	wire [4-1:0] node21456;
	wire [4-1:0] node21457;
	wire [4-1:0] node21462;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21469;
	wire [4-1:0] node21470;
	wire [4-1:0] node21473;
	wire [4-1:0] node21476;
	wire [4-1:0] node21478;
	wire [4-1:0] node21481;
	wire [4-1:0] node21482;
	wire [4-1:0] node21483;
	wire [4-1:0] node21484;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21487;
	wire [4-1:0] node21488;
	wire [4-1:0] node21492;
	wire [4-1:0] node21493;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21510;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21518;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21523;
	wire [4-1:0] node21527;
	wire [4-1:0] node21528;
	wire [4-1:0] node21530;
	wire [4-1:0] node21533;
	wire [4-1:0] node21535;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21542;
	wire [4-1:0] node21544;
	wire [4-1:0] node21545;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21552;
	wire [4-1:0] node21553;
	wire [4-1:0] node21557;
	wire [4-1:0] node21559;
	wire [4-1:0] node21560;
	wire [4-1:0] node21564;
	wire [4-1:0] node21565;
	wire [4-1:0] node21566;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21571;
	wire [4-1:0] node21575;
	wire [4-1:0] node21576;
	wire [4-1:0] node21580;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21589;
	wire [4-1:0] node21593;
	wire [4-1:0] node21594;
	wire [4-1:0] node21596;
	wire [4-1:0] node21598;
	wire [4-1:0] node21602;
	wire [4-1:0] node21603;
	wire [4-1:0] node21604;
	wire [4-1:0] node21605;
	wire [4-1:0] node21608;
	wire [4-1:0] node21609;
	wire [4-1:0] node21613;
	wire [4-1:0] node21615;
	wire [4-1:0] node21617;
	wire [4-1:0] node21620;
	wire [4-1:0] node21623;
	wire [4-1:0] node21624;
	wire [4-1:0] node21625;
	wire [4-1:0] node21627;
	wire [4-1:0] node21628;
	wire [4-1:0] node21630;
	wire [4-1:0] node21633;
	wire [4-1:0] node21636;
	wire [4-1:0] node21637;
	wire [4-1:0] node21639;
	wire [4-1:0] node21640;
	wire [4-1:0] node21643;
	wire [4-1:0] node21646;
	wire [4-1:0] node21647;
	wire [4-1:0] node21651;
	wire [4-1:0] node21652;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21656;
	wire [4-1:0] node21659;
	wire [4-1:0] node21662;
	wire [4-1:0] node21663;
	wire [4-1:0] node21667;
	wire [4-1:0] node21668;
	wire [4-1:0] node21669;
	wire [4-1:0] node21673;
	wire [4-1:0] node21674;
	wire [4-1:0] node21677;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21683;
	wire [4-1:0] node21684;
	wire [4-1:0] node21685;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21689;
	wire [4-1:0] node21692;
	wire [4-1:0] node21694;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21701;
	wire [4-1:0] node21704;
	wire [4-1:0] node21705;
	wire [4-1:0] node21708;
	wire [4-1:0] node21711;
	wire [4-1:0] node21712;
	wire [4-1:0] node21713;
	wire [4-1:0] node21715;
	wire [4-1:0] node21719;
	wire [4-1:0] node21720;
	wire [4-1:0] node21722;
	wire [4-1:0] node21725;
	wire [4-1:0] node21727;
	wire [4-1:0] node21728;
	wire [4-1:0] node21731;
	wire [4-1:0] node21734;
	wire [4-1:0] node21735;
	wire [4-1:0] node21736;
	wire [4-1:0] node21739;
	wire [4-1:0] node21740;
	wire [4-1:0] node21741;
	wire [4-1:0] node21742;
	wire [4-1:0] node21745;
	wire [4-1:0] node21748;
	wire [4-1:0] node21750;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21756;
	wire [4-1:0] node21757;
	wire [4-1:0] node21761;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21768;
	wire [4-1:0] node21769;
	wire [4-1:0] node21770;
	wire [4-1:0] node21774;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21779;
	wire [4-1:0] node21780;
	wire [4-1:0] node21781;
	wire [4-1:0] node21783;
	wire [4-1:0] node21786;
	wire [4-1:0] node21788;
	wire [4-1:0] node21791;
	wire [4-1:0] node21792;
	wire [4-1:0] node21793;
	wire [4-1:0] node21796;
	wire [4-1:0] node21800;
	wire [4-1:0] node21801;
	wire [4-1:0] node21803;
	wire [4-1:0] node21805;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21810;
	wire [4-1:0] node21811;
	wire [4-1:0] node21814;
	wire [4-1:0] node21819;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21823;
	wire [4-1:0] node21826;
	wire [4-1:0] node21829;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21838;
	wire [4-1:0] node21839;
	wire [4-1:0] node21842;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21849;
	wire [4-1:0] node21853;
	wire [4-1:0] node21855;
	wire [4-1:0] node21856;
	wire [4-1:0] node21858;
	wire [4-1:0] node21862;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21865;
	wire [4-1:0] node21866;
	wire [4-1:0] node21868;
	wire [4-1:0] node21870;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21875;
	wire [4-1:0] node21879;
	wire [4-1:0] node21880;
	wire [4-1:0] node21881;
	wire [4-1:0] node21884;
	wire [4-1:0] node21887;
	wire [4-1:0] node21888;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21899;
	wire [4-1:0] node21902;
	wire [4-1:0] node21904;
	wire [4-1:0] node21905;
	wire [4-1:0] node21909;
	wire [4-1:0] node21910;
	wire [4-1:0] node21911;
	wire [4-1:0] node21912;
	wire [4-1:0] node21915;
	wire [4-1:0] node21918;
	wire [4-1:0] node21919;
	wire [4-1:0] node21920;
	wire [4-1:0] node21923;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21931;
	wire [4-1:0] node21932;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21939;
	wire [4-1:0] node21943;
	wire [4-1:0] node21944;
	wire [4-1:0] node21945;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21954;
	wire [4-1:0] node21957;
	wire [4-1:0] node21958;
	wire [4-1:0] node21961;
	wire [4-1:0] node21964;
	wire [4-1:0] node21965;
	wire [4-1:0] node21966;
	wire [4-1:0] node21967;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21970;
	wire [4-1:0] node21973;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21981;
	wire [4-1:0] node21983;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21990;
	wire [4-1:0] node21993;
	wire [4-1:0] node21994;
	wire [4-1:0] node21995;
	wire [4-1:0] node21998;
	wire [4-1:0] node22001;
	wire [4-1:0] node22002;
	wire [4-1:0] node22003;
	wire [4-1:0] node22006;
	wire [4-1:0] node22009;
	wire [4-1:0] node22010;
	wire [4-1:0] node22013;
	wire [4-1:0] node22016;
	wire [4-1:0] node22017;
	wire [4-1:0] node22019;
	wire [4-1:0] node22020;
	wire [4-1:0] node22021;
	wire [4-1:0] node22024;
	wire [4-1:0] node22027;
	wire [4-1:0] node22028;
	wire [4-1:0] node22032;
	wire [4-1:0] node22033;
	wire [4-1:0] node22034;
	wire [4-1:0] node22035;
	wire [4-1:0] node22036;
	wire [4-1:0] node22039;
	wire [4-1:0] node22044;
	wire [4-1:0] node22045;
	wire [4-1:0] node22046;
	wire [4-1:0] node22051;
	wire [4-1:0] node22052;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22056;
	wire [4-1:0] node22057;
	wire [4-1:0] node22059;
	wire [4-1:0] node22060;
	wire [4-1:0] node22061;
	wire [4-1:0] node22064;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22073;
	wire [4-1:0] node22074;
	wire [4-1:0] node22075;
	wire [4-1:0] node22077;
	wire [4-1:0] node22080;
	wire [4-1:0] node22082;
	wire [4-1:0] node22084;
	wire [4-1:0] node22087;
	wire [4-1:0] node22088;
	wire [4-1:0] node22089;
	wire [4-1:0] node22090;
	wire [4-1:0] node22093;
	wire [4-1:0] node22096;
	wire [4-1:0] node22098;
	wire [4-1:0] node22101;
	wire [4-1:0] node22102;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22108;
	wire [4-1:0] node22109;
	wire [4-1:0] node22110;
	wire [4-1:0] node22113;
	wire [4-1:0] node22117;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22123;
	wire [4-1:0] node22124;
	wire [4-1:0] node22125;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22132;
	wire [4-1:0] node22136;
	wire [4-1:0] node22138;
	wire [4-1:0] node22140;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22145;
	wire [4-1:0] node22146;
	wire [4-1:0] node22147;
	wire [4-1:0] node22148;
	wire [4-1:0] node22149;
	wire [4-1:0] node22152;
	wire [4-1:0] node22156;
	wire [4-1:0] node22157;
	wire [4-1:0] node22158;
	wire [4-1:0] node22161;
	wire [4-1:0] node22165;
	wire [4-1:0] node22166;
	wire [4-1:0] node22170;
	wire [4-1:0] node22171;
	wire [4-1:0] node22172;
	wire [4-1:0] node22175;
	wire [4-1:0] node22177;
	wire [4-1:0] node22180;
	wire [4-1:0] node22182;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22188;
	wire [4-1:0] node22189;
	wire [4-1:0] node22193;
	wire [4-1:0] node22195;
	wire [4-1:0] node22197;
	wire [4-1:0] node22200;
	wire [4-1:0] node22202;
	wire [4-1:0] node22203;
	wire [4-1:0] node22206;
	wire [4-1:0] node22209;
	wire [4-1:0] node22210;
	wire [4-1:0] node22211;
	wire [4-1:0] node22212;
	wire [4-1:0] node22214;
	wire [4-1:0] node22217;
	wire [4-1:0] node22219;
	wire [4-1:0] node22223;
	wire [4-1:0] node22224;
	wire [4-1:0] node22225;
	wire [4-1:0] node22226;
	wire [4-1:0] node22231;
	wire [4-1:0] node22232;
	wire [4-1:0] node22236;
	wire [4-1:0] node22237;
	wire [4-1:0] node22238;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22242;
	wire [4-1:0] node22244;
	wire [4-1:0] node22247;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22252;
	wire [4-1:0] node22254;
	wire [4-1:0] node22258;
	wire [4-1:0] node22259;
	wire [4-1:0] node22260;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22266;
	wire [4-1:0] node22268;
	wire [4-1:0] node22271;
	wire [4-1:0] node22272;
	wire [4-1:0] node22276;
	wire [4-1:0] node22278;
	wire [4-1:0] node22281;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22284;
	wire [4-1:0] node22286;
	wire [4-1:0] node22289;
	wire [4-1:0] node22291;
	wire [4-1:0] node22292;
	wire [4-1:0] node22296;
	wire [4-1:0] node22297;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22303;
	wire [4-1:0] node22307;
	wire [4-1:0] node22308;
	wire [4-1:0] node22309;
	wire [4-1:0] node22311;
	wire [4-1:0] node22312;
	wire [4-1:0] node22316;
	wire [4-1:0] node22317;
	wire [4-1:0] node22318;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22325;
	wire [4-1:0] node22329;
	wire [4-1:0] node22330;
	wire [4-1:0] node22332;
	wire [4-1:0] node22336;
	wire [4-1:0] node22337;
	wire [4-1:0] node22338;
	wire [4-1:0] node22339;
	wire [4-1:0] node22340;
	wire [4-1:0] node22341;
	wire [4-1:0] node22346;
	wire [4-1:0] node22347;
	wire [4-1:0] node22348;
	wire [4-1:0] node22349;
	wire [4-1:0] node22352;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22361;
	wire [4-1:0] node22362;
	wire [4-1:0] node22366;
	wire [4-1:0] node22367;
	wire [4-1:0] node22371;
	wire [4-1:0] node22373;
	wire [4-1:0] node22374;
	wire [4-1:0] node22376;
	wire [4-1:0] node22380;
	wire [4-1:0] node22381;
	wire [4-1:0] node22382;
	wire [4-1:0] node22383;
	wire [4-1:0] node22385;
	wire [4-1:0] node22389;
	wire [4-1:0] node22390;
	wire [4-1:0] node22393;
	wire [4-1:0] node22395;
	wire [4-1:0] node22396;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22402;
	wire [4-1:0] node22403;
	wire [4-1:0] node22406;
	wire [4-1:0] node22410;
	wire [4-1:0] node22412;
	wire [4-1:0] node22414;
	wire [4-1:0] node22415;
	wire [4-1:0] node22419;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22423;
	wire [4-1:0] node22424;
	wire [4-1:0] node22425;
	wire [4-1:0] node22426;
	wire [4-1:0] node22429;
	wire [4-1:0] node22432;
	wire [4-1:0] node22433;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22440;
	wire [4-1:0] node22443;
	wire [4-1:0] node22444;
	wire [4-1:0] node22447;
	wire [4-1:0] node22450;
	wire [4-1:0] node22451;
	wire [4-1:0] node22452;
	wire [4-1:0] node22454;
	wire [4-1:0] node22457;
	wire [4-1:0] node22460;
	wire [4-1:0] node22461;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22466;
	wire [4-1:0] node22470;
	wire [4-1:0] node22471;
	wire [4-1:0] node22472;
	wire [4-1:0] node22475;
	wire [4-1:0] node22478;
	wire [4-1:0] node22479;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22485;
	wire [4-1:0] node22486;
	wire [4-1:0] node22487;
	wire [4-1:0] node22489;
	wire [4-1:0] node22493;
	wire [4-1:0] node22494;
	wire [4-1:0] node22497;
	wire [4-1:0] node22498;
	wire [4-1:0] node22502;
	wire [4-1:0] node22503;
	wire [4-1:0] node22507;
	wire [4-1:0] node22508;
	wire [4-1:0] node22509;
	wire [4-1:0] node22511;
	wire [4-1:0] node22512;
	wire [4-1:0] node22516;
	wire [4-1:0] node22517;
	wire [4-1:0] node22521;
	wire [4-1:0] node22522;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22529;
	wire [4-1:0] node22531;
	wire [4-1:0] node22534;
	wire [4-1:0] node22535;
	wire [4-1:0] node22536;
	wire [4-1:0] node22537;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22540;
	wire [4-1:0] node22546;
	wire [4-1:0] node22547;
	wire [4-1:0] node22548;
	wire [4-1:0] node22553;
	wire [4-1:0] node22554;
	wire [4-1:0] node22555;
	wire [4-1:0] node22557;
	wire [4-1:0] node22558;
	wire [4-1:0] node22562;
	wire [4-1:0] node22563;
	wire [4-1:0] node22565;
	wire [4-1:0] node22569;
	wire [4-1:0] node22570;
	wire [4-1:0] node22571;
	wire [4-1:0] node22575;
	wire [4-1:0] node22578;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22581;
	wire [4-1:0] node22582;
	wire [4-1:0] node22586;
	wire [4-1:0] node22589;
	wire [4-1:0] node22590;
	wire [4-1:0] node22592;
	wire [4-1:0] node22596;
	wire [4-1:0] node22597;
	wire [4-1:0] node22599;
	wire [4-1:0] node22601;
	wire [4-1:0] node22602;
	wire [4-1:0] node22606;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22610;
	wire [4-1:0] node22613;
	wire [4-1:0] node22617;
	wire [4-1:0] node22618;
	wire [4-1:0] node22619;
	wire [4-1:0] node22620;
	wire [4-1:0] node22621;
	wire [4-1:0] node22623;
	wire [4-1:0] node22626;
	wire [4-1:0] node22627;
	wire [4-1:0] node22628;
	wire [4-1:0] node22630;
	wire [4-1:0] node22635;
	wire [4-1:0] node22636;
	wire [4-1:0] node22638;
	wire [4-1:0] node22641;
	wire [4-1:0] node22643;
	wire [4-1:0] node22645;
	wire [4-1:0] node22648;
	wire [4-1:0] node22649;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22655;
	wire [4-1:0] node22657;
	wire [4-1:0] node22658;
	wire [4-1:0] node22661;
	wire [4-1:0] node22664;
	wire [4-1:0] node22665;
	wire [4-1:0] node22666;
	wire [4-1:0] node22668;
	wire [4-1:0] node22671;
	wire [4-1:0] node22672;
	wire [4-1:0] node22674;
	wire [4-1:0] node22678;
	wire [4-1:0] node22679;
	wire [4-1:0] node22680;
	wire [4-1:0] node22682;
	wire [4-1:0] node22685;
	wire [4-1:0] node22688;
	wire [4-1:0] node22689;
	wire [4-1:0] node22693;
	wire [4-1:0] node22694;
	wire [4-1:0] node22695;
	wire [4-1:0] node22696;
	wire [4-1:0] node22697;
	wire [4-1:0] node22698;
	wire [4-1:0] node22701;
	wire [4-1:0] node22705;
	wire [4-1:0] node22706;
	wire [4-1:0] node22707;
	wire [4-1:0] node22710;
	wire [4-1:0] node22714;
	wire [4-1:0] node22715;
	wire [4-1:0] node22717;
	wire [4-1:0] node22720;
	wire [4-1:0] node22721;
	wire [4-1:0] node22724;
	wire [4-1:0] node22727;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22731;
	wire [4-1:0] node22735;
	wire [4-1:0] node22737;
	wire [4-1:0] node22740;
	wire [4-1:0] node22742;
	wire [4-1:0] node22745;
	wire [4-1:0] node22746;
	wire [4-1:0] node22747;
	wire [4-1:0] node22748;
	wire [4-1:0] node22751;
	wire [4-1:0] node22755;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22760;
	wire [4-1:0] node22761;
	wire [4-1:0] node22762;
	wire [4-1:0] node22763;
	wire [4-1:0] node22764;
	wire [4-1:0] node22765;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22771;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22779;
	wire [4-1:0] node22782;
	wire [4-1:0] node22783;
	wire [4-1:0] node22785;
	wire [4-1:0] node22786;
	wire [4-1:0] node22787;
	wire [4-1:0] node22790;
	wire [4-1:0] node22794;
	wire [4-1:0] node22796;
	wire [4-1:0] node22797;
	wire [4-1:0] node22800;
	wire [4-1:0] node22803;
	wire [4-1:0] node22804;
	wire [4-1:0] node22805;
	wire [4-1:0] node22806;
	wire [4-1:0] node22810;
	wire [4-1:0] node22812;
	wire [4-1:0] node22813;
	wire [4-1:0] node22816;
	wire [4-1:0] node22819;
	wire [4-1:0] node22820;
	wire [4-1:0] node22821;
	wire [4-1:0] node22823;
	wire [4-1:0] node22827;
	wire [4-1:0] node22829;
	wire [4-1:0] node22831;
	wire [4-1:0] node22832;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22838;
	wire [4-1:0] node22839;
	wire [4-1:0] node22840;
	wire [4-1:0] node22841;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22849;
	wire [4-1:0] node22852;
	wire [4-1:0] node22855;
	wire [4-1:0] node22856;
	wire [4-1:0] node22857;
	wire [4-1:0] node22858;
	wire [4-1:0] node22859;
	wire [4-1:0] node22863;
	wire [4-1:0] node22864;
	wire [4-1:0] node22867;
	wire [4-1:0] node22870;
	wire [4-1:0] node22872;
	wire [4-1:0] node22875;
	wire [4-1:0] node22876;
	wire [4-1:0] node22877;
	wire [4-1:0] node22881;
	wire [4-1:0] node22883;
	wire [4-1:0] node22886;
	wire [4-1:0] node22887;
	wire [4-1:0] node22888;
	wire [4-1:0] node22890;
	wire [4-1:0] node22891;
	wire [4-1:0] node22894;
	wire [4-1:0] node22897;
	wire [4-1:0] node22898;
	wire [4-1:0] node22899;
	wire [4-1:0] node22902;
	wire [4-1:0] node22906;
	wire [4-1:0] node22907;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22911;
	wire [4-1:0] node22914;
	wire [4-1:0] node22917;
	wire [4-1:0] node22919;
	wire [4-1:0] node22922;
	wire [4-1:0] node22923;
	wire [4-1:0] node22924;
	wire [4-1:0] node22927;
	wire [4-1:0] node22930;
	wire [4-1:0] node22932;
	wire [4-1:0] node22933;
	wire [4-1:0] node22937;
	wire [4-1:0] node22938;
	wire [4-1:0] node22939;
	wire [4-1:0] node22940;
	wire [4-1:0] node22941;
	wire [4-1:0] node22942;
	wire [4-1:0] node22944;
	wire [4-1:0] node22947;
	wire [4-1:0] node22949;
	wire [4-1:0] node22951;
	wire [4-1:0] node22954;
	wire [4-1:0] node22955;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22960;
	wire [4-1:0] node22964;
	wire [4-1:0] node22965;
	wire [4-1:0] node22967;
	wire [4-1:0] node22970;
	wire [4-1:0] node22973;
	wire [4-1:0] node22974;
	wire [4-1:0] node22975;
	wire [4-1:0] node22976;
	wire [4-1:0] node22980;
	wire [4-1:0] node22981;
	wire [4-1:0] node22985;
	wire [4-1:0] node22987;
	wire [4-1:0] node22988;
	wire [4-1:0] node22989;
	wire [4-1:0] node22992;
	wire [4-1:0] node22996;
	wire [4-1:0] node22997;
	wire [4-1:0] node22998;
	wire [4-1:0] node22999;
	wire [4-1:0] node23002;
	wire [4-1:0] node23004;
	wire [4-1:0] node23007;
	wire [4-1:0] node23008;
	wire [4-1:0] node23009;
	wire [4-1:0] node23010;
	wire [4-1:0] node23013;
	wire [4-1:0] node23017;
	wire [4-1:0] node23018;
	wire [4-1:0] node23022;
	wire [4-1:0] node23023;
	wire [4-1:0] node23024;
	wire [4-1:0] node23025;
	wire [4-1:0] node23029;
	wire [4-1:0] node23030;
	wire [4-1:0] node23034;
	wire [4-1:0] node23035;
	wire [4-1:0] node23036;
	wire [4-1:0] node23041;
	wire [4-1:0] node23042;
	wire [4-1:0] node23043;
	wire [4-1:0] node23044;
	wire [4-1:0] node23045;
	wire [4-1:0] node23047;
	wire [4-1:0] node23050;
	wire [4-1:0] node23051;
	wire [4-1:0] node23052;
	wire [4-1:0] node23056;
	wire [4-1:0] node23057;
	wire [4-1:0] node23061;
	wire [4-1:0] node23062;
	wire [4-1:0] node23063;
	wire [4-1:0] node23064;
	wire [4-1:0] node23067;
	wire [4-1:0] node23071;
	wire [4-1:0] node23072;
	wire [4-1:0] node23076;
	wire [4-1:0] node23077;
	wire [4-1:0] node23079;
	wire [4-1:0] node23080;
	wire [4-1:0] node23081;
	wire [4-1:0] node23084;
	wire [4-1:0] node23088;
	wire [4-1:0] node23090;
	wire [4-1:0] node23091;
	wire [4-1:0] node23093;
	wire [4-1:0] node23096;
	wire [4-1:0] node23099;
	wire [4-1:0] node23100;
	wire [4-1:0] node23101;
	wire [4-1:0] node23102;
	wire [4-1:0] node23105;
	wire [4-1:0] node23106;
	wire [4-1:0] node23107;
	wire [4-1:0] node23111;
	wire [4-1:0] node23113;
	wire [4-1:0] node23116;
	wire [4-1:0] node23118;
	wire [4-1:0] node23119;
	wire [4-1:0] node23122;
	wire [4-1:0] node23125;
	wire [4-1:0] node23126;
	wire [4-1:0] node23127;
	wire [4-1:0] node23128;
	wire [4-1:0] node23131;
	wire [4-1:0] node23133;
	wire [4-1:0] node23136;
	wire [4-1:0] node23138;
	wire [4-1:0] node23141;
	wire [4-1:0] node23142;
	wire [4-1:0] node23144;
	wire [4-1:0] node23146;
	wire [4-1:0] node23149;
	wire [4-1:0] node23152;
	wire [4-1:0] node23153;
	wire [4-1:0] node23154;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23159;
	wire [4-1:0] node23162;
	wire [4-1:0] node23163;
	wire [4-1:0] node23166;
	wire [4-1:0] node23169;
	wire [4-1:0] node23170;
	wire [4-1:0] node23171;
	wire [4-1:0] node23172;
	wire [4-1:0] node23176;
	wire [4-1:0] node23177;
	wire [4-1:0] node23181;
	wire [4-1:0] node23182;
	wire [4-1:0] node23183;
	wire [4-1:0] node23186;
	wire [4-1:0] node23189;
	wire [4-1:0] node23191;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23196;
	wire [4-1:0] node23197;
	wire [4-1:0] node23199;
	wire [4-1:0] node23203;
	wire [4-1:0] node23205;
	wire [4-1:0] node23208;
	wire [4-1:0] node23209;
	wire [4-1:0] node23210;
	wire [4-1:0] node23211;
	wire [4-1:0] node23212;
	wire [4-1:0] node23215;
	wire [4-1:0] node23219;
	wire [4-1:0] node23221;
	wire [4-1:0] node23223;
	wire [4-1:0] node23226;
	wire [4-1:0] node23229;
	wire [4-1:0] node23230;
	wire [4-1:0] node23231;
	wire [4-1:0] node23232;
	wire [4-1:0] node23233;
	wire [4-1:0] node23236;
	wire [4-1:0] node23239;
	wire [4-1:0] node23240;
	wire [4-1:0] node23241;
	wire [4-1:0] node23244;
	wire [4-1:0] node23246;
	wire [4-1:0] node23250;
	wire [4-1:0] node23251;
	wire [4-1:0] node23252;
	wire [4-1:0] node23253;
	wire [4-1:0] node23254;
	wire [4-1:0] node23258;
	wire [4-1:0] node23260;
	wire [4-1:0] node23263;
	wire [4-1:0] node23266;
	wire [4-1:0] node23267;
	wire [4-1:0] node23268;
	wire [4-1:0] node23272;
	wire [4-1:0] node23273;
	wire [4-1:0] node23276;
	wire [4-1:0] node23279;
	wire [4-1:0] node23280;
	wire [4-1:0] node23281;
	wire [4-1:0] node23283;
	wire [4-1:0] node23285;
	wire [4-1:0] node23287;
	wire [4-1:0] node23290;
	wire [4-1:0] node23292;
	wire [4-1:0] node23294;
	wire [4-1:0] node23295;
	wire [4-1:0] node23299;
	wire [4-1:0] node23300;
	wire [4-1:0] node23301;
	wire [4-1:0] node23303;
	wire [4-1:0] node23306;
	wire [4-1:0] node23307;
	wire [4-1:0] node23310;
	wire [4-1:0] node23313;
	wire [4-1:0] node23314;
	wire [4-1:0] node23316;
	wire [4-1:0] node23320;
	wire [4-1:0] node23321;
	wire [4-1:0] node23322;
	wire [4-1:0] node23323;
	wire [4-1:0] node23324;
	wire [4-1:0] node23326;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23332;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23338;
	wire [4-1:0] node23341;
	wire [4-1:0] node23343;
	wire [4-1:0] node23346;
	wire [4-1:0] node23347;
	wire [4-1:0] node23348;
	wire [4-1:0] node23349;
	wire [4-1:0] node23353;
	wire [4-1:0] node23354;
	wire [4-1:0] node23355;
	wire [4-1:0] node23358;
	wire [4-1:0] node23362;
	wire [4-1:0] node23363;
	wire [4-1:0] node23367;
	wire [4-1:0] node23368;
	wire [4-1:0] node23369;
	wire [4-1:0] node23370;
	wire [4-1:0] node23371;
	wire [4-1:0] node23372;
	wire [4-1:0] node23375;
	wire [4-1:0] node23380;
	wire [4-1:0] node23381;
	wire [4-1:0] node23382;
	wire [4-1:0] node23387;
	wire [4-1:0] node23388;
	wire [4-1:0] node23389;
	wire [4-1:0] node23391;
	wire [4-1:0] node23394;
	wire [4-1:0] node23395;
	wire [4-1:0] node23399;
	wire [4-1:0] node23400;
	wire [4-1:0] node23401;
	wire [4-1:0] node23403;
	wire [4-1:0] node23406;
	wire [4-1:0] node23408;
	wire [4-1:0] node23411;
	wire [4-1:0] node23413;
	wire [4-1:0] node23416;
	wire [4-1:0] node23417;
	wire [4-1:0] node23418;
	wire [4-1:0] node23420;
	wire [4-1:0] node23421;
	wire [4-1:0] node23423;
	wire [4-1:0] node23426;
	wire [4-1:0] node23428;
	wire [4-1:0] node23431;
	wire [4-1:0] node23433;
	wire [4-1:0] node23436;
	wire [4-1:0] node23437;
	wire [4-1:0] node23438;
	wire [4-1:0] node23440;
	wire [4-1:0] node23443;
	wire [4-1:0] node23445;
	wire [4-1:0] node23448;
	wire [4-1:0] node23449;
	wire [4-1:0] node23451;
	wire [4-1:0] node23454;
	wire [4-1:0] node23456;
	wire [4-1:0] node23459;
	wire [4-1:0] node23460;
	wire [4-1:0] node23461;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23464;
	wire [4-1:0] node23465;
	wire [4-1:0] node23466;
	wire [4-1:0] node23469;
	wire [4-1:0] node23472;
	wire [4-1:0] node23473;
	wire [4-1:0] node23474;
	wire [4-1:0] node23475;
	wire [4-1:0] node23479;
	wire [4-1:0] node23480;
	wire [4-1:0] node23483;
	wire [4-1:0] node23486;
	wire [4-1:0] node23488;
	wire [4-1:0] node23491;
	wire [4-1:0] node23492;
	wire [4-1:0] node23493;
	wire [4-1:0] node23495;
	wire [4-1:0] node23498;
	wire [4-1:0] node23501;
	wire [4-1:0] node23502;
	wire [4-1:0] node23504;
	wire [4-1:0] node23506;
	wire [4-1:0] node23510;
	wire [4-1:0] node23511;
	wire [4-1:0] node23512;
	wire [4-1:0] node23513;
	wire [4-1:0] node23514;
	wire [4-1:0] node23517;
	wire [4-1:0] node23521;
	wire [4-1:0] node23522;
	wire [4-1:0] node23523;
	wire [4-1:0] node23524;
	wire [4-1:0] node23528;
	wire [4-1:0] node23529;
	wire [4-1:0] node23534;
	wire [4-1:0] node23535;
	wire [4-1:0] node23536;
	wire [4-1:0] node23537;
	wire [4-1:0] node23541;
	wire [4-1:0] node23542;
	wire [4-1:0] node23546;
	wire [4-1:0] node23547;
	wire [4-1:0] node23550;
	wire [4-1:0] node23551;
	wire [4-1:0] node23555;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23559;
	wire [4-1:0] node23560;
	wire [4-1:0] node23564;
	wire [4-1:0] node23565;
	wire [4-1:0] node23569;
	wire [4-1:0] node23571;
	wire [4-1:0] node23574;
	wire [4-1:0] node23575;
	wire [4-1:0] node23576;
	wire [4-1:0] node23578;
	wire [4-1:0] node23582;
	wire [4-1:0] node23583;
	wire [4-1:0] node23584;
	wire [4-1:0] node23585;
	wire [4-1:0] node23588;
	wire [4-1:0] node23593;
	wire [4-1:0] node23594;
	wire [4-1:0] node23595;
	wire [4-1:0] node23596;
	wire [4-1:0] node23599;
	wire [4-1:0] node23601;
	wire [4-1:0] node23602;
	wire [4-1:0] node23605;
	wire [4-1:0] node23608;
	wire [4-1:0] node23611;
	wire [4-1:0] node23612;
	wire [4-1:0] node23613;
	wire [4-1:0] node23616;
	wire [4-1:0] node23617;
	wire [4-1:0] node23620;
	wire [4-1:0] node23623;
	wire [4-1:0] node23625;
	wire [4-1:0] node23627;
	wire [4-1:0] node23630;
	wire [4-1:0] node23631;
	wire [4-1:0] node23632;
	wire [4-1:0] node23633;
	wire [4-1:0] node23634;
	wire [4-1:0] node23635;
	wire [4-1:0] node23636;
	wire [4-1:0] node23638;
	wire [4-1:0] node23643;
	wire [4-1:0] node23645;
	wire [4-1:0] node23647;
	wire [4-1:0] node23649;
	wire [4-1:0] node23652;
	wire [4-1:0] node23653;
	wire [4-1:0] node23654;
	wire [4-1:0] node23657;
	wire [4-1:0] node23659;
	wire [4-1:0] node23662;
	wire [4-1:0] node23663;
	wire [4-1:0] node23664;
	wire [4-1:0] node23668;
	wire [4-1:0] node23669;
	wire [4-1:0] node23672;
	wire [4-1:0] node23675;
	wire [4-1:0] node23676;
	wire [4-1:0] node23677;
	wire [4-1:0] node23678;
	wire [4-1:0] node23679;
	wire [4-1:0] node23683;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23690;
	wire [4-1:0] node23692;
	wire [4-1:0] node23694;
	wire [4-1:0] node23695;
	wire [4-1:0] node23698;
	wire [4-1:0] node23701;
	wire [4-1:0] node23702;
	wire [4-1:0] node23703;
	wire [4-1:0] node23704;
	wire [4-1:0] node23708;
	wire [4-1:0] node23709;
	wire [4-1:0] node23713;
	wire [4-1:0] node23714;
	wire [4-1:0] node23715;
	wire [4-1:0] node23720;
	wire [4-1:0] node23721;
	wire [4-1:0] node23722;
	wire [4-1:0] node23723;
	wire [4-1:0] node23724;
	wire [4-1:0] node23727;
	wire [4-1:0] node23728;
	wire [4-1:0] node23730;
	wire [4-1:0] node23734;
	wire [4-1:0] node23736;
	wire [4-1:0] node23737;
	wire [4-1:0] node23738;
	wire [4-1:0] node23743;
	wire [4-1:0] node23744;
	wire [4-1:0] node23745;
	wire [4-1:0] node23747;
	wire [4-1:0] node23750;
	wire [4-1:0] node23751;
	wire [4-1:0] node23755;
	wire [4-1:0] node23756;
	wire [4-1:0] node23758;
	wire [4-1:0] node23761;
	wire [4-1:0] node23763;
	wire [4-1:0] node23764;
	wire [4-1:0] node23767;
	wire [4-1:0] node23770;
	wire [4-1:0] node23771;
	wire [4-1:0] node23772;
	wire [4-1:0] node23774;
	wire [4-1:0] node23775;
	wire [4-1:0] node23779;
	wire [4-1:0] node23781;
	wire [4-1:0] node23782;
	wire [4-1:0] node23786;
	wire [4-1:0] node23787;
	wire [4-1:0] node23788;
	wire [4-1:0] node23789;
	wire [4-1:0] node23791;
	wire [4-1:0] node23795;
	wire [4-1:0] node23796;
	wire [4-1:0] node23800;
	wire [4-1:0] node23801;
	wire [4-1:0] node23802;
	wire [4-1:0] node23806;
	wire [4-1:0] node23807;
	wire [4-1:0] node23811;
	wire [4-1:0] node23812;
	wire [4-1:0] node23813;
	wire [4-1:0] node23814;
	wire [4-1:0] node23815;
	wire [4-1:0] node23816;
	wire [4-1:0] node23817;
	wire [4-1:0] node23818;
	wire [4-1:0] node23823;
	wire [4-1:0] node23824;
	wire [4-1:0] node23826;
	wire [4-1:0] node23828;
	wire [4-1:0] node23832;
	wire [4-1:0] node23833;
	wire [4-1:0] node23835;
	wire [4-1:0] node23836;
	wire [4-1:0] node23839;
	wire [4-1:0] node23842;
	wire [4-1:0] node23843;
	wire [4-1:0] node23845;
	wire [4-1:0] node23846;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23852;
	wire [4-1:0] node23855;
	wire [4-1:0] node23859;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23863;
	wire [4-1:0] node23864;
	wire [4-1:0] node23868;
	wire [4-1:0] node23870;
	wire [4-1:0] node23872;
	wire [4-1:0] node23873;
	wire [4-1:0] node23877;
	wire [4-1:0] node23878;
	wire [4-1:0] node23879;
	wire [4-1:0] node23880;
	wire [4-1:0] node23881;
	wire [4-1:0] node23887;
	wire [4-1:0] node23888;
	wire [4-1:0] node23890;
	wire [4-1:0] node23893;
	wire [4-1:0] node23895;
	wire [4-1:0] node23898;
	wire [4-1:0] node23899;
	wire [4-1:0] node23900;
	wire [4-1:0] node23901;
	wire [4-1:0] node23903;
	wire [4-1:0] node23904;
	wire [4-1:0] node23908;
	wire [4-1:0] node23909;
	wire [4-1:0] node23910;
	wire [4-1:0] node23912;
	wire [4-1:0] node23915;
	wire [4-1:0] node23918;
	wire [4-1:0] node23920;
	wire [4-1:0] node23923;
	wire [4-1:0] node23924;
	wire [4-1:0] node23926;
	wire [4-1:0] node23929;
	wire [4-1:0] node23930;
	wire [4-1:0] node23933;
	wire [4-1:0] node23936;
	wire [4-1:0] node23937;
	wire [4-1:0] node23938;
	wire [4-1:0] node23940;
	wire [4-1:0] node23943;
	wire [4-1:0] node23945;
	wire [4-1:0] node23946;
	wire [4-1:0] node23949;
	wire [4-1:0] node23952;
	wire [4-1:0] node23953;
	wire [4-1:0] node23955;
	wire [4-1:0] node23958;
	wire [4-1:0] node23959;
	wire [4-1:0] node23960;
	wire [4-1:0] node23964;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23970;
	wire [4-1:0] node23971;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23979;
	wire [4-1:0] node23983;
	wire [4-1:0] node23984;
	wire [4-1:0] node23985;
	wire [4-1:0] node23986;
	wire [4-1:0] node23987;
	wire [4-1:0] node23990;
	wire [4-1:0] node23996;
	wire [4-1:0] node23997;
	wire [4-1:0] node23998;
	wire [4-1:0] node24002;
	wire [4-1:0] node24003;
	wire [4-1:0] node24007;
	wire [4-1:0] node24008;
	wire [4-1:0] node24009;
	wire [4-1:0] node24010;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24023;
	wire [4-1:0] node24024;
	wire [4-1:0] node24025;
	wire [4-1:0] node24026;
	wire [4-1:0] node24027;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24034;
	wire [4-1:0] node24037;
	wire [4-1:0] node24041;
	wire [4-1:0] node24042;
	wire [4-1:0] node24046;
	wire [4-1:0] node24047;
	wire [4-1:0] node24048;
	wire [4-1:0] node24049;
	wire [4-1:0] node24050;
	wire [4-1:0] node24051;
	wire [4-1:0] node24052;
	wire [4-1:0] node24053;
	wire [4-1:0] node24054;
	wire [4-1:0] node24055;
	wire [4-1:0] node24060;
	wire [4-1:0] node24061;
	wire [4-1:0] node24062;
	wire [4-1:0] node24064;
	wire [4-1:0] node24068;
	wire [4-1:0] node24070;
	wire [4-1:0] node24073;
	wire [4-1:0] node24074;
	wire [4-1:0] node24075;
	wire [4-1:0] node24078;
	wire [4-1:0] node24080;
	wire [4-1:0] node24083;
	wire [4-1:0] node24084;
	wire [4-1:0] node24085;
	wire [4-1:0] node24086;
	wire [4-1:0] node24089;
	wire [4-1:0] node24094;
	wire [4-1:0] node24095;
	wire [4-1:0] node24096;
	wire [4-1:0] node24097;
	wire [4-1:0] node24099;
	wire [4-1:0] node24102;
	wire [4-1:0] node24103;
	wire [4-1:0] node24105;
	wire [4-1:0] node24108;
	wire [4-1:0] node24110;
	wire [4-1:0] node24113;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24118;
	wire [4-1:0] node24122;
	wire [4-1:0] node24123;
	wire [4-1:0] node24124;
	wire [4-1:0] node24125;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24131;
	wire [4-1:0] node24135;
	wire [4-1:0] node24138;
	wire [4-1:0] node24139;
	wire [4-1:0] node24140;
	wire [4-1:0] node24143;
	wire [4-1:0] node24147;
	wire [4-1:0] node24148;
	wire [4-1:0] node24149;
	wire [4-1:0] node24150;
	wire [4-1:0] node24151;
	wire [4-1:0] node24152;
	wire [4-1:0] node24153;
	wire [4-1:0] node24156;
	wire [4-1:0] node24160;
	wire [4-1:0] node24162;
	wire [4-1:0] node24165;
	wire [4-1:0] node24166;
	wire [4-1:0] node24167;
	wire [4-1:0] node24168;
	wire [4-1:0] node24173;
	wire [4-1:0] node24176;
	wire [4-1:0] node24177;
	wire [4-1:0] node24178;
	wire [4-1:0] node24179;
	wire [4-1:0] node24180;
	wire [4-1:0] node24183;
	wire [4-1:0] node24188;
	wire [4-1:0] node24189;
	wire [4-1:0] node24191;
	wire [4-1:0] node24195;
	wire [4-1:0] node24196;
	wire [4-1:0] node24197;
	wire [4-1:0] node24198;
	wire [4-1:0] node24201;
	wire [4-1:0] node24202;
	wire [4-1:0] node24203;
	wire [4-1:0] node24208;
	wire [4-1:0] node24210;
	wire [4-1:0] node24213;
	wire [4-1:0] node24214;
	wire [4-1:0] node24215;
	wire [4-1:0] node24217;
	wire [4-1:0] node24218;
	wire [4-1:0] node24221;
	wire [4-1:0] node24224;
	wire [4-1:0] node24226;
	wire [4-1:0] node24228;
	wire [4-1:0] node24231;
	wire [4-1:0] node24233;
	wire [4-1:0] node24236;
	wire [4-1:0] node24237;
	wire [4-1:0] node24238;
	wire [4-1:0] node24239;
	wire [4-1:0] node24240;
	wire [4-1:0] node24242;
	wire [4-1:0] node24244;
	wire [4-1:0] node24247;
	wire [4-1:0] node24249;
	wire [4-1:0] node24250;
	wire [4-1:0] node24253;
	wire [4-1:0] node24256;
	wire [4-1:0] node24257;
	wire [4-1:0] node24259;
	wire [4-1:0] node24260;
	wire [4-1:0] node24262;
	wire [4-1:0] node24265;
	wire [4-1:0] node24266;
	wire [4-1:0] node24270;
	wire [4-1:0] node24272;
	wire [4-1:0] node24274;
	wire [4-1:0] node24275;
	wire [4-1:0] node24278;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24283;
	wire [4-1:0] node24284;
	wire [4-1:0] node24285;
	wire [4-1:0] node24289;
	wire [4-1:0] node24290;
	wire [4-1:0] node24293;
	wire [4-1:0] node24296;
	wire [4-1:0] node24297;
	wire [4-1:0] node24298;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24306;
	wire [4-1:0] node24307;
	wire [4-1:0] node24312;
	wire [4-1:0] node24314;
	wire [4-1:0] node24317;
	wire [4-1:0] node24318;
	wire [4-1:0] node24319;
	wire [4-1:0] node24323;
	wire [4-1:0] node24324;
	wire [4-1:0] node24325;
	wire [4-1:0] node24328;
	wire [4-1:0] node24331;
	wire [4-1:0] node24332;
	wire [4-1:0] node24336;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24339;
	wire [4-1:0] node24340;
	wire [4-1:0] node24342;
	wire [4-1:0] node24346;
	wire [4-1:0] node24347;
	wire [4-1:0] node24350;
	wire [4-1:0] node24351;
	wire [4-1:0] node24355;
	wire [4-1:0] node24356;
	wire [4-1:0] node24357;
	wire [4-1:0] node24359;
	wire [4-1:0] node24360;
	wire [4-1:0] node24365;
	wire [4-1:0] node24366;
	wire [4-1:0] node24367;
	wire [4-1:0] node24369;
	wire [4-1:0] node24373;
	wire [4-1:0] node24375;
	wire [4-1:0] node24378;
	wire [4-1:0] node24379;
	wire [4-1:0] node24380;
	wire [4-1:0] node24381;
	wire [4-1:0] node24382;
	wire [4-1:0] node24383;
	wire [4-1:0] node24386;
	wire [4-1:0] node24389;
	wire [4-1:0] node24390;
	wire [4-1:0] node24394;
	wire [4-1:0] node24395;
	wire [4-1:0] node24397;
	wire [4-1:0] node24401;
	wire [4-1:0] node24403;
	wire [4-1:0] node24406;
	wire [4-1:0] node24407;
	wire [4-1:0] node24408;
	wire [4-1:0] node24411;
	wire [4-1:0] node24412;
	wire [4-1:0] node24415;
	wire [4-1:0] node24417;
	wire [4-1:0] node24420;
	wire [4-1:0] node24421;
	wire [4-1:0] node24422;
	wire [4-1:0] node24423;
	wire [4-1:0] node24426;
	wire [4-1:0] node24431;
	wire [4-1:0] node24432;
	wire [4-1:0] node24433;
	wire [4-1:0] node24434;
	wire [4-1:0] node24435;
	wire [4-1:0] node24437;
	wire [4-1:0] node24438;
	wire [4-1:0] node24440;
	wire [4-1:0] node24442;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24450;
	wire [4-1:0] node24451;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24458;
	wire [4-1:0] node24460;
	wire [4-1:0] node24463;
	wire [4-1:0] node24464;
	wire [4-1:0] node24465;
	wire [4-1:0] node24467;
	wire [4-1:0] node24470;
	wire [4-1:0] node24472;
	wire [4-1:0] node24475;
	wire [4-1:0] node24476;
	wire [4-1:0] node24478;
	wire [4-1:0] node24481;
	wire [4-1:0] node24483;
	wire [4-1:0] node24486;
	wire [4-1:0] node24487;
	wire [4-1:0] node24488;
	wire [4-1:0] node24489;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24493;
	wire [4-1:0] node24496;
	wire [4-1:0] node24498;
	wire [4-1:0] node24501;
	wire [4-1:0] node24502;
	wire [4-1:0] node24506;
	wire [4-1:0] node24508;
	wire [4-1:0] node24510;
	wire [4-1:0] node24512;
	wire [4-1:0] node24515;
	wire [4-1:0] node24516;
	wire [4-1:0] node24518;
	wire [4-1:0] node24521;
	wire [4-1:0] node24523;
	wire [4-1:0] node24525;
	wire [4-1:0] node24527;
	wire [4-1:0] node24530;
	wire [4-1:0] node24531;
	wire [4-1:0] node24532;
	wire [4-1:0] node24533;
	wire [4-1:0] node24534;
	wire [4-1:0] node24536;
	wire [4-1:0] node24541;
	wire [4-1:0] node24542;
	wire [4-1:0] node24545;
	wire [4-1:0] node24548;
	wire [4-1:0] node24549;
	wire [4-1:0] node24550;
	wire [4-1:0] node24552;
	wire [4-1:0] node24553;
	wire [4-1:0] node24558;
	wire [4-1:0] node24559;
	wire [4-1:0] node24562;
	wire [4-1:0] node24565;
	wire [4-1:0] node24566;
	wire [4-1:0] node24567;
	wire [4-1:0] node24568;
	wire [4-1:0] node24569;
	wire [4-1:0] node24570;
	wire [4-1:0] node24574;
	wire [4-1:0] node24576;
	wire [4-1:0] node24577;
	wire [4-1:0] node24581;
	wire [4-1:0] node24582;
	wire [4-1:0] node24583;
	wire [4-1:0] node24586;
	wire [4-1:0] node24589;
	wire [4-1:0] node24590;
	wire [4-1:0] node24591;
	wire [4-1:0] node24595;
	wire [4-1:0] node24596;
	wire [4-1:0] node24600;
	wire [4-1:0] node24601;
	wire [4-1:0] node24602;
	wire [4-1:0] node24603;
	wire [4-1:0] node24605;
	wire [4-1:0] node24609;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24613;
	wire [4-1:0] node24618;
	wire [4-1:0] node24619;
	wire [4-1:0] node24621;
	wire [4-1:0] node24622;
	wire [4-1:0] node24625;
	wire [4-1:0] node24628;
	wire [4-1:0] node24629;
	wire [4-1:0] node24630;
	wire [4-1:0] node24633;
	wire [4-1:0] node24636;
	wire [4-1:0] node24637;
	wire [4-1:0] node24641;
	wire [4-1:0] node24642;
	wire [4-1:0] node24643;
	wire [4-1:0] node24644;
	wire [4-1:0] node24645;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24653;
	wire [4-1:0] node24654;
	wire [4-1:0] node24655;
	wire [4-1:0] node24658;
	wire [4-1:0] node24661;
	wire [4-1:0] node24662;
	wire [4-1:0] node24665;
	wire [4-1:0] node24668;
	wire [4-1:0] node24669;
	wire [4-1:0] node24670;
	wire [4-1:0] node24674;
	wire [4-1:0] node24675;
	wire [4-1:0] node24676;
	wire [4-1:0] node24677;
	wire [4-1:0] node24680;
	wire [4-1:0] node24684;
	wire [4-1:0] node24685;
	wire [4-1:0] node24687;
	wire [4-1:0] node24690;
	wire [4-1:0] node24691;
	wire [4-1:0] node24695;
	wire [4-1:0] node24696;
	wire [4-1:0] node24697;
	wire [4-1:0] node24698;
	wire [4-1:0] node24699;
	wire [4-1:0] node24703;
	wire [4-1:0] node24704;
	wire [4-1:0] node24708;
	wire [4-1:0] node24710;
	wire [4-1:0] node24713;
	wire [4-1:0] node24714;
	wire [4-1:0] node24717;
	wire [4-1:0] node24720;
	wire [4-1:0] node24721;
	wire [4-1:0] node24722;
	wire [4-1:0] node24723;
	wire [4-1:0] node24724;
	wire [4-1:0] node24725;
	wire [4-1:0] node24726;
	wire [4-1:0] node24727;
	wire [4-1:0] node24729;
	wire [4-1:0] node24732;
	wire [4-1:0] node24735;
	wire [4-1:0] node24736;
	wire [4-1:0] node24739;
	wire [4-1:0] node24740;
	wire [4-1:0] node24744;
	wire [4-1:0] node24745;
	wire [4-1:0] node24747;
	wire [4-1:0] node24750;
	wire [4-1:0] node24751;
	wire [4-1:0] node24754;
	wire [4-1:0] node24757;
	wire [4-1:0] node24758;
	wire [4-1:0] node24759;
	wire [4-1:0] node24760;
	wire [4-1:0] node24761;
	wire [4-1:0] node24764;
	wire [4-1:0] node24767;
	wire [4-1:0] node24770;
	wire [4-1:0] node24771;
	wire [4-1:0] node24772;
	wire [4-1:0] node24773;
	wire [4-1:0] node24776;
	wire [4-1:0] node24781;
	wire [4-1:0] node24782;
	wire [4-1:0] node24784;
	wire [4-1:0] node24785;
	wire [4-1:0] node24789;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24795;
	wire [4-1:0] node24798;
	wire [4-1:0] node24799;
	wire [4-1:0] node24800;
	wire [4-1:0] node24801;
	wire [4-1:0] node24802;
	wire [4-1:0] node24804;
	wire [4-1:0] node24807;
	wire [4-1:0] node24808;
	wire [4-1:0] node24811;
	wire [4-1:0] node24814;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24817;
	wire [4-1:0] node24820;
	wire [4-1:0] node24823;
	wire [4-1:0] node24824;
	wire [4-1:0] node24827;
	wire [4-1:0] node24830;
	wire [4-1:0] node24831;
	wire [4-1:0] node24835;
	wire [4-1:0] node24836;
	wire [4-1:0] node24837;
	wire [4-1:0] node24838;
	wire [4-1:0] node24843;
	wire [4-1:0] node24844;
	wire [4-1:0] node24846;
	wire [4-1:0] node24849;
	wire [4-1:0] node24851;
	wire [4-1:0] node24852;
	wire [4-1:0] node24856;
	wire [4-1:0] node24857;
	wire [4-1:0] node24858;
	wire [4-1:0] node24859;
	wire [4-1:0] node24861;
	wire [4-1:0] node24864;
	wire [4-1:0] node24865;
	wire [4-1:0] node24869;
	wire [4-1:0] node24870;
	wire [4-1:0] node24871;
	wire [4-1:0] node24875;
	wire [4-1:0] node24876;
	wire [4-1:0] node24880;
	wire [4-1:0] node24881;
	wire [4-1:0] node24882;
	wire [4-1:0] node24885;
	wire [4-1:0] node24888;
	wire [4-1:0] node24889;
	wire [4-1:0] node24891;
	wire [4-1:0] node24894;
	wire [4-1:0] node24895;
	wire [4-1:0] node24899;
	wire [4-1:0] node24900;
	wire [4-1:0] node24901;
	wire [4-1:0] node24902;
	wire [4-1:0] node24903;
	wire [4-1:0] node24904;
	wire [4-1:0] node24905;
	wire [4-1:0] node24909;
	wire [4-1:0] node24910;
	wire [4-1:0] node24914;
	wire [4-1:0] node24917;
	wire [4-1:0] node24918;
	wire [4-1:0] node24919;
	wire [4-1:0] node24920;
	wire [4-1:0] node24924;
	wire [4-1:0] node24925;
	wire [4-1:0] node24928;
	wire [4-1:0] node24931;
	wire [4-1:0] node24932;
	wire [4-1:0] node24933;
	wire [4-1:0] node24937;
	wire [4-1:0] node24938;
	wire [4-1:0] node24942;
	wire [4-1:0] node24943;
	wire [4-1:0] node24944;
	wire [4-1:0] node24945;
	wire [4-1:0] node24947;
	wire [4-1:0] node24949;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24957;
	wire [4-1:0] node24958;
	wire [4-1:0] node24961;
	wire [4-1:0] node24962;
	wire [4-1:0] node24963;
	wire [4-1:0] node24967;
	wire [4-1:0] node24970;
	wire [4-1:0] node24972;
	wire [4-1:0] node24973;
	wire [4-1:0] node24974;
	wire [4-1:0] node24975;
	wire [4-1:0] node24980;
	wire [4-1:0] node24982;
	wire [4-1:0] node24984;
	wire [4-1:0] node24987;
	wire [4-1:0] node24988;
	wire [4-1:0] node24989;
	wire [4-1:0] node24990;
	wire [4-1:0] node24992;
	wire [4-1:0] node24993;
	wire [4-1:0] node24996;
	wire [4-1:0] node24999;
	wire [4-1:0] node25000;
	wire [4-1:0] node25002;
	wire [4-1:0] node25005;
	wire [4-1:0] node25006;
	wire [4-1:0] node25009;
	wire [4-1:0] node25012;
	wire [4-1:0] node25013;
	wire [4-1:0] node25015;
	wire [4-1:0] node25016;
	wire [4-1:0] node25020;
	wire [4-1:0] node25021;
	wire [4-1:0] node25024;
	wire [4-1:0] node25027;
	wire [4-1:0] node25028;
	wire [4-1:0] node25029;
	wire [4-1:0] node25030;
	wire [4-1:0] node25031;
	wire [4-1:0] node25036;
	wire [4-1:0] node25037;
	wire [4-1:0] node25038;
	wire [4-1:0] node25041;
	wire [4-1:0] node25045;
	wire [4-1:0] node25046;
	wire [4-1:0] node25047;
	wire [4-1:0] node25050;
	wire [4-1:0] node25053;
	wire [4-1:0] node25054;
	wire [4-1:0] node25056;
	wire [4-1:0] node25057;
	wire [4-1:0] node25061;
	wire [4-1:0] node25062;
	wire [4-1:0] node25065;
	wire [4-1:0] node25068;
	wire [4-1:0] node25069;
	wire [4-1:0] node25070;
	wire [4-1:0] node25071;
	wire [4-1:0] node25072;
	wire [4-1:0] node25073;
	wire [4-1:0] node25076;
	wire [4-1:0] node25077;
	wire [4-1:0] node25078;
	wire [4-1:0] node25080;
	wire [4-1:0] node25083;
	wire [4-1:0] node25085;
	wire [4-1:0] node25088;
	wire [4-1:0] node25091;
	wire [4-1:0] node25092;
	wire [4-1:0] node25093;
	wire [4-1:0] node25096;
	wire [4-1:0] node25099;
	wire [4-1:0] node25100;
	wire [4-1:0] node25104;
	wire [4-1:0] node25105;
	wire [4-1:0] node25106;
	wire [4-1:0] node25108;
	wire [4-1:0] node25110;
	wire [4-1:0] node25113;
	wire [4-1:0] node25115;
	wire [4-1:0] node25117;
	wire [4-1:0] node25120;
	wire [4-1:0] node25121;
	wire [4-1:0] node25123;
	wire [4-1:0] node25124;
	wire [4-1:0] node25127;
	wire [4-1:0] node25130;
	wire [4-1:0] node25131;
	wire [4-1:0] node25132;
	wire [4-1:0] node25133;
	wire [4-1:0] node25136;
	wire [4-1:0] node25141;
	wire [4-1:0] node25142;
	wire [4-1:0] node25143;
	wire [4-1:0] node25144;
	wire [4-1:0] node25145;
	wire [4-1:0] node25146;
	wire [4-1:0] node25148;
	wire [4-1:0] node25153;
	wire [4-1:0] node25154;
	wire [4-1:0] node25155;
	wire [4-1:0] node25159;
	wire [4-1:0] node25160;
	wire [4-1:0] node25163;
	wire [4-1:0] node25165;
	wire [4-1:0] node25168;
	wire [4-1:0] node25169;
	wire [4-1:0] node25170;
	wire [4-1:0] node25171;
	wire [4-1:0] node25174;
	wire [4-1:0] node25177;
	wire [4-1:0] node25178;
	wire [4-1:0] node25182;
	wire [4-1:0] node25183;
	wire [4-1:0] node25186;
	wire [4-1:0] node25189;
	wire [4-1:0] node25190;
	wire [4-1:0] node25191;
	wire [4-1:0] node25192;
	wire [4-1:0] node25195;
	wire [4-1:0] node25196;
	wire [4-1:0] node25199;
	wire [4-1:0] node25200;
	wire [4-1:0] node25204;
	wire [4-1:0] node25205;
	wire [4-1:0] node25206;
	wire [4-1:0] node25209;
	wire [4-1:0] node25212;
	wire [4-1:0] node25213;
	wire [4-1:0] node25216;
	wire [4-1:0] node25219;
	wire [4-1:0] node25220;
	wire [4-1:0] node25221;
	wire [4-1:0] node25222;
	wire [4-1:0] node25227;
	wire [4-1:0] node25228;
	wire [4-1:0] node25232;
	wire [4-1:0] node25233;
	wire [4-1:0] node25234;
	wire [4-1:0] node25235;
	wire [4-1:0] node25236;
	wire [4-1:0] node25237;
	wire [4-1:0] node25238;
	wire [4-1:0] node25239;
	wire [4-1:0] node25243;
	wire [4-1:0] node25247;
	wire [4-1:0] node25248;
	wire [4-1:0] node25252;
	wire [4-1:0] node25253;
	wire [4-1:0] node25254;
	wire [4-1:0] node25256;
	wire [4-1:0] node25260;
	wire [4-1:0] node25263;
	wire [4-1:0] node25264;
	wire [4-1:0] node25265;
	wire [4-1:0] node25266;
	wire [4-1:0] node25268;
	wire [4-1:0] node25272;
	wire [4-1:0] node25273;
	wire [4-1:0] node25277;
	wire [4-1:0] node25278;
	wire [4-1:0] node25279;
	wire [4-1:0] node25281;
	wire [4-1:0] node25285;
	wire [4-1:0] node25286;
	wire [4-1:0] node25290;
	wire [4-1:0] node25291;
	wire [4-1:0] node25292;
	wire [4-1:0] node25293;
	wire [4-1:0] node25295;
	wire [4-1:0] node25297;
	wire [4-1:0] node25299;
	wire [4-1:0] node25303;
	wire [4-1:0] node25304;
	wire [4-1:0] node25308;
	wire [4-1:0] node25309;
	wire [4-1:0] node25310;
	wire [4-1:0] node25311;
	wire [4-1:0] node25312;
	wire [4-1:0] node25314;
	wire [4-1:0] node25320;
	wire [4-1:0] node25321;
	wire [4-1:0] node25325;
	wire [4-1:0] node25326;
	wire [4-1:0] node25327;
	wire [4-1:0] node25328;
	wire [4-1:0] node25329;
	wire [4-1:0] node25330;
	wire [4-1:0] node25331;
	wire [4-1:0] node25332;
	wire [4-1:0] node25333;
	wire [4-1:0] node25334;
	wire [4-1:0] node25335;
	wire [4-1:0] node25336;
	wire [4-1:0] node25340;
	wire [4-1:0] node25343;
	wire [4-1:0] node25345;
	wire [4-1:0] node25348;
	wire [4-1:0] node25349;
	wire [4-1:0] node25350;
	wire [4-1:0] node25351;
	wire [4-1:0] node25354;
	wire [4-1:0] node25356;
	wire [4-1:0] node25359;
	wire [4-1:0] node25361;
	wire [4-1:0] node25364;
	wire [4-1:0] node25365;
	wire [4-1:0] node25367;
	wire [4-1:0] node25370;
	wire [4-1:0] node25373;
	wire [4-1:0] node25374;
	wire [4-1:0] node25375;
	wire [4-1:0] node25376;
	wire [4-1:0] node25377;
	wire [4-1:0] node25378;
	wire [4-1:0] node25382;
	wire [4-1:0] node25385;
	wire [4-1:0] node25386;
	wire [4-1:0] node25389;
	wire [4-1:0] node25391;
	wire [4-1:0] node25394;
	wire [4-1:0] node25395;
	wire [4-1:0] node25396;
	wire [4-1:0] node25399;
	wire [4-1:0] node25400;
	wire [4-1:0] node25403;
	wire [4-1:0] node25406;
	wire [4-1:0] node25407;
	wire [4-1:0] node25411;
	wire [4-1:0] node25412;
	wire [4-1:0] node25413;
	wire [4-1:0] node25415;
	wire [4-1:0] node25419;
	wire [4-1:0] node25420;
	wire [4-1:0] node25424;
	wire [4-1:0] node25425;
	wire [4-1:0] node25426;
	wire [4-1:0] node25427;
	wire [4-1:0] node25428;
	wire [4-1:0] node25429;
	wire [4-1:0] node25432;
	wire [4-1:0] node25436;
	wire [4-1:0] node25437;
	wire [4-1:0] node25439;
	wire [4-1:0] node25440;
	wire [4-1:0] node25443;
	wire [4-1:0] node25446;
	wire [4-1:0] node25447;
	wire [4-1:0] node25449;
	wire [4-1:0] node25452;
	wire [4-1:0] node25455;
	wire [4-1:0] node25456;
	wire [4-1:0] node25458;
	wire [4-1:0] node25459;
	wire [4-1:0] node25462;
	wire [4-1:0] node25465;
	wire [4-1:0] node25466;
	wire [4-1:0] node25468;
	wire [4-1:0] node25471;
	wire [4-1:0] node25473;
	wire [4-1:0] node25475;
	wire [4-1:0] node25478;
	wire [4-1:0] node25479;
	wire [4-1:0] node25480;
	wire [4-1:0] node25481;
	wire [4-1:0] node25482;
	wire [4-1:0] node25483;
	wire [4-1:0] node25486;
	wire [4-1:0] node25491;
	wire [4-1:0] node25493;
	wire [4-1:0] node25495;
	wire [4-1:0] node25498;
	wire [4-1:0] node25499;
	wire [4-1:0] node25500;
	wire [4-1:0] node25503;
	wire [4-1:0] node25504;
	wire [4-1:0] node25505;
	wire [4-1:0] node25508;
	wire [4-1:0] node25512;
	wire [4-1:0] node25513;
	wire [4-1:0] node25514;
	wire [4-1:0] node25515;
	wire [4-1:0] node25519;
	wire [4-1:0] node25520;
	wire [4-1:0] node25523;
	wire [4-1:0] node25526;
	wire [4-1:0] node25529;
	wire [4-1:0] node25530;
	wire [4-1:0] node25531;
	wire [4-1:0] node25532;
	wire [4-1:0] node25533;
	wire [4-1:0] node25534;
	wire [4-1:0] node25536;
	wire [4-1:0] node25539;
	wire [4-1:0] node25540;
	wire [4-1:0] node25543;
	wire [4-1:0] node25546;
	wire [4-1:0] node25547;
	wire [4-1:0] node25549;
	wire [4-1:0] node25552;
	wire [4-1:0] node25553;
	wire [4-1:0] node25556;
	wire [4-1:0] node25559;
	wire [4-1:0] node25560;
	wire [4-1:0] node25562;
	wire [4-1:0] node25563;
	wire [4-1:0] node25566;
	wire [4-1:0] node25568;
	wire [4-1:0] node25571;
	wire [4-1:0] node25572;
	wire [4-1:0] node25573;
	wire [4-1:0] node25576;
	wire [4-1:0] node25577;
	wire [4-1:0] node25581;
	wire [4-1:0] node25584;
	wire [4-1:0] node25585;
	wire [4-1:0] node25586;
	wire [4-1:0] node25587;
	wire [4-1:0] node25589;
	wire [4-1:0] node25592;
	wire [4-1:0] node25593;
	wire [4-1:0] node25597;
	wire [4-1:0] node25599;
	wire [4-1:0] node25600;
	wire [4-1:0] node25604;
	wire [4-1:0] node25605;
	wire [4-1:0] node25606;
	wire [4-1:0] node25607;
	wire [4-1:0] node25611;
	wire [4-1:0] node25612;
	wire [4-1:0] node25616;
	wire [4-1:0] node25617;
	wire [4-1:0] node25618;
	wire [4-1:0] node25621;
	wire [4-1:0] node25622;
	wire [4-1:0] node25626;
	wire [4-1:0] node25627;
	wire [4-1:0] node25631;
	wire [4-1:0] node25632;
	wire [4-1:0] node25633;
	wire [4-1:0] node25634;
	wire [4-1:0] node25635;
	wire [4-1:0] node25637;
	wire [4-1:0] node25638;
	wire [4-1:0] node25641;
	wire [4-1:0] node25645;
	wire [4-1:0] node25647;
	wire [4-1:0] node25650;
	wire [4-1:0] node25651;
	wire [4-1:0] node25652;
	wire [4-1:0] node25656;
	wire [4-1:0] node25658;
	wire [4-1:0] node25659;
	wire [4-1:0] node25661;
	wire [4-1:0] node25664;
	wire [4-1:0] node25666;
	wire [4-1:0] node25669;
	wire [4-1:0] node25670;
	wire [4-1:0] node25671;
	wire [4-1:0] node25672;
	wire [4-1:0] node25674;
	wire [4-1:0] node25678;
	wire [4-1:0] node25680;
	wire [4-1:0] node25681;
	wire [4-1:0] node25685;
	wire [4-1:0] node25686;
	wire [4-1:0] node25688;
	wire [4-1:0] node25689;
	wire [4-1:0] node25692;
	wire [4-1:0] node25694;
	wire [4-1:0] node25697;
	wire [4-1:0] node25699;
	wire [4-1:0] node25702;
	wire [4-1:0] node25703;
	wire [4-1:0] node25704;
	wire [4-1:0] node25705;
	wire [4-1:0] node25706;
	wire [4-1:0] node25707;
	wire [4-1:0] node25708;
	wire [4-1:0] node25709;
	wire [4-1:0] node25712;
	wire [4-1:0] node25715;
	wire [4-1:0] node25718;
	wire [4-1:0] node25719;
	wire [4-1:0] node25721;
	wire [4-1:0] node25724;
	wire [4-1:0] node25725;
	wire [4-1:0] node25729;
	wire [4-1:0] node25730;
	wire [4-1:0] node25731;
	wire [4-1:0] node25732;
	wire [4-1:0] node25736;
	wire [4-1:0] node25737;
	wire [4-1:0] node25741;
	wire [4-1:0] node25744;
	wire [4-1:0] node25745;
	wire [4-1:0] node25746;
	wire [4-1:0] node25747;
	wire [4-1:0] node25748;
	wire [4-1:0] node25750;
	wire [4-1:0] node25753;
	wire [4-1:0] node25756;
	wire [4-1:0] node25758;
	wire [4-1:0] node25761;
	wire [4-1:0] node25762;
	wire [4-1:0] node25764;
	wire [4-1:0] node25768;
	wire [4-1:0] node25769;
	wire [4-1:0] node25770;
	wire [4-1:0] node25771;
	wire [4-1:0] node25775;
	wire [4-1:0] node25776;
	wire [4-1:0] node25777;
	wire [4-1:0] node25780;
	wire [4-1:0] node25783;
	wire [4-1:0] node25785;
	wire [4-1:0] node25788;
	wire [4-1:0] node25789;
	wire [4-1:0] node25791;
	wire [4-1:0] node25792;
	wire [4-1:0] node25796;
	wire [4-1:0] node25797;
	wire [4-1:0] node25800;
	wire [4-1:0] node25803;
	wire [4-1:0] node25804;
	wire [4-1:0] node25805;
	wire [4-1:0] node25806;
	wire [4-1:0] node25807;
	wire [4-1:0] node25809;
	wire [4-1:0] node25811;
	wire [4-1:0] node25814;
	wire [4-1:0] node25815;
	wire [4-1:0] node25818;
	wire [4-1:0] node25819;
	wire [4-1:0] node25823;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25830;
	wire [4-1:0] node25833;
	wire [4-1:0] node25835;
	wire [4-1:0] node25838;
	wire [4-1:0] node25839;
	wire [4-1:0] node25840;
	wire [4-1:0] node25842;
	wire [4-1:0] node25843;
	wire [4-1:0] node25847;
	wire [4-1:0] node25849;
	wire [4-1:0] node25852;
	wire [4-1:0] node25853;
	wire [4-1:0] node25854;
	wire [4-1:0] node25855;
	wire [4-1:0] node25860;
	wire [4-1:0] node25861;
	wire [4-1:0] node25864;
	wire [4-1:0] node25866;
	wire [4-1:0] node25869;
	wire [4-1:0] node25870;
	wire [4-1:0] node25871;
	wire [4-1:0] node25872;
	wire [4-1:0] node25875;
	wire [4-1:0] node25876;
	wire [4-1:0] node25880;
	wire [4-1:0] node25882;
	wire [4-1:0] node25883;
	wire [4-1:0] node25887;
	wire [4-1:0] node25888;
	wire [4-1:0] node25890;
	wire [4-1:0] node25893;
	wire [4-1:0] node25894;
	wire [4-1:0] node25895;
	wire [4-1:0] node25898;
	wire [4-1:0] node25901;
	wire [4-1:0] node25902;
	wire [4-1:0] node25905;
	wire [4-1:0] node25906;
	wire [4-1:0] node25909;
	wire [4-1:0] node25912;
	wire [4-1:0] node25913;
	wire [4-1:0] node25914;
	wire [4-1:0] node25915;
	wire [4-1:0] node25916;
	wire [4-1:0] node25917;
	wire [4-1:0] node25918;
	wire [4-1:0] node25921;
	wire [4-1:0] node25925;
	wire [4-1:0] node25926;
	wire [4-1:0] node25927;
	wire [4-1:0] node25931;
	wire [4-1:0] node25932;
	wire [4-1:0] node25936;
	wire [4-1:0] node25937;
	wire [4-1:0] node25938;
	wire [4-1:0] node25940;
	wire [4-1:0] node25943;
	wire [4-1:0] node25944;
	wire [4-1:0] node25945;
	wire [4-1:0] node25949;
	wire [4-1:0] node25951;
	wire [4-1:0] node25955;
	wire [4-1:0] node25956;
	wire [4-1:0] node25957;
	wire [4-1:0] node25959;
	wire [4-1:0] node25960;
	wire [4-1:0] node25963;
	wire [4-1:0] node25966;
	wire [4-1:0] node25967;
	wire [4-1:0] node25968;
	wire [4-1:0] node25972;
	wire [4-1:0] node25973;
	wire [4-1:0] node25977;
	wire [4-1:0] node25978;
	wire [4-1:0] node25979;
	wire [4-1:0] node25980;
	wire [4-1:0] node25983;
	wire [4-1:0] node25986;
	wire [4-1:0] node25987;
	wire [4-1:0] node25990;
	wire [4-1:0] node25993;
	wire [4-1:0] node25994;
	wire [4-1:0] node25995;
	wire [4-1:0] node25996;
	wire [4-1:0] node26000;
	wire [4-1:0] node26002;
	wire [4-1:0] node26005;
	wire [4-1:0] node26006;
	wire [4-1:0] node26009;
	wire [4-1:0] node26012;
	wire [4-1:0] node26013;
	wire [4-1:0] node26014;
	wire [4-1:0] node26015;
	wire [4-1:0] node26016;
	wire [4-1:0] node26017;
	wire [4-1:0] node26021;
	wire [4-1:0] node26022;
	wire [4-1:0] node26025;
	wire [4-1:0] node26026;
	wire [4-1:0] node26030;
	wire [4-1:0] node26031;
	wire [4-1:0] node26032;
	wire [4-1:0] node26033;
	wire [4-1:0] node26036;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26044;
	wire [4-1:0] node26047;
	wire [4-1:0] node26048;
	wire [4-1:0] node26051;
	wire [4-1:0] node26052;
	wire [4-1:0] node26054;
	wire [4-1:0] node26055;
	wire [4-1:0] node26058;
	wire [4-1:0] node26061;
	wire [4-1:0] node26062;
	wire [4-1:0] node26064;
	wire [4-1:0] node26067;
	wire [4-1:0] node26070;
	wire [4-1:0] node26071;
	wire [4-1:0] node26072;
	wire [4-1:0] node26074;
	wire [4-1:0] node26077;
	wire [4-1:0] node26078;
	wire [4-1:0] node26079;
	wire [4-1:0] node26081;
	wire [4-1:0] node26085;
	wire [4-1:0] node26088;
	wire [4-1:0] node26089;
	wire [4-1:0] node26091;
	wire [4-1:0] node26093;
	wire [4-1:0] node26094;
	wire [4-1:0] node26098;
	wire [4-1:0] node26099;
	wire [4-1:0] node26101;
	wire [4-1:0] node26103;
	wire [4-1:0] node26106;
	wire [4-1:0] node26108;
	wire [4-1:0] node26111;
	wire [4-1:0] node26112;
	wire [4-1:0] node26113;
	wire [4-1:0] node26114;
	wire [4-1:0] node26115;
	wire [4-1:0] node26116;
	wire [4-1:0] node26117;
	wire [4-1:0] node26118;
	wire [4-1:0] node26119;
	wire [4-1:0] node26124;
	wire [4-1:0] node26125;
	wire [4-1:0] node26126;
	wire [4-1:0] node26127;
	wire [4-1:0] node26132;
	wire [4-1:0] node26135;
	wire [4-1:0] node26136;
	wire [4-1:0] node26137;
	wire [4-1:0] node26138;
	wire [4-1:0] node26141;
	wire [4-1:0] node26142;
	wire [4-1:0] node26146;
	wire [4-1:0] node26147;
	wire [4-1:0] node26149;
	wire [4-1:0] node26152;
	wire [4-1:0] node26155;
	wire [4-1:0] node26156;
	wire [4-1:0] node26157;
	wire [4-1:0] node26160;
	wire [4-1:0] node26162;
	wire [4-1:0] node26165;
	wire [4-1:0] node26166;
	wire [4-1:0] node26170;
	wire [4-1:0] node26171;
	wire [4-1:0] node26172;
	wire [4-1:0] node26174;
	wire [4-1:0] node26176;
	wire [4-1:0] node26179;
	wire [4-1:0] node26180;
	wire [4-1:0] node26181;
	wire [4-1:0] node26182;
	wire [4-1:0] node26185;
	wire [4-1:0] node26189;
	wire [4-1:0] node26190;
	wire [4-1:0] node26194;
	wire [4-1:0] node26195;
	wire [4-1:0] node26196;
	wire [4-1:0] node26198;
	wire [4-1:0] node26201;
	wire [4-1:0] node26202;
	wire [4-1:0] node26203;
	wire [4-1:0] node26206;
	wire [4-1:0] node26209;
	wire [4-1:0] node26210;
	wire [4-1:0] node26214;
	wire [4-1:0] node26215;
	wire [4-1:0] node26217;
	wire [4-1:0] node26220;
	wire [4-1:0] node26221;
	wire [4-1:0] node26223;
	wire [4-1:0] node26226;
	wire [4-1:0] node26229;
	wire [4-1:0] node26230;
	wire [4-1:0] node26231;
	wire [4-1:0] node26232;
	wire [4-1:0] node26233;
	wire [4-1:0] node26237;
	wire [4-1:0] node26238;
	wire [4-1:0] node26240;
	wire [4-1:0] node26243;
	wire [4-1:0] node26244;
	wire [4-1:0] node26247;
	wire [4-1:0] node26250;
	wire [4-1:0] node26251;
	wire [4-1:0] node26252;
	wire [4-1:0] node26254;
	wire [4-1:0] node26257;
	wire [4-1:0] node26259;
	wire [4-1:0] node26260;
	wire [4-1:0] node26263;
	wire [4-1:0] node26266;
	wire [4-1:0] node26267;
	wire [4-1:0] node26268;
	wire [4-1:0] node26272;
	wire [4-1:0] node26275;
	wire [4-1:0] node26276;
	wire [4-1:0] node26277;
	wire [4-1:0] node26278;
	wire [4-1:0] node26281;
	wire [4-1:0] node26282;
	wire [4-1:0] node26286;
	wire [4-1:0] node26289;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26292;
	wire [4-1:0] node26296;
	wire [4-1:0] node26297;
	wire [4-1:0] node26300;
	wire [4-1:0] node26302;
	wire [4-1:0] node26305;
	wire [4-1:0] node26306;
	wire [4-1:0] node26307;
	wire [4-1:0] node26308;
	wire [4-1:0] node26311;
	wire [4-1:0] node26314;
	wire [4-1:0] node26317;
	wire [4-1:0] node26319;
	wire [4-1:0] node26321;
	wire [4-1:0] node26324;
	wire [4-1:0] node26325;
	wire [4-1:0] node26326;
	wire [4-1:0] node26327;
	wire [4-1:0] node26328;
	wire [4-1:0] node26329;
	wire [4-1:0] node26330;
	wire [4-1:0] node26332;
	wire [4-1:0] node26335;
	wire [4-1:0] node26337;
	wire [4-1:0] node26341;
	wire [4-1:0] node26342;
	wire [4-1:0] node26343;
	wire [4-1:0] node26347;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26352;
	wire [4-1:0] node26353;
	wire [4-1:0] node26357;
	wire [4-1:0] node26358;
	wire [4-1:0] node26361;
	wire [4-1:0] node26364;
	wire [4-1:0] node26365;
	wire [4-1:0] node26367;
	wire [4-1:0] node26370;
	wire [4-1:0] node26372;
	wire [4-1:0] node26375;
	wire [4-1:0] node26376;
	wire [4-1:0] node26377;
	wire [4-1:0] node26378;
	wire [4-1:0] node26381;
	wire [4-1:0] node26383;
	wire [4-1:0] node26386;
	wire [4-1:0] node26387;
	wire [4-1:0] node26388;
	wire [4-1:0] node26390;
	wire [4-1:0] node26393;
	wire [4-1:0] node26397;
	wire [4-1:0] node26398;
	wire [4-1:0] node26399;
	wire [4-1:0] node26400;
	wire [4-1:0] node26401;
	wire [4-1:0] node26405;
	wire [4-1:0] node26406;
	wire [4-1:0] node26410;
	wire [4-1:0] node26413;
	wire [4-1:0] node26414;
	wire [4-1:0] node26417;
	wire [4-1:0] node26419;
	wire [4-1:0] node26422;
	wire [4-1:0] node26423;
	wire [4-1:0] node26424;
	wire [4-1:0] node26425;
	wire [4-1:0] node26426;
	wire [4-1:0] node26429;
	wire [4-1:0] node26432;
	wire [4-1:0] node26433;
	wire [4-1:0] node26434;
	wire [4-1:0] node26435;
	wire [4-1:0] node26441;
	wire [4-1:0] node26442;
	wire [4-1:0] node26443;
	wire [4-1:0] node26445;
	wire [4-1:0] node26446;
	wire [4-1:0] node26450;
	wire [4-1:0] node26452;
	wire [4-1:0] node26455;
	wire [4-1:0] node26457;
	wire [4-1:0] node26459;
	wire [4-1:0] node26461;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26466;
	wire [4-1:0] node26467;
	wire [4-1:0] node26471;
	wire [4-1:0] node26472;
	wire [4-1:0] node26475;
	wire [4-1:0] node26476;
	wire [4-1:0] node26479;
	wire [4-1:0] node26482;
	wire [4-1:0] node26483;
	wire [4-1:0] node26484;
	wire [4-1:0] node26487;
	wire [4-1:0] node26488;
	wire [4-1:0] node26492;
	wire [4-1:0] node26493;
	wire [4-1:0] node26496;
	wire [4-1:0] node26498;
	wire [4-1:0] node26501;
	wire [4-1:0] node26502;
	wire [4-1:0] node26503;
	wire [4-1:0] node26504;
	wire [4-1:0] node26505;
	wire [4-1:0] node26506;
	wire [4-1:0] node26507;
	wire [4-1:0] node26509;
	wire [4-1:0] node26511;
	wire [4-1:0] node26514;
	wire [4-1:0] node26516;
	wire [4-1:0] node26519;
	wire [4-1:0] node26520;
	wire [4-1:0] node26522;
	wire [4-1:0] node26526;
	wire [4-1:0] node26527;
	wire [4-1:0] node26528;
	wire [4-1:0] node26530;
	wire [4-1:0] node26533;
	wire [4-1:0] node26534;
	wire [4-1:0] node26537;
	wire [4-1:0] node26540;
	wire [4-1:0] node26541;
	wire [4-1:0] node26543;
	wire [4-1:0] node26544;
	wire [4-1:0] node26547;
	wire [4-1:0] node26551;
	wire [4-1:0] node26552;
	wire [4-1:0] node26553;
	wire [4-1:0] node26554;
	wire [4-1:0] node26555;
	wire [4-1:0] node26557;
	wire [4-1:0] node26560;
	wire [4-1:0] node26563;
	wire [4-1:0] node26565;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26571;
	wire [4-1:0] node26572;
	wire [4-1:0] node26576;
	wire [4-1:0] node26578;
	wire [4-1:0] node26580;
	wire [4-1:0] node26583;
	wire [4-1:0] node26584;
	wire [4-1:0] node26585;
	wire [4-1:0] node26587;
	wire [4-1:0] node26589;
	wire [4-1:0] node26592;
	wire [4-1:0] node26593;
	wire [4-1:0] node26597;
	wire [4-1:0] node26598;
	wire [4-1:0] node26601;
	wire [4-1:0] node26604;
	wire [4-1:0] node26605;
	wire [4-1:0] node26606;
	wire [4-1:0] node26607;
	wire [4-1:0] node26608;
	wire [4-1:0] node26610;
	wire [4-1:0] node26612;
	wire [4-1:0] node26615;
	wire [4-1:0] node26616;
	wire [4-1:0] node26617;
	wire [4-1:0] node26620;
	wire [4-1:0] node26624;
	wire [4-1:0] node26625;
	wire [4-1:0] node26627;
	wire [4-1:0] node26630;
	wire [4-1:0] node26631;
	wire [4-1:0] node26632;
	wire [4-1:0] node26636;
	wire [4-1:0] node26639;
	wire [4-1:0] node26640;
	wire [4-1:0] node26642;
	wire [4-1:0] node26643;
	wire [4-1:0] node26646;
	wire [4-1:0] node26648;
	wire [4-1:0] node26651;
	wire [4-1:0] node26652;
	wire [4-1:0] node26653;
	wire [4-1:0] node26657;
	wire [4-1:0] node26658;
	wire [4-1:0] node26661;
	wire [4-1:0] node26664;
	wire [4-1:0] node26665;
	wire [4-1:0] node26666;
	wire [4-1:0] node26667;
	wire [4-1:0] node26668;
	wire [4-1:0] node26671;
	wire [4-1:0] node26675;
	wire [4-1:0] node26676;
	wire [4-1:0] node26679;
	wire [4-1:0] node26680;
	wire [4-1:0] node26681;
	wire [4-1:0] node26685;
	wire [4-1:0] node26687;
	wire [4-1:0] node26690;
	wire [4-1:0] node26691;
	wire [4-1:0] node26692;
	wire [4-1:0] node26693;
	wire [4-1:0] node26694;
	wire [4-1:0] node26698;
	wire [4-1:0] node26701;
	wire [4-1:0] node26702;
	wire [4-1:0] node26705;
	wire [4-1:0] node26707;
	wire [4-1:0] node26710;
	wire [4-1:0] node26711;
	wire [4-1:0] node26714;
	wire [4-1:0] node26717;
	wire [4-1:0] node26718;
	wire [4-1:0] node26719;
	wire [4-1:0] node26720;
	wire [4-1:0] node26721;
	wire [4-1:0] node26722;
	wire [4-1:0] node26723;
	wire [4-1:0] node26726;
	wire [4-1:0] node26729;
	wire [4-1:0] node26730;
	wire [4-1:0] node26734;
	wire [4-1:0] node26735;
	wire [4-1:0] node26736;
	wire [4-1:0] node26738;
	wire [4-1:0] node26741;
	wire [4-1:0] node26742;
	wire [4-1:0] node26746;
	wire [4-1:0] node26747;
	wire [4-1:0] node26750;
	wire [4-1:0] node26753;
	wire [4-1:0] node26754;
	wire [4-1:0] node26755;
	wire [4-1:0] node26759;
	wire [4-1:0] node26760;
	wire [4-1:0] node26762;
	wire [4-1:0] node26764;
	wire [4-1:0] node26767;
	wire [4-1:0] node26768;
	wire [4-1:0] node26771;
	wire [4-1:0] node26774;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26777;
	wire [4-1:0] node26778;
	wire [4-1:0] node26781;
	wire [4-1:0] node26784;
	wire [4-1:0] node26785;
	wire [4-1:0] node26788;
	wire [4-1:0] node26791;
	wire [4-1:0] node26793;
	wire [4-1:0] node26794;
	wire [4-1:0] node26797;
	wire [4-1:0] node26800;
	wire [4-1:0] node26801;
	wire [4-1:0] node26802;
	wire [4-1:0] node26804;
	wire [4-1:0] node26808;
	wire [4-1:0] node26809;
	wire [4-1:0] node26810;
	wire [4-1:0] node26813;
	wire [4-1:0] node26815;
	wire [4-1:0] node26818;
	wire [4-1:0] node26820;
	wire [4-1:0] node26823;
	wire [4-1:0] node26824;
	wire [4-1:0] node26825;
	wire [4-1:0] node26826;
	wire [4-1:0] node26827;
	wire [4-1:0] node26829;
	wire [4-1:0] node26830;
	wire [4-1:0] node26834;
	wire [4-1:0] node26835;
	wire [4-1:0] node26838;
	wire [4-1:0] node26840;
	wire [4-1:0] node26843;
	wire [4-1:0] node26844;
	wire [4-1:0] node26845;
	wire [4-1:0] node26846;
	wire [4-1:0] node26851;
	wire [4-1:0] node26854;
	wire [4-1:0] node26855;
	wire [4-1:0] node26856;
	wire [4-1:0] node26857;
	wire [4-1:0] node26860;
	wire [4-1:0] node26861;
	wire [4-1:0] node26865;
	wire [4-1:0] node26866;
	wire [4-1:0] node26867;
	wire [4-1:0] node26872;
	wire [4-1:0] node26873;
	wire [4-1:0] node26874;
	wire [4-1:0] node26878;
	wire [4-1:0] node26880;
	wire [4-1:0] node26883;
	wire [4-1:0] node26884;
	wire [4-1:0] node26885;
	wire [4-1:0] node26886;
	wire [4-1:0] node26887;
	wire [4-1:0] node26890;
	wire [4-1:0] node26892;
	wire [4-1:0] node26895;
	wire [4-1:0] node26896;
	wire [4-1:0] node26897;
	wire [4-1:0] node26902;
	wire [4-1:0] node26903;
	wire [4-1:0] node26904;
	wire [4-1:0] node26905;
	wire [4-1:0] node26909;
	wire [4-1:0] node26911;
	wire [4-1:0] node26914;
	wire [4-1:0] node26917;
	wire [4-1:0] node26918;
	wire [4-1:0] node26920;
	wire [4-1:0] node26921;
	wire [4-1:0] node26925;
	wire [4-1:0] node26926;
	wire [4-1:0] node26927;
	wire [4-1:0] node26929;
	wire [4-1:0] node26932;
	wire [4-1:0] node26935;
	wire [4-1:0] node26938;
	wire [4-1:0] node26939;
	wire [4-1:0] node26940;
	wire [4-1:0] node26941;
	wire [4-1:0] node26942;
	wire [4-1:0] node26943;
	wire [4-1:0] node26944;
	wire [4-1:0] node26945;
	wire [4-1:0] node26946;
	wire [4-1:0] node26950;
	wire [4-1:0] node26951;
	wire [4-1:0] node26954;
	wire [4-1:0] node26957;
	wire [4-1:0] node26958;
	wire [4-1:0] node26961;
	wire [4-1:0] node26962;
	wire [4-1:0] node26965;
	wire [4-1:0] node26968;
	wire [4-1:0] node26969;
	wire [4-1:0] node26970;
	wire [4-1:0] node26973;
	wire [4-1:0] node26974;
	wire [4-1:0] node26977;
	wire [4-1:0] node26980;
	wire [4-1:0] node26981;
	wire [4-1:0] node26984;
	wire [4-1:0] node26985;
	wire [4-1:0] node26988;
	wire [4-1:0] node26991;
	wire [4-1:0] node26992;
	wire [4-1:0] node26993;
	wire [4-1:0] node26994;
	wire [4-1:0] node26995;
	wire [4-1:0] node26996;
	wire [4-1:0] node26999;
	wire [4-1:0] node27003;
	wire [4-1:0] node27004;
	wire [4-1:0] node27007;
	wire [4-1:0] node27008;
	wire [4-1:0] node27012;
	wire [4-1:0] node27013;
	wire [4-1:0] node27014;
	wire [4-1:0] node27015;
	wire [4-1:0] node27016;
	wire [4-1:0] node27019;
	wire [4-1:0] node27024;
	wire [4-1:0] node27025;
	wire [4-1:0] node27028;
	wire [4-1:0] node27029;
	wire [4-1:0] node27033;
	wire [4-1:0] node27034;
	wire [4-1:0] node27035;
	wire [4-1:0] node27036;
	wire [4-1:0] node27037;
	wire [4-1:0] node27041;
	wire [4-1:0] node27042;
	wire [4-1:0] node27046;
	wire [4-1:0] node27047;
	wire [4-1:0] node27048;
	wire [4-1:0] node27052;
	wire [4-1:0] node27053;
	wire [4-1:0] node27056;
	wire [4-1:0] node27059;
	wire [4-1:0] node27060;
	wire [4-1:0] node27061;
	wire [4-1:0] node27063;
	wire [4-1:0] node27066;
	wire [4-1:0] node27067;
	wire [4-1:0] node27070;
	wire [4-1:0] node27073;
	wire [4-1:0] node27074;
	wire [4-1:0] node27075;
	wire [4-1:0] node27076;
	wire [4-1:0] node27079;
	wire [4-1:0] node27082;
	wire [4-1:0] node27084;
	wire [4-1:0] node27087;
	wire [4-1:0] node27088;
	wire [4-1:0] node27091;
	wire [4-1:0] node27094;
	wire [4-1:0] node27095;
	wire [4-1:0] node27096;
	wire [4-1:0] node27097;
	wire [4-1:0] node27099;
	wire [4-1:0] node27102;
	wire [4-1:0] node27103;
	wire [4-1:0] node27107;
	wire [4-1:0] node27108;
	wire [4-1:0] node27109;
	wire [4-1:0] node27110;
	wire [4-1:0] node27112;
	wire [4-1:0] node27113;
	wire [4-1:0] node27117;
	wire [4-1:0] node27118;
	wire [4-1:0] node27122;
	wire [4-1:0] node27123;
	wire [4-1:0] node27126;
	wire [4-1:0] node27128;
	wire [4-1:0] node27131;
	wire [4-1:0] node27132;
	wire [4-1:0] node27135;
	wire [4-1:0] node27138;
	wire [4-1:0] node27139;
	wire [4-1:0] node27140;
	wire [4-1:0] node27142;
	wire [4-1:0] node27145;
	wire [4-1:0] node27146;
	wire [4-1:0] node27150;
	wire [4-1:0] node27153;
	wire [4-1:0] node27154;
	wire [4-1:0] node27155;
	wire [4-1:0] node27156;
	wire [4-1:0] node27157;
	wire [4-1:0] node27158;
	wire [4-1:0] node27159;
	wire [4-1:0] node27162;
	wire [4-1:0] node27165;
	wire [4-1:0] node27166;
	wire [4-1:0] node27170;
	wire [4-1:0] node27171;
	wire [4-1:0] node27172;
	wire [4-1:0] node27175;
	wire [4-1:0] node27178;
	wire [4-1:0] node27181;
	wire [4-1:0] node27182;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27185;
	wire [4-1:0] node27186;
	wire [4-1:0] node27189;
	wire [4-1:0] node27193;
	wire [4-1:0] node27194;
	wire [4-1:0] node27198;
	wire [4-1:0] node27199;
	wire [4-1:0] node27200;
	wire [4-1:0] node27202;
	wire [4-1:0] node27206;
	wire [4-1:0] node27208;
	wire [4-1:0] node27209;
	wire [4-1:0] node27212;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27217;
	wire [4-1:0] node27220;
	wire [4-1:0] node27221;
	wire [4-1:0] node27225;
	wire [4-1:0] node27226;
	wire [4-1:0] node27227;
	wire [4-1:0] node27230;
	wire [4-1:0] node27231;
	wire [4-1:0] node27235;
	wire [4-1:0] node27238;
	wire [4-1:0] node27239;
	wire [4-1:0] node27240;
	wire [4-1:0] node27241;
	wire [4-1:0] node27242;
	wire [4-1:0] node27245;
	wire [4-1:0] node27248;
	wire [4-1:0] node27249;
	wire [4-1:0] node27252;
	wire [4-1:0] node27255;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27261;
	wire [4-1:0] node27264;
	wire [4-1:0] node27265;
	wire [4-1:0] node27266;
	wire [4-1:0] node27267;
	wire [4-1:0] node27270;
	wire [4-1:0] node27273;
	wire [4-1:0] node27275;
	wire [4-1:0] node27278;
	wire [4-1:0] node27279;
	wire [4-1:0] node27280;
	wire [4-1:0] node27283;
	wire [4-1:0] node27286;
	wire [4-1:0] node27288;
	wire [4-1:0] node27291;
	wire [4-1:0] node27292;
	wire [4-1:0] node27293;
	wire [4-1:0] node27294;
	wire [4-1:0] node27295;
	wire [4-1:0] node27299;
	wire [4-1:0] node27300;
	wire [4-1:0] node27304;
	wire [4-1:0] node27305;
	wire [4-1:0] node27306;
	wire [4-1:0] node27307;
	wire [4-1:0] node27310;
	wire [4-1:0] node27313;
	wire [4-1:0] node27315;
	wire [4-1:0] node27316;
	wire [4-1:0] node27320;
	wire [4-1:0] node27321;
	wire [4-1:0] node27324;
	wire [4-1:0] node27327;
	wire [4-1:0] node27328;
	wire [4-1:0] node27329;
	wire [4-1:0] node27331;
	wire [4-1:0] node27334;
	wire [4-1:0] node27335;
	wire [4-1:0] node27339;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27344;
	wire [4-1:0] node27345;
	wire [4-1:0] node27346;
	wire [4-1:0] node27347;
	wire [4-1:0] node27349;
	wire [4-1:0] node27352;
	wire [4-1:0] node27353;
	wire [4-1:0] node27354;
	wire [4-1:0] node27357;
	wire [4-1:0] node27360;
	wire [4-1:0] node27363;
	wire [4-1:0] node27364;
	wire [4-1:0] node27365;
	wire [4-1:0] node27368;
	wire [4-1:0] node27369;
	wire [4-1:0] node27373;
	wire [4-1:0] node27376;
	wire [4-1:0] node27377;
	wire [4-1:0] node27378;
	wire [4-1:0] node27379;
	wire [4-1:0] node27382;
	wire [4-1:0] node27385;
	wire [4-1:0] node27386;
	wire [4-1:0] node27387;
	wire [4-1:0] node27391;
	wire [4-1:0] node27392;
	wire [4-1:0] node27394;
	wire [4-1:0] node27397;
	wire [4-1:0] node27398;
	wire [4-1:0] node27402;
	wire [4-1:0] node27403;
	wire [4-1:0] node27404;
	wire [4-1:0] node27407;
	wire [4-1:0] node27408;
	wire [4-1:0] node27412;
	wire [4-1:0] node27415;
	wire [4-1:0] node27416;
	wire [4-1:0] node27417;
	wire [4-1:0] node27418;
	wire [4-1:0] node27420;
	wire [4-1:0] node27423;
	wire [4-1:0] node27424;
	wire [4-1:0] node27428;
	wire [4-1:0] node27429;
	wire [4-1:0] node27430;
	wire [4-1:0] node27431;
	wire [4-1:0] node27434;
	wire [4-1:0] node27437;
	wire [4-1:0] node27439;
	wire [4-1:0] node27440;
	wire [4-1:0] node27444;
	wire [4-1:0] node27445;
	wire [4-1:0] node27446;
	wire [4-1:0] node27447;
	wire [4-1:0] node27450;
	wire [4-1:0] node27451;
	wire [4-1:0] node27456;
	wire [4-1:0] node27457;
	wire [4-1:0] node27458;
	wire [4-1:0] node27462;
	wire [4-1:0] node27463;
	wire [4-1:0] node27465;
	wire [4-1:0] node27468;
	wire [4-1:0] node27469;
	wire [4-1:0] node27473;
	wire [4-1:0] node27474;
	wire [4-1:0] node27475;
	wire [4-1:0] node27477;
	wire [4-1:0] node27480;
	wire [4-1:0] node27481;
	wire [4-1:0] node27485;
	wire [4-1:0] node27488;
	wire [4-1:0] node27489;
	wire [4-1:0] node27490;
	wire [4-1:0] node27491;
	wire [4-1:0] node27492;
	wire [4-1:0] node27494;
	wire [4-1:0] node27497;
	wire [4-1:0] node27498;
	wire [4-1:0] node27501;
	wire [4-1:0] node27503;
	wire [4-1:0] node27505;
	wire [4-1:0] node27506;
	wire [4-1:0] node27509;
	wire [4-1:0] node27512;
	wire [4-1:0] node27513;
	wire [4-1:0] node27514;
	wire [4-1:0] node27515;
	wire [4-1:0] node27518;
	wire [4-1:0] node27521;
	wire [4-1:0] node27522;
	wire [4-1:0] node27523;
	wire [4-1:0] node27526;
	wire [4-1:0] node27529;
	wire [4-1:0] node27530;
	wire [4-1:0] node27532;
	wire [4-1:0] node27535;
	wire [4-1:0] node27536;
	wire [4-1:0] node27539;
	wire [4-1:0] node27542;
	wire [4-1:0] node27545;
	wire [4-1:0] node27546;
	wire [4-1:0] node27547;
	wire [4-1:0] node27548;
	wire [4-1:0] node27549;
	wire [4-1:0] node27551;
	wire [4-1:0] node27554;
	wire [4-1:0] node27555;
	wire [4-1:0] node27556;
	wire [4-1:0] node27559;
	wire [4-1:0] node27562;
	wire [4-1:0] node27565;
	wire [4-1:0] node27566;
	wire [4-1:0] node27569;
	wire [4-1:0] node27572;
	wire [4-1:0] node27573;
	wire [4-1:0] node27574;
	wire [4-1:0] node27575;
	wire [4-1:0] node27578;
	wire [4-1:0] node27582;
	wire [4-1:0] node27584;
	wire [4-1:0] node27585;
	wire [4-1:0] node27589;
	wire [4-1:0] node27590;
	wire [4-1:0] node27591;
	wire [4-1:0] node27592;
	wire [4-1:0] node27595;
	wire [4-1:0] node27598;
	wire [4-1:0] node27599;
	wire [4-1:0] node27600;
	wire [4-1:0] node27602;
	wire [4-1:0] node27605;
	wire [4-1:0] node27606;
	wire [4-1:0] node27610;
	wire [4-1:0] node27612;
	wire [4-1:0] node27615;
	wire [4-1:0] node27616;
	wire [4-1:0] node27617;
	wire [4-1:0] node27620;
	wire [4-1:0] node27623;
	wire [4-1:0] node27624;
	wire [4-1:0] node27625;
	wire [4-1:0] node27627;
	wire [4-1:0] node27630;
	wire [4-1:0] node27632;
	wire [4-1:0] node27635;
	wire [4-1:0] node27638;
	wire [4-1:0] node27639;
	wire [4-1:0] node27640;
	wire [4-1:0] node27641;
	wire [4-1:0] node27642;
	wire [4-1:0] node27645;
	wire [4-1:0] node27647;
	wire [4-1:0] node27650;
	wire [4-1:0] node27651;
	wire [4-1:0] node27654;
	wire [4-1:0] node27655;
	wire [4-1:0] node27657;
	wire [4-1:0] node27660;
	wire [4-1:0] node27662;
	wire [4-1:0] node27665;
	wire [4-1:0] node27666;
	wire [4-1:0] node27667;
	wire [4-1:0] node27668;
	wire [4-1:0] node27669;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27678;
	wire [4-1:0] node27680;
	wire [4-1:0] node27683;
	wire [4-1:0] node27684;
	wire [4-1:0] node27685;
	wire [4-1:0] node27689;
	wire [4-1:0] node27690;
	wire [4-1:0] node27693;
	wire [4-1:0] node27694;
	wire [4-1:0] node27698;
	wire [4-1:0] node27699;
	wire [4-1:0] node27700;
	wire [4-1:0] node27701;
	wire [4-1:0] node27704;
	wire [4-1:0] node27706;
	wire [4-1:0] node27710;
	wire [4-1:0] node27711;
	wire [4-1:0] node27712;
	wire [4-1:0] node27714;
	wire [4-1:0] node27719;
	wire [4-1:0] node27720;
	wire [4-1:0] node27721;
	wire [4-1:0] node27722;
	wire [4-1:0] node27723;
	wire [4-1:0] node27724;
	wire [4-1:0] node27725;
	wire [4-1:0] node27726;
	wire [4-1:0] node27727;
	wire [4-1:0] node27729;
	wire [4-1:0] node27730;
	wire [4-1:0] node27734;
	wire [4-1:0] node27735;
	wire [4-1:0] node27737;
	wire [4-1:0] node27740;
	wire [4-1:0] node27743;
	wire [4-1:0] node27744;
	wire [4-1:0] node27747;
	wire [4-1:0] node27748;
	wire [4-1:0] node27749;
	wire [4-1:0] node27750;
	wire [4-1:0] node27756;
	wire [4-1:0] node27757;
	wire [4-1:0] node27758;
	wire [4-1:0] node27759;
	wire [4-1:0] node27760;
	wire [4-1:0] node27764;
	wire [4-1:0] node27767;
	wire [4-1:0] node27768;
	wire [4-1:0] node27771;
	wire [4-1:0] node27774;
	wire [4-1:0] node27775;
	wire [4-1:0] node27776;
	wire [4-1:0] node27778;
	wire [4-1:0] node27779;
	wire [4-1:0] node27782;
	wire [4-1:0] node27785;
	wire [4-1:0] node27786;
	wire [4-1:0] node27789;
	wire [4-1:0] node27792;
	wire [4-1:0] node27793;
	wire [4-1:0] node27794;
	wire [4-1:0] node27798;
	wire [4-1:0] node27801;
	wire [4-1:0] node27802;
	wire [4-1:0] node27803;
	wire [4-1:0] node27804;
	wire [4-1:0] node27805;
	wire [4-1:0] node27806;
	wire [4-1:0] node27809;
	wire [4-1:0] node27811;
	wire [4-1:0] node27814;
	wire [4-1:0] node27815;
	wire [4-1:0] node27818;
	wire [4-1:0] node27821;
	wire [4-1:0] node27822;
	wire [4-1:0] node27824;
	wire [4-1:0] node27827;
	wire [4-1:0] node27828;
	wire [4-1:0] node27829;
	wire [4-1:0] node27833;
	wire [4-1:0] node27836;
	wire [4-1:0] node27837;
	wire [4-1:0] node27838;
	wire [4-1:0] node27839;
	wire [4-1:0] node27842;
	wire [4-1:0] node27846;
	wire [4-1:0] node27847;
	wire [4-1:0] node27848;
	wire [4-1:0] node27849;
	wire [4-1:0] node27852;
	wire [4-1:0] node27855;
	wire [4-1:0] node27856;
	wire [4-1:0] node27859;
	wire [4-1:0] node27862;
	wire [4-1:0] node27865;
	wire [4-1:0] node27866;
	wire [4-1:0] node27867;
	wire [4-1:0] node27868;
	wire [4-1:0] node27871;
	wire [4-1:0] node27872;
	wire [4-1:0] node27875;
	wire [4-1:0] node27876;
	wire [4-1:0] node27879;
	wire [4-1:0] node27882;
	wire [4-1:0] node27883;
	wire [4-1:0] node27887;
	wire [4-1:0] node27888;
	wire [4-1:0] node27890;
	wire [4-1:0] node27891;
	wire [4-1:0] node27892;
	wire [4-1:0] node27897;
	wire [4-1:0] node27898;
	wire [4-1:0] node27901;
	wire [4-1:0] node27902;
	wire [4-1:0] node27905;
	wire [4-1:0] node27906;
	wire [4-1:0] node27910;
	wire [4-1:0] node27911;
	wire [4-1:0] node27912;
	wire [4-1:0] node27913;
	wire [4-1:0] node27914;
	wire [4-1:0] node27915;
	wire [4-1:0] node27916;
	wire [4-1:0] node27917;
	wire [4-1:0] node27921;
	wire [4-1:0] node27925;
	wire [4-1:0] node27926;
	wire [4-1:0] node27929;
	wire [4-1:0] node27932;
	wire [4-1:0] node27933;
	wire [4-1:0] node27935;
	wire [4-1:0] node27938;
	wire [4-1:0] node27939;
	wire [4-1:0] node27942;
	wire [4-1:0] node27943;
	wire [4-1:0] node27945;
	wire [4-1:0] node27948;
	wire [4-1:0] node27951;
	wire [4-1:0] node27952;
	wire [4-1:0] node27953;
	wire [4-1:0] node27955;
	wire [4-1:0] node27956;
	wire [4-1:0] node27959;
	wire [4-1:0] node27962;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27968;
	wire [4-1:0] node27970;
	wire [4-1:0] node27973;
	wire [4-1:0] node27974;
	wire [4-1:0] node27975;
	wire [4-1:0] node27978;
	wire [4-1:0] node27979;
	wire [4-1:0] node27982;
	wire [4-1:0] node27985;
	wire [4-1:0] node27986;
	wire [4-1:0] node27989;
	wire [4-1:0] node27991;
	wire [4-1:0] node27994;
	wire [4-1:0] node27995;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node28000;
	wire [4-1:0] node28003;
	wire [4-1:0] node28006;
	wire [4-1:0] node28007;
	wire [4-1:0] node28008;
	wire [4-1:0] node28009;
	wire [4-1:0] node28013;
	wire [4-1:0] node28014;
	wire [4-1:0] node28018;
	wire [4-1:0] node28020;
	wire [4-1:0] node28023;
	wire [4-1:0] node28024;
	wire [4-1:0] node28026;
	wire [4-1:0] node28028;
	wire [4-1:0] node28031;
	wire [4-1:0] node28032;
	wire [4-1:0] node28033;
	wire [4-1:0] node28035;
	wire [4-1:0] node28040;
	wire [4-1:0] node28041;
	wire [4-1:0] node28042;
	wire [4-1:0] node28043;
	wire [4-1:0] node28046;
	wire [4-1:0] node28049;
	wire [4-1:0] node28050;
	wire [4-1:0] node28052;
	wire [4-1:0] node28056;
	wire [4-1:0] node28057;
	wire [4-1:0] node28058;
	wire [4-1:0] node28059;
	wire [4-1:0] node28062;
	wire [4-1:0] node28066;
	wire [4-1:0] node28069;
	wire [4-1:0] node28070;
	wire [4-1:0] node28071;
	wire [4-1:0] node28072;
	wire [4-1:0] node28073;
	wire [4-1:0] node28074;
	wire [4-1:0] node28075;
	wire [4-1:0] node28076;
	wire [4-1:0] node28078;
	wire [4-1:0] node28082;
	wire [4-1:0] node28086;
	wire [4-1:0] node28087;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28092;
	wire [4-1:0] node28095;
	wire [4-1:0] node28098;
	wire [4-1:0] node28099;
	wire [4-1:0] node28100;
	wire [4-1:0] node28102;
	wire [4-1:0] node28105;
	wire [4-1:0] node28108;
	wire [4-1:0] node28110;
	wire [4-1:0] node28111;
	wire [4-1:0] node28115;
	wire [4-1:0] node28116;
	wire [4-1:0] node28117;
	wire [4-1:0] node28118;
	wire [4-1:0] node28119;
	wire [4-1:0] node28123;
	wire [4-1:0] node28124;
	wire [4-1:0] node28126;
	wire [4-1:0] node28129;
	wire [4-1:0] node28132;
	wire [4-1:0] node28133;
	wire [4-1:0] node28134;
	wire [4-1:0] node28135;
	wire [4-1:0] node28138;
	wire [4-1:0] node28141;
	wire [4-1:0] node28145;
	wire [4-1:0] node28146;
	wire [4-1:0] node28148;
	wire [4-1:0] node28149;
	wire [4-1:0] node28153;
	wire [4-1:0] node28154;
	wire [4-1:0] node28155;
	wire [4-1:0] node28158;
	wire [4-1:0] node28162;
	wire [4-1:0] node28163;
	wire [4-1:0] node28164;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28168;
	wire [4-1:0] node28171;
	wire [4-1:0] node28172;
	wire [4-1:0] node28175;
	wire [4-1:0] node28176;
	wire [4-1:0] node28180;
	wire [4-1:0] node28181;
	wire [4-1:0] node28184;
	wire [4-1:0] node28186;
	wire [4-1:0] node28187;
	wire [4-1:0] node28190;
	wire [4-1:0] node28193;
	wire [4-1:0] node28194;
	wire [4-1:0] node28195;
	wire [4-1:0] node28198;
	wire [4-1:0] node28199;
	wire [4-1:0] node28200;
	wire [4-1:0] node28203;
	wire [4-1:0] node28206;
	wire [4-1:0] node28207;
	wire [4-1:0] node28211;
	wire [4-1:0] node28212;
	wire [4-1:0] node28213;
	wire [4-1:0] node28217;
	wire [4-1:0] node28218;
	wire [4-1:0] node28219;
	wire [4-1:0] node28222;
	wire [4-1:0] node28226;
	wire [4-1:0] node28227;
	wire [4-1:0] node28228;
	wire [4-1:0] node28229;
	wire [4-1:0] node28230;
	wire [4-1:0] node28234;
	wire [4-1:0] node28235;
	wire [4-1:0] node28236;
	wire [4-1:0] node28240;
	wire [4-1:0] node28243;
	wire [4-1:0] node28244;
	wire [4-1:0] node28246;
	wire [4-1:0] node28249;
	wire [4-1:0] node28250;
	wire [4-1:0] node28253;
	wire [4-1:0] node28256;
	wire [4-1:0] node28257;
	wire [4-1:0] node28258;
	wire [4-1:0] node28261;
	wire [4-1:0] node28263;
	wire [4-1:0] node28264;
	wire [4-1:0] node28267;
	wire [4-1:0] node28270;
	wire [4-1:0] node28271;
	wire [4-1:0] node28273;
	wire [4-1:0] node28276;
	wire [4-1:0] node28277;
	wire [4-1:0] node28281;
	wire [4-1:0] node28282;
	wire [4-1:0] node28283;
	wire [4-1:0] node28284;
	wire [4-1:0] node28285;
	wire [4-1:0] node28286;
	wire [4-1:0] node28288;
	wire [4-1:0] node28289;
	wire [4-1:0] node28292;
	wire [4-1:0] node28295;
	wire [4-1:0] node28296;
	wire [4-1:0] node28297;
	wire [4-1:0] node28301;
	wire [4-1:0] node28304;
	wire [4-1:0] node28305;
	wire [4-1:0] node28308;
	wire [4-1:0] node28309;
	wire [4-1:0] node28312;
	wire [4-1:0] node28313;
	wire [4-1:0] node28316;
	wire [4-1:0] node28319;
	wire [4-1:0] node28320;
	wire [4-1:0] node28321;
	wire [4-1:0] node28323;
	wire [4-1:0] node28324;
	wire [4-1:0] node28327;
	wire [4-1:0] node28330;
	wire [4-1:0] node28332;
	wire [4-1:0] node28335;
	wire [4-1:0] node28336;
	wire [4-1:0] node28339;
	wire [4-1:0] node28341;
	wire [4-1:0] node28344;
	wire [4-1:0] node28345;
	wire [4-1:0] node28346;
	wire [4-1:0] node28347;
	wire [4-1:0] node28350;
	wire [4-1:0] node28352;
	wire [4-1:0] node28353;
	wire [4-1:0] node28357;
	wire [4-1:0] node28359;
	wire [4-1:0] node28362;
	wire [4-1:0] node28363;
	wire [4-1:0] node28365;
	wire [4-1:0] node28366;
	wire [4-1:0] node28370;
	wire [4-1:0] node28371;
	wire [4-1:0] node28372;
	wire [4-1:0] node28375;
	wire [4-1:0] node28378;
	wire [4-1:0] node28381;
	wire [4-1:0] node28382;
	wire [4-1:0] node28383;
	wire [4-1:0] node28384;
	wire [4-1:0] node28385;
	wire [4-1:0] node28386;
	wire [4-1:0] node28389;
	wire [4-1:0] node28392;
	wire [4-1:0] node28393;
	wire [4-1:0] node28395;
	wire [4-1:0] node28399;
	wire [4-1:0] node28401;
	wire [4-1:0] node28402;
	wire [4-1:0] node28403;
	wire [4-1:0] node28406;
	wire [4-1:0] node28409;
	wire [4-1:0] node28411;
	wire [4-1:0] node28414;
	wire [4-1:0] node28415;
	wire [4-1:0] node28416;
	wire [4-1:0] node28418;
	wire [4-1:0] node28419;
	wire [4-1:0] node28422;
	wire [4-1:0] node28425;
	wire [4-1:0] node28426;
	wire [4-1:0] node28427;
	wire [4-1:0] node28430;
	wire [4-1:0] node28433;
	wire [4-1:0] node28434;
	wire [4-1:0] node28437;
	wire [4-1:0] node28440;
	wire [4-1:0] node28442;
	wire [4-1:0] node28443;
	wire [4-1:0] node28446;
	wire [4-1:0] node28449;
	wire [4-1:0] node28450;
	wire [4-1:0] node28451;
	wire [4-1:0] node28452;
	wire [4-1:0] node28455;
	wire [4-1:0] node28457;
	wire [4-1:0] node28459;
	wire [4-1:0] node28462;
	wire [4-1:0] node28463;
	wire [4-1:0] node28465;
	wire [4-1:0] node28469;
	wire [4-1:0] node28471;
	wire [4-1:0] node28472;
	wire [4-1:0] node28473;
	wire [4-1:0] node28476;
	wire [4-1:0] node28479;
	wire [4-1:0] node28480;
	wire [4-1:0] node28483;
	wire [4-1:0] node28486;
	wire [4-1:0] node28487;
	wire [4-1:0] node28488;
	wire [4-1:0] node28489;
	wire [4-1:0] node28490;
	wire [4-1:0] node28491;
	wire [4-1:0] node28492;
	wire [4-1:0] node28493;
	wire [4-1:0] node28495;
	wire [4-1:0] node28498;
	wire [4-1:0] node28499;
	wire [4-1:0] node28501;
	wire [4-1:0] node28504;
	wire [4-1:0] node28505;
	wire [4-1:0] node28509;
	wire [4-1:0] node28510;
	wire [4-1:0] node28512;
	wire [4-1:0] node28515;
	wire [4-1:0] node28516;
	wire [4-1:0] node28520;
	wire [4-1:0] node28521;
	wire [4-1:0] node28523;
	wire [4-1:0] node28525;
	wire [4-1:0] node28528;
	wire [4-1:0] node28531;
	wire [4-1:0] node28532;
	wire [4-1:0] node28533;
	wire [4-1:0] node28534;
	wire [4-1:0] node28536;
	wire [4-1:0] node28538;
	wire [4-1:0] node28542;
	wire [4-1:0] node28543;
	wire [4-1:0] node28546;
	wire [4-1:0] node28548;
	wire [4-1:0] node28551;
	wire [4-1:0] node28552;
	wire [4-1:0] node28554;
	wire [4-1:0] node28555;
	wire [4-1:0] node28558;
	wire [4-1:0] node28561;
	wire [4-1:0] node28562;
	wire [4-1:0] node28563;
	wire [4-1:0] node28567;
	wire [4-1:0] node28568;
	wire [4-1:0] node28571;
	wire [4-1:0] node28574;
	wire [4-1:0] node28575;
	wire [4-1:0] node28576;
	wire [4-1:0] node28577;
	wire [4-1:0] node28579;
	wire [4-1:0] node28582;
	wire [4-1:0] node28583;
	wire [4-1:0] node28585;
	wire [4-1:0] node28588;
	wire [4-1:0] node28591;
	wire [4-1:0] node28592;
	wire [4-1:0] node28594;
	wire [4-1:0] node28595;
	wire [4-1:0] node28598;
	wire [4-1:0] node28601;
	wire [4-1:0] node28602;
	wire [4-1:0] node28603;
	wire [4-1:0] node28604;
	wire [4-1:0] node28609;
	wire [4-1:0] node28610;
	wire [4-1:0] node28614;
	wire [4-1:0] node28615;
	wire [4-1:0] node28616;
	wire [4-1:0] node28617;
	wire [4-1:0] node28619;
	wire [4-1:0] node28623;
	wire [4-1:0] node28625;
	wire [4-1:0] node28628;
	wire [4-1:0] node28629;
	wire [4-1:0] node28630;
	wire [4-1:0] node28632;
	wire [4-1:0] node28636;
	wire [4-1:0] node28637;
	wire [4-1:0] node28638;
	wire [4-1:0] node28641;
	wire [4-1:0] node28642;
	wire [4-1:0] node28646;
	wire [4-1:0] node28647;
	wire [4-1:0] node28648;
	wire [4-1:0] node28653;
	wire [4-1:0] node28654;
	wire [4-1:0] node28655;
	wire [4-1:0] node28656;
	wire [4-1:0] node28657;
	wire [4-1:0] node28658;
	wire [4-1:0] node28660;
	wire [4-1:0] node28662;
	wire [4-1:0] node28665;
	wire [4-1:0] node28668;
	wire [4-1:0] node28669;
	wire [4-1:0] node28672;
	wire [4-1:0] node28675;
	wire [4-1:0] node28676;
	wire [4-1:0] node28677;
	wire [4-1:0] node28679;
	wire [4-1:0] node28680;
	wire [4-1:0] node28683;
	wire [4-1:0] node28686;
	wire [4-1:0] node28687;
	wire [4-1:0] node28691;
	wire [4-1:0] node28692;
	wire [4-1:0] node28693;
	wire [4-1:0] node28698;
	wire [4-1:0] node28699;
	wire [4-1:0] node28700;
	wire [4-1:0] node28701;
	wire [4-1:0] node28702;
	wire [4-1:0] node28706;
	wire [4-1:0] node28708;
	wire [4-1:0] node28711;
	wire [4-1:0] node28712;
	wire [4-1:0] node28714;
	wire [4-1:0] node28715;
	wire [4-1:0] node28719;
	wire [4-1:0] node28720;
	wire [4-1:0] node28721;
	wire [4-1:0] node28725;
	wire [4-1:0] node28726;
	wire [4-1:0] node28730;
	wire [4-1:0] node28731;
	wire [4-1:0] node28732;
	wire [4-1:0] node28733;
	wire [4-1:0] node28736;
	wire [4-1:0] node28739;
	wire [4-1:0] node28742;
	wire [4-1:0] node28743;
	wire [4-1:0] node28744;
	wire [4-1:0] node28747;
	wire [4-1:0] node28750;
	wire [4-1:0] node28751;
	wire [4-1:0] node28755;
	wire [4-1:0] node28756;
	wire [4-1:0] node28757;
	wire [4-1:0] node28758;
	wire [4-1:0] node28759;
	wire [4-1:0] node28760;
	wire [4-1:0] node28761;
	wire [4-1:0] node28765;
	wire [4-1:0] node28766;
	wire [4-1:0] node28769;
	wire [4-1:0] node28772;
	wire [4-1:0] node28775;
	wire [4-1:0] node28776;
	wire [4-1:0] node28778;
	wire [4-1:0] node28781;
	wire [4-1:0] node28782;
	wire [4-1:0] node28786;
	wire [4-1:0] node28787;
	wire [4-1:0] node28788;
	wire [4-1:0] node28789;
	wire [4-1:0] node28792;
	wire [4-1:0] node28795;
	wire [4-1:0] node28797;
	wire [4-1:0] node28799;
	wire [4-1:0] node28802;
	wire [4-1:0] node28803;
	wire [4-1:0] node28804;
	wire [4-1:0] node28807;
	wire [4-1:0] node28810;
	wire [4-1:0] node28811;
	wire [4-1:0] node28815;
	wire [4-1:0] node28816;
	wire [4-1:0] node28817;
	wire [4-1:0] node28818;
	wire [4-1:0] node28820;
	wire [4-1:0] node28824;
	wire [4-1:0] node28825;
	wire [4-1:0] node28828;
	wire [4-1:0] node28831;
	wire [4-1:0] node28832;
	wire [4-1:0] node28833;
	wire [4-1:0] node28834;
	wire [4-1:0] node28836;
	wire [4-1:0] node28841;
	wire [4-1:0] node28842;
	wire [4-1:0] node28846;
	wire [4-1:0] node28847;
	wire [4-1:0] node28848;
	wire [4-1:0] node28849;
	wire [4-1:0] node28850;
	wire [4-1:0] node28851;
	wire [4-1:0] node28852;
	wire [4-1:0] node28853;
	wire [4-1:0] node28856;
	wire [4-1:0] node28859;
	wire [4-1:0] node28860;
	wire [4-1:0] node28861;
	wire [4-1:0] node28865;
	wire [4-1:0] node28868;
	wire [4-1:0] node28869;
	wire [4-1:0] node28870;
	wire [4-1:0] node28873;
	wire [4-1:0] node28877;
	wire [4-1:0] node28878;
	wire [4-1:0] node28880;
	wire [4-1:0] node28881;
	wire [4-1:0] node28883;
	wire [4-1:0] node28886;
	wire [4-1:0] node28889;
	wire [4-1:0] node28890;
	wire [4-1:0] node28892;
	wire [4-1:0] node28895;
	wire [4-1:0] node28896;
	wire [4-1:0] node28899;
	wire [4-1:0] node28900;
	wire [4-1:0] node28903;
	wire [4-1:0] node28906;
	wire [4-1:0] node28907;
	wire [4-1:0] node28908;
	wire [4-1:0] node28909;
	wire [4-1:0] node28910;
	wire [4-1:0] node28913;
	wire [4-1:0] node28914;
	wire [4-1:0] node28917;
	wire [4-1:0] node28920;
	wire [4-1:0] node28922;
	wire [4-1:0] node28923;
	wire [4-1:0] node28927;
	wire [4-1:0] node28928;
	wire [4-1:0] node28931;
	wire [4-1:0] node28932;
	wire [4-1:0] node28936;
	wire [4-1:0] node28937;
	wire [4-1:0] node28938;
	wire [4-1:0] node28939;
	wire [4-1:0] node28943;
	wire [4-1:0] node28946;
	wire [4-1:0] node28947;
	wire [4-1:0] node28948;
	wire [4-1:0] node28949;
	wire [4-1:0] node28953;
	wire [4-1:0] node28954;
	wire [4-1:0] node28958;
	wire [4-1:0] node28959;
	wire [4-1:0] node28962;
	wire [4-1:0] node28964;
	wire [4-1:0] node28967;
	wire [4-1:0] node28968;
	wire [4-1:0] node28969;
	wire [4-1:0] node28970;
	wire [4-1:0] node28971;
	wire [4-1:0] node28973;
	wire [4-1:0] node28974;
	wire [4-1:0] node28977;
	wire [4-1:0] node28980;
	wire [4-1:0] node28981;
	wire [4-1:0] node28982;
	wire [4-1:0] node28985;
	wire [4-1:0] node28989;
	wire [4-1:0] node28990;
	wire [4-1:0] node28993;
	wire [4-1:0] node28996;
	wire [4-1:0] node28997;
	wire [4-1:0] node28998;
	wire [4-1:0] node29000;
	wire [4-1:0] node29002;
	wire [4-1:0] node29006;
	wire [4-1:0] node29008;
	wire [4-1:0] node29010;
	wire [4-1:0] node29013;
	wire [4-1:0] node29014;
	wire [4-1:0] node29015;
	wire [4-1:0] node29016;
	wire [4-1:0] node29017;
	wire [4-1:0] node29019;
	wire [4-1:0] node29022;
	wire [4-1:0] node29025;
	wire [4-1:0] node29026;
	wire [4-1:0] node29027;
	wire [4-1:0] node29031;
	wire [4-1:0] node29034;
	wire [4-1:0] node29035;
	wire [4-1:0] node29036;
	wire [4-1:0] node29039;
	wire [4-1:0] node29040;
	wire [4-1:0] node29044;
	wire [4-1:0] node29045;
	wire [4-1:0] node29046;
	wire [4-1:0] node29051;
	wire [4-1:0] node29052;
	wire [4-1:0] node29053;
	wire [4-1:0] node29055;
	wire [4-1:0] node29058;
	wire [4-1:0] node29060;
	wire [4-1:0] node29063;
	wire [4-1:0] node29064;
	wire [4-1:0] node29065;
	wire [4-1:0] node29068;
	wire [4-1:0] node29071;
	wire [4-1:0] node29072;
	wire [4-1:0] node29073;
	wire [4-1:0] node29078;
	wire [4-1:0] node29079;
	wire [4-1:0] node29080;
	wire [4-1:0] node29081;
	wire [4-1:0] node29082;
	wire [4-1:0] node29083;
	wire [4-1:0] node29084;
	wire [4-1:0] node29087;
	wire [4-1:0] node29090;
	wire [4-1:0] node29091;
	wire [4-1:0] node29095;
	wire [4-1:0] node29096;
	wire [4-1:0] node29099;
	wire [4-1:0] node29100;
	wire [4-1:0] node29104;
	wire [4-1:0] node29105;
	wire [4-1:0] node29106;
	wire [4-1:0] node29108;
	wire [4-1:0] node29111;
	wire [4-1:0] node29113;
	wire [4-1:0] node29116;
	wire [4-1:0] node29117;
	wire [4-1:0] node29118;
	wire [4-1:0] node29122;
	wire [4-1:0] node29124;
	wire [4-1:0] node29127;
	wire [4-1:0] node29128;
	wire [4-1:0] node29129;
	wire [4-1:0] node29130;
	wire [4-1:0] node29133;
	wire [4-1:0] node29136;
	wire [4-1:0] node29139;
	wire [4-1:0] node29140;
	wire [4-1:0] node29141;
	wire [4-1:0] node29143;
	wire [4-1:0] node29145;
	wire [4-1:0] node29148;
	wire [4-1:0] node29150;
	wire [4-1:0] node29153;
	wire [4-1:0] node29154;
	wire [4-1:0] node29155;
	wire [4-1:0] node29158;
	wire [4-1:0] node29161;
	wire [4-1:0] node29162;
	wire [4-1:0] node29165;
	wire [4-1:0] node29168;
	wire [4-1:0] node29169;
	wire [4-1:0] node29170;
	wire [4-1:0] node29171;
	wire [4-1:0] node29172;
	wire [4-1:0] node29174;
	wire [4-1:0] node29177;
	wire [4-1:0] node29178;
	wire [4-1:0] node29181;
	wire [4-1:0] node29184;
	wire [4-1:0] node29185;
	wire [4-1:0] node29187;
	wire [4-1:0] node29191;
	wire [4-1:0] node29192;
	wire [4-1:0] node29194;
	wire [4-1:0] node29196;
	wire [4-1:0] node29199;
	wire [4-1:0] node29200;
	wire [4-1:0] node29201;
	wire [4-1:0] node29205;
	wire [4-1:0] node29206;
	wire [4-1:0] node29209;
	wire [4-1:0] node29212;
	wire [4-1:0] node29213;
	wire [4-1:0] node29214;
	wire [4-1:0] node29216;
	wire [4-1:0] node29217;
	wire [4-1:0] node29220;
	wire [4-1:0] node29223;
	wire [4-1:0] node29224;
	wire [4-1:0] node29227;
	wire [4-1:0] node29230;
	wire [4-1:0] node29231;
	wire [4-1:0] node29232;
	wire [4-1:0] node29233;
	wire [4-1:0] node29237;
	wire [4-1:0] node29238;
	wire [4-1:0] node29242;
	wire [4-1:0] node29243;
	wire [4-1:0] node29244;
	wire [4-1:0] node29245;
	wire [4-1:0] node29250;
	wire [4-1:0] node29252;
	wire [4-1:0] node29253;
	wire [4-1:0] node29257;
	wire [4-1:0] node29258;
	wire [4-1:0] node29259;
	wire [4-1:0] node29260;
	wire [4-1:0] node29261;
	wire [4-1:0] node29262;
	wire [4-1:0] node29263;
	wire [4-1:0] node29264;
	wire [4-1:0] node29265;
	wire [4-1:0] node29267;
	wire [4-1:0] node29270;
	wire [4-1:0] node29272;
	wire [4-1:0] node29275;
	wire [4-1:0] node29276;
	wire [4-1:0] node29279;
	wire [4-1:0] node29280;
	wire [4-1:0] node29283;
	wire [4-1:0] node29286;
	wire [4-1:0] node29287;
	wire [4-1:0] node29290;
	wire [4-1:0] node29293;
	wire [4-1:0] node29294;
	wire [4-1:0] node29295;
	wire [4-1:0] node29298;
	wire [4-1:0] node29301;
	wire [4-1:0] node29303;
	wire [4-1:0] node29304;
	wire [4-1:0] node29307;
	wire [4-1:0] node29310;
	wire [4-1:0] node29311;
	wire [4-1:0] node29312;
	wire [4-1:0] node29313;
	wire [4-1:0] node29314;
	wire [4-1:0] node29316;
	wire [4-1:0] node29319;
	wire [4-1:0] node29321;
	wire [4-1:0] node29324;
	wire [4-1:0] node29325;
	wire [4-1:0] node29327;
	wire [4-1:0] node29331;
	wire [4-1:0] node29332;
	wire [4-1:0] node29334;
	wire [4-1:0] node29336;
	wire [4-1:0] node29337;
	wire [4-1:0] node29341;
	wire [4-1:0] node29342;
	wire [4-1:0] node29344;
	wire [4-1:0] node29345;
	wire [4-1:0] node29348;
	wire [4-1:0] node29351;
	wire [4-1:0] node29352;
	wire [4-1:0] node29355;
	wire [4-1:0] node29358;
	wire [4-1:0] node29359;
	wire [4-1:0] node29360;
	wire [4-1:0] node29362;
	wire [4-1:0] node29365;
	wire [4-1:0] node29367;
	wire [4-1:0] node29370;
	wire [4-1:0] node29371;
	wire [4-1:0] node29373;
	wire [4-1:0] node29376;
	wire [4-1:0] node29378;
	wire [4-1:0] node29381;
	wire [4-1:0] node29382;
	wire [4-1:0] node29383;
	wire [4-1:0] node29384;
	wire [4-1:0] node29386;
	wire [4-1:0] node29387;
	wire [4-1:0] node29390;
	wire [4-1:0] node29393;
	wire [4-1:0] node29394;
	wire [4-1:0] node29395;
	wire [4-1:0] node29399;
	wire [4-1:0] node29400;
	wire [4-1:0] node29401;
	wire [4-1:0] node29405;
	wire [4-1:0] node29406;
	wire [4-1:0] node29407;
	wire [4-1:0] node29412;
	wire [4-1:0] node29413;
	wire [4-1:0] node29414;
	wire [4-1:0] node29415;
	wire [4-1:0] node29418;
	wire [4-1:0] node29421;
	wire [4-1:0] node29424;
	wire [4-1:0] node29425;
	wire [4-1:0] node29426;
	wire [4-1:0] node29429;
	wire [4-1:0] node29430;
	wire [4-1:0] node29435;
	wire [4-1:0] node29436;
	wire [4-1:0] node29437;
	wire [4-1:0] node29439;
	wire [4-1:0] node29440;
	wire [4-1:0] node29442;
	wire [4-1:0] node29443;
	wire [4-1:0] node29447;
	wire [4-1:0] node29448;
	wire [4-1:0] node29452;
	wire [4-1:0] node29453;
	wire [4-1:0] node29455;
	wire [4-1:0] node29456;
	wire [4-1:0] node29457;
	wire [4-1:0] node29461;
	wire [4-1:0] node29462;
	wire [4-1:0] node29466;
	wire [4-1:0] node29467;
	wire [4-1:0] node29468;
	wire [4-1:0] node29469;
	wire [4-1:0] node29472;
	wire [4-1:0] node29476;
	wire [4-1:0] node29478;
	wire [4-1:0] node29481;
	wire [4-1:0] node29482;
	wire [4-1:0] node29483;
	wire [4-1:0] node29484;
	wire [4-1:0] node29485;
	wire [4-1:0] node29488;
	wire [4-1:0] node29491;
	wire [4-1:0] node29492;
	wire [4-1:0] node29496;
	wire [4-1:0] node29497;
	wire [4-1:0] node29500;
	wire [4-1:0] node29503;
	wire [4-1:0] node29504;
	wire [4-1:0] node29505;
	wire [4-1:0] node29507;
	wire [4-1:0] node29509;
	wire [4-1:0] node29512;
	wire [4-1:0] node29515;
	wire [4-1:0] node29516;
	wire [4-1:0] node29519;
	wire [4-1:0] node29521;
	wire [4-1:0] node29524;
	wire [4-1:0] node29525;
	wire [4-1:0] node29526;
	wire [4-1:0] node29527;
	wire [4-1:0] node29528;
	wire [4-1:0] node29529;
	wire [4-1:0] node29530;
	wire [4-1:0] node29534;
	wire [4-1:0] node29535;
	wire [4-1:0] node29539;
	wire [4-1:0] node29541;
	wire [4-1:0] node29542;
	wire [4-1:0] node29546;
	wire [4-1:0] node29547;
	wire [4-1:0] node29548;
	wire [4-1:0] node29550;
	wire [4-1:0] node29553;
	wire [4-1:0] node29554;
	wire [4-1:0] node29558;
	wire [4-1:0] node29559;
	wire [4-1:0] node29561;
	wire [4-1:0] node29564;
	wire [4-1:0] node29566;
	wire [4-1:0] node29569;
	wire [4-1:0] node29570;
	wire [4-1:0] node29571;
	wire [4-1:0] node29573;
	wire [4-1:0] node29576;
	wire [4-1:0] node29578;
	wire [4-1:0] node29581;
	wire [4-1:0] node29582;
	wire [4-1:0] node29583;
	wire [4-1:0] node29587;
	wire [4-1:0] node29588;
	wire [4-1:0] node29592;
	wire [4-1:0] node29593;
	wire [4-1:0] node29594;
	wire [4-1:0] node29595;
	wire [4-1:0] node29596;
	wire [4-1:0] node29597;
	wire [4-1:0] node29599;
	wire [4-1:0] node29602;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29609;
	wire [4-1:0] node29610;
	wire [4-1:0] node29614;
	wire [4-1:0] node29615;
	wire [4-1:0] node29618;
	wire [4-1:0] node29621;
	wire [4-1:0] node29622;
	wire [4-1:0] node29623;
	wire [4-1:0] node29624;
	wire [4-1:0] node29625;
	wire [4-1:0] node29628;
	wire [4-1:0] node29631;
	wire [4-1:0] node29632;
	wire [4-1:0] node29633;
	wire [4-1:0] node29636;
	wire [4-1:0] node29640;
	wire [4-1:0] node29642;
	wire [4-1:0] node29645;
	wire [4-1:0] node29646;
	wire [4-1:0] node29647;
	wire [4-1:0] node29650;
	wire [4-1:0] node29652;
	wire [4-1:0] node29654;
	wire [4-1:0] node29657;
	wire [4-1:0] node29658;
	wire [4-1:0] node29661;
	wire [4-1:0] node29664;
	wire [4-1:0] node29665;
	wire [4-1:0] node29666;
	wire [4-1:0] node29667;
	wire [4-1:0] node29668;
	wire [4-1:0] node29669;
	wire [4-1:0] node29671;
	wire [4-1:0] node29674;
	wire [4-1:0] node29676;
	wire [4-1:0] node29680;
	wire [4-1:0] node29681;
	wire [4-1:0] node29684;
	wire [4-1:0] node29687;
	wire [4-1:0] node29688;
	wire [4-1:0] node29691;
	wire [4-1:0] node29694;
	wire [4-1:0] node29695;
	wire [4-1:0] node29696;
	wire [4-1:0] node29698;
	wire [4-1:0] node29701;
	wire [4-1:0] node29702;
	wire [4-1:0] node29705;
	wire [4-1:0] node29708;
	wire [4-1:0] node29709;
	wire [4-1:0] node29712;
	wire [4-1:0] node29715;
	wire [4-1:0] node29716;
	wire [4-1:0] node29717;
	wire [4-1:0] node29718;
	wire [4-1:0] node29719;
	wire [4-1:0] node29720;
	wire [4-1:0] node29721;
	wire [4-1:0] node29722;
	wire [4-1:0] node29724;
	wire [4-1:0] node29727;
	wire [4-1:0] node29728;
	wire [4-1:0] node29732;
	wire [4-1:0] node29733;
	wire [4-1:0] node29737;
	wire [4-1:0] node29738;
	wire [4-1:0] node29741;
	wire [4-1:0] node29742;
	wire [4-1:0] node29743;
	wire [4-1:0] node29747;
	wire [4-1:0] node29748;
	wire [4-1:0] node29752;
	wire [4-1:0] node29753;
	wire [4-1:0] node29754;
	wire [4-1:0] node29756;
	wire [4-1:0] node29757;
	wire [4-1:0] node29760;
	wire [4-1:0] node29763;
	wire [4-1:0] node29764;
	wire [4-1:0] node29767;
	wire [4-1:0] node29768;
	wire [4-1:0] node29772;
	wire [4-1:0] node29773;
	wire [4-1:0] node29775;
	wire [4-1:0] node29776;
	wire [4-1:0] node29780;
	wire [4-1:0] node29781;
	wire [4-1:0] node29784;
	wire [4-1:0] node29787;
	wire [4-1:0] node29788;
	wire [4-1:0] node29789;
	wire [4-1:0] node29790;
	wire [4-1:0] node29791;
	wire [4-1:0] node29792;
	wire [4-1:0] node29797;
	wire [4-1:0] node29798;
	wire [4-1:0] node29799;
	wire [4-1:0] node29800;
	wire [4-1:0] node29803;
	wire [4-1:0] node29807;
	wire [4-1:0] node29808;
	wire [4-1:0] node29809;
	wire [4-1:0] node29812;
	wire [4-1:0] node29816;
	wire [4-1:0] node29817;
	wire [4-1:0] node29818;
	wire [4-1:0] node29819;
	wire [4-1:0] node29822;
	wire [4-1:0] node29825;
	wire [4-1:0] node29827;
	wire [4-1:0] node29830;
	wire [4-1:0] node29832;
	wire [4-1:0] node29833;
	wire [4-1:0] node29836;
	wire [4-1:0] node29839;
	wire [4-1:0] node29840;
	wire [4-1:0] node29841;
	wire [4-1:0] node29842;
	wire [4-1:0] node29845;
	wire [4-1:0] node29847;
	wire [4-1:0] node29850;
	wire [4-1:0] node29851;
	wire [4-1:0] node29852;
	wire [4-1:0] node29853;
	wire [4-1:0] node29857;
	wire [4-1:0] node29858;
	wire [4-1:0] node29863;
	wire [4-1:0] node29864;
	wire [4-1:0] node29865;
	wire [4-1:0] node29866;
	wire [4-1:0] node29867;
	wire [4-1:0] node29870;
	wire [4-1:0] node29875;
	wire [4-1:0] node29877;
	wire [4-1:0] node29880;
	wire [4-1:0] node29881;
	wire [4-1:0] node29882;
	wire [4-1:0] node29883;
	wire [4-1:0] node29885;
	wire [4-1:0] node29888;
	wire [4-1:0] node29889;
	wire [4-1:0] node29891;
	wire [4-1:0] node29894;
	wire [4-1:0] node29897;
	wire [4-1:0] node29898;
	wire [4-1:0] node29899;
	wire [4-1:0] node29900;
	wire [4-1:0] node29904;
	wire [4-1:0] node29905;
	wire [4-1:0] node29909;
	wire [4-1:0] node29910;
	wire [4-1:0] node29911;
	wire [4-1:0] node29915;
	wire [4-1:0] node29916;
	wire [4-1:0] node29920;
	wire [4-1:0] node29921;
	wire [4-1:0] node29922;
	wire [4-1:0] node29924;
	wire [4-1:0] node29925;
	wire [4-1:0] node29927;
	wire [4-1:0] node29930;
	wire [4-1:0] node29931;
	wire [4-1:0] node29935;
	wire [4-1:0] node29936;
	wire [4-1:0] node29937;
	wire [4-1:0] node29938;
	wire [4-1:0] node29941;
	wire [4-1:0] node29945;
	wire [4-1:0] node29946;
	wire [4-1:0] node29949;
	wire [4-1:0] node29952;
	wire [4-1:0] node29953;
	wire [4-1:0] node29954;
	wire [4-1:0] node29955;
	wire [4-1:0] node29956;
	wire [4-1:0] node29957;
	wire [4-1:0] node29960;
	wire [4-1:0] node29963;
	wire [4-1:0] node29965;
	wire [4-1:0] node29968;
	wire [4-1:0] node29969;
	wire [4-1:0] node29972;
	wire [4-1:0] node29975;
	wire [4-1:0] node29976;
	wire [4-1:0] node29977;
	wire [4-1:0] node29981;
	wire [4-1:0] node29982;
	wire [4-1:0] node29983;
	wire [4-1:0] node29987;
	wire [4-1:0] node29990;
	wire [4-1:0] node29991;
	wire [4-1:0] node29992;
	wire [4-1:0] node29994;
	wire [4-1:0] node29998;
	wire [4-1:0] node29999;
	wire [4-1:0] node30001;
	wire [4-1:0] node30005;
	wire [4-1:0] node30006;
	wire [4-1:0] node30007;
	wire [4-1:0] node30008;
	wire [4-1:0] node30009;
	wire [4-1:0] node30013;
	wire [4-1:0] node30014;
	wire [4-1:0] node30019;
	wire [4-1:0] node30020;
	wire [4-1:0] node30021;
	wire [4-1:0] node30022;
	wire [4-1:0] node30026;
	wire [4-1:0] node30027;
	wire [4-1:0] node30032;
	wire [4-1:0] node30033;
	wire [4-1:0] node30034;
	wire [4-1:0] node30035;
	wire [4-1:0] node30036;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30039;
	wire [4-1:0] node30040;
	wire [4-1:0] node30041;
	wire [4-1:0] node30042;
	wire [4-1:0] node30044;
	wire [4-1:0] node30047;
	wire [4-1:0] node30049;
	wire [4-1:0] node30052;
	wire [4-1:0] node30053;
	wire [4-1:0] node30055;
	wire [4-1:0] node30058;
	wire [4-1:0] node30060;
	wire [4-1:0] node30063;
	wire [4-1:0] node30064;
	wire [4-1:0] node30065;
	wire [4-1:0] node30067;
	wire [4-1:0] node30070;
	wire [4-1:0] node30072;
	wire [4-1:0] node30075;
	wire [4-1:0] node30076;
	wire [4-1:0] node30078;
	wire [4-1:0] node30081;
	wire [4-1:0] node30083;
	wire [4-1:0] node30086;
	wire [4-1:0] node30087;
	wire [4-1:0] node30088;
	wire [4-1:0] node30089;
	wire [4-1:0] node30091;
	wire [4-1:0] node30094;
	wire [4-1:0] node30096;
	wire [4-1:0] node30099;
	wire [4-1:0] node30101;
	wire [4-1:0] node30102;
	wire [4-1:0] node30105;
	wire [4-1:0] node30108;
	wire [4-1:0] node30109;
	wire [4-1:0] node30110;
	wire [4-1:0] node30112;
	wire [4-1:0] node30115;
	wire [4-1:0] node30116;
	wire [4-1:0] node30117;
	wire [4-1:0] node30118;
	wire [4-1:0] node30122;
	wire [4-1:0] node30123;
	wire [4-1:0] node30127;
	wire [4-1:0] node30129;
	wire [4-1:0] node30132;
	wire [4-1:0] node30133;
	wire [4-1:0] node30134;
	wire [4-1:0] node30135;
	wire [4-1:0] node30137;
	wire [4-1:0] node30141;
	wire [4-1:0] node30143;
	wire [4-1:0] node30146;
	wire [4-1:0] node30147;
	wire [4-1:0] node30148;
	wire [4-1:0] node30150;
	wire [4-1:0] node30153;
	wire [4-1:0] node30154;
	wire [4-1:0] node30159;
	wire [4-1:0] node30160;
	wire [4-1:0] node30161;
	wire [4-1:0] node30162;
	wire [4-1:0] node30164;
	wire [4-1:0] node30165;
	wire [4-1:0] node30166;
	wire [4-1:0] node30170;
	wire [4-1:0] node30171;
	wire [4-1:0] node30175;
	wire [4-1:0] node30176;
	wire [4-1:0] node30178;
	wire [4-1:0] node30181;
	wire [4-1:0] node30183;
	wire [4-1:0] node30184;
	wire [4-1:0] node30187;
	wire [4-1:0] node30190;
	wire [4-1:0] node30191;
	wire [4-1:0] node30192;
	wire [4-1:0] node30195;
	wire [4-1:0] node30198;
	wire [4-1:0] node30199;
	wire [4-1:0] node30201;
	wire [4-1:0] node30203;
	wire [4-1:0] node30204;
	wire [4-1:0] node30207;
	wire [4-1:0] node30210;
	wire [4-1:0] node30211;
	wire [4-1:0] node30212;
	wire [4-1:0] node30215;
	wire [4-1:0] node30219;
	wire [4-1:0] node30220;
	wire [4-1:0] node30221;
	wire [4-1:0] node30222;
	wire [4-1:0] node30225;
	wire [4-1:0] node30228;
	wire [4-1:0] node30229;
	wire [4-1:0] node30231;
	wire [4-1:0] node30234;
	wire [4-1:0] node30236;
	wire [4-1:0] node30239;
	wire [4-1:0] node30240;
	wire [4-1:0] node30241;
	wire [4-1:0] node30243;
	wire [4-1:0] node30246;
	wire [4-1:0] node30248;
	wire [4-1:0] node30251;
	wire [4-1:0] node30252;
	wire [4-1:0] node30254;
	wire [4-1:0] node30257;
	wire [4-1:0] node30260;
	wire [4-1:0] node30261;
	wire [4-1:0] node30262;
	wire [4-1:0] node30263;
	wire [4-1:0] node30264;
	wire [4-1:0] node30265;
	wire [4-1:0] node30268;
	wire [4-1:0] node30271;
	wire [4-1:0] node30272;
	wire [4-1:0] node30275;
	wire [4-1:0] node30278;
	wire [4-1:0] node30279;
	wire [4-1:0] node30280;
	wire [4-1:0] node30281;
	wire [4-1:0] node30282;
	wire [4-1:0] node30283;
	wire [4-1:0] node30286;
	wire [4-1:0] node30290;
	wire [4-1:0] node30291;
	wire [4-1:0] node30295;
	wire [4-1:0] node30296;
	wire [4-1:0] node30298;
	wire [4-1:0] node30301;
	wire [4-1:0] node30303;
	wire [4-1:0] node30304;
	wire [4-1:0] node30308;
	wire [4-1:0] node30309;
	wire [4-1:0] node30310;
	wire [4-1:0] node30313;
	wire [4-1:0] node30314;
	wire [4-1:0] node30317;
	wire [4-1:0] node30320;
	wire [4-1:0] node30321;
	wire [4-1:0] node30322;
	wire [4-1:0] node30325;
	wire [4-1:0] node30328;
	wire [4-1:0] node30330;
	wire [4-1:0] node30333;
	wire [4-1:0] node30334;
	wire [4-1:0] node30335;
	wire [4-1:0] node30336;
	wire [4-1:0] node30337;
	wire [4-1:0] node30340;
	wire [4-1:0] node30343;
	wire [4-1:0] node30345;
	wire [4-1:0] node30346;
	wire [4-1:0] node30349;
	wire [4-1:0] node30352;
	wire [4-1:0] node30353;
	wire [4-1:0] node30354;
	wire [4-1:0] node30356;
	wire [4-1:0] node30357;
	wire [4-1:0] node30360;
	wire [4-1:0] node30364;
	wire [4-1:0] node30366;
	wire [4-1:0] node30368;
	wire [4-1:0] node30369;
	wire [4-1:0] node30373;
	wire [4-1:0] node30374;
	wire [4-1:0] node30375;
	wire [4-1:0] node30376;
	wire [4-1:0] node30379;
	wire [4-1:0] node30382;
	wire [4-1:0] node30383;
	wire [4-1:0] node30384;
	wire [4-1:0] node30387;
	wire [4-1:0] node30391;
	wire [4-1:0] node30392;
	wire [4-1:0] node30395;
	wire [4-1:0] node30396;
	wire [4-1:0] node30398;
	wire [4-1:0] node30401;
	wire [4-1:0] node30403;
	wire [4-1:0] node30406;
	wire [4-1:0] node30407;
	wire [4-1:0] node30408;
	wire [4-1:0] node30409;
	wire [4-1:0] node30410;
	wire [4-1:0] node30411;
	wire [4-1:0] node30412;
	wire [4-1:0] node30415;
	wire [4-1:0] node30418;
	wire [4-1:0] node30419;
	wire [4-1:0] node30422;
	wire [4-1:0] node30425;
	wire [4-1:0] node30427;
	wire [4-1:0] node30428;
	wire [4-1:0] node30432;
	wire [4-1:0] node30433;
	wire [4-1:0] node30434;
	wire [4-1:0] node30436;
	wire [4-1:0] node30438;
	wire [4-1:0] node30442;
	wire [4-1:0] node30443;
	wire [4-1:0] node30444;
	wire [4-1:0] node30446;
	wire [4-1:0] node30449;
	wire [4-1:0] node30453;
	wire [4-1:0] node30454;
	wire [4-1:0] node30455;
	wire [4-1:0] node30456;
	wire [4-1:0] node30459;
	wire [4-1:0] node30462;
	wire [4-1:0] node30463;
	wire [4-1:0] node30467;
	wire [4-1:0] node30468;
	wire [4-1:0] node30469;
	wire [4-1:0] node30472;
	wire [4-1:0] node30475;
	wire [4-1:0] node30476;
	wire [4-1:0] node30477;
	wire [4-1:0] node30481;
	wire [4-1:0] node30483;
	wire [4-1:0] node30484;
	wire [4-1:0] node30487;
	wire [4-1:0] node30490;
	wire [4-1:0] node30491;
	wire [4-1:0] node30492;
	wire [4-1:0] node30493;
	wire [4-1:0] node30494;
	wire [4-1:0] node30498;
	wire [4-1:0] node30499;
	wire [4-1:0] node30503;
	wire [4-1:0] node30504;
	wire [4-1:0] node30505;
	wire [4-1:0] node30509;
	wire [4-1:0] node30510;
	wire [4-1:0] node30514;
	wire [4-1:0] node30515;
	wire [4-1:0] node30516;
	wire [4-1:0] node30517;
	wire [4-1:0] node30519;
	wire [4-1:0] node30521;
	wire [4-1:0] node30524;
	wire [4-1:0] node30526;
	wire [4-1:0] node30527;
	wire [4-1:0] node30530;
	wire [4-1:0] node30533;
	wire [4-1:0] node30534;
	wire [4-1:0] node30535;
	wire [4-1:0] node30538;
	wire [4-1:0] node30541;
	wire [4-1:0] node30542;
	wire [4-1:0] node30545;
	wire [4-1:0] node30548;
	wire [4-1:0] node30549;
	wire [4-1:0] node30550;
	wire [4-1:0] node30551;
	wire [4-1:0] node30554;
	wire [4-1:0] node30555;
	wire [4-1:0] node30559;
	wire [4-1:0] node30560;
	wire [4-1:0] node30562;
	wire [4-1:0] node30565;
	wire [4-1:0] node30566;
	wire [4-1:0] node30571;
	wire [4-1:0] node30572;
	wire [4-1:0] node30573;
	wire [4-1:0] node30574;
	wire [4-1:0] node30575;
	wire [4-1:0] node30578;
	wire [4-1:0] node30579;
	wire [4-1:0] node30581;
	wire [4-1:0] node30584;
	wire [4-1:0] node30585;
	wire [4-1:0] node30589;
	wire [4-1:0] node30590;
	wire [4-1:0] node30591;
	wire [4-1:0] node30592;
	wire [4-1:0] node30593;
	wire [4-1:0] node30594;
	wire [4-1:0] node30598;
	wire [4-1:0] node30599;
	wire [4-1:0] node30602;
	wire [4-1:0] node30605;
	wire [4-1:0] node30606;
	wire [4-1:0] node30609;
	wire [4-1:0] node30612;
	wire [4-1:0] node30613;
	wire [4-1:0] node30614;
	wire [4-1:0] node30617;
	wire [4-1:0] node30620;
	wire [4-1:0] node30621;
	wire [4-1:0] node30623;
	wire [4-1:0] node30624;
	wire [4-1:0] node30628;
	wire [4-1:0] node30629;
	wire [4-1:0] node30633;
	wire [4-1:0] node30634;
	wire [4-1:0] node30636;
	wire [4-1:0] node30639;
	wire [4-1:0] node30640;
	wire [4-1:0] node30644;
	wire [4-1:0] node30645;
	wire [4-1:0] node30646;
	wire [4-1:0] node30649;
	wire [4-1:0] node30650;
	wire [4-1:0] node30652;
	wire [4-1:0] node30655;
	wire [4-1:0] node30656;
	wire [4-1:0] node30660;
	wire [4-1:0] node30661;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30664;
	wire [4-1:0] node30665;
	wire [4-1:0] node30668;
	wire [4-1:0] node30672;
	wire [4-1:0] node30673;
	wire [4-1:0] node30676;
	wire [4-1:0] node30679;
	wire [4-1:0] node30680;
	wire [4-1:0] node30681;
	wire [4-1:0] node30682;
	wire [4-1:0] node30683;
	wire [4-1:0] node30686;
	wire [4-1:0] node30691;
	wire [4-1:0] node30693;
	wire [4-1:0] node30694;
	wire [4-1:0] node30697;
	wire [4-1:0] node30700;
	wire [4-1:0] node30701;
	wire [4-1:0] node30702;
	wire [4-1:0] node30706;
	wire [4-1:0] node30707;
	wire [4-1:0] node30711;
	wire [4-1:0] node30712;
	wire [4-1:0] node30713;
	wire [4-1:0] node30714;
	wire [4-1:0] node30717;
	wire [4-1:0] node30718;
	wire [4-1:0] node30720;
	wire [4-1:0] node30723;
	wire [4-1:0] node30724;
	wire [4-1:0] node30728;
	wire [4-1:0] node30729;
	wire [4-1:0] node30730;
	wire [4-1:0] node30731;
	wire [4-1:0] node30734;
	wire [4-1:0] node30737;
	wire [4-1:0] node30738;
	wire [4-1:0] node30739;
	wire [4-1:0] node30742;
	wire [4-1:0] node30745;
	wire [4-1:0] node30746;
	wire [4-1:0] node30748;
	wire [4-1:0] node30749;
	wire [4-1:0] node30753;
	wire [4-1:0] node30754;
	wire [4-1:0] node30755;
	wire [4-1:0] node30758;
	wire [4-1:0] node30762;
	wire [4-1:0] node30763;
	wire [4-1:0] node30764;
	wire [4-1:0] node30768;
	wire [4-1:0] node30769;
	wire [4-1:0] node30773;
	wire [4-1:0] node30774;
	wire [4-1:0] node30775;
	wire [4-1:0] node30778;
	wire [4-1:0] node30779;
	wire [4-1:0] node30781;
	wire [4-1:0] node30784;
	wire [4-1:0] node30785;
	wire [4-1:0] node30789;
	wire [4-1:0] node30790;
	wire [4-1:0] node30791;
	wire [4-1:0] node30792;
	wire [4-1:0] node30793;
	wire [4-1:0] node30796;
	wire [4-1:0] node30799;
	wire [4-1:0] node30800;
	wire [4-1:0] node30804;
	wire [4-1:0] node30805;
	wire [4-1:0] node30806;
	wire [4-1:0] node30810;
	wire [4-1:0] node30813;
	wire [4-1:0] node30814;
	wire [4-1:0] node30815;
	wire [4-1:0] node30816;
	wire [4-1:0] node30817;
	wire [4-1:0] node30822;
	wire [4-1:0] node30823;
	wire [4-1:0] node30824;
	wire [4-1:0] node30827;
	wire [4-1:0] node30829;
	wire [4-1:0] node30832;
	wire [4-1:0] node30834;
	wire [4-1:0] node30837;
	wire [4-1:0] node30838;
	wire [4-1:0] node30840;
	wire [4-1:0] node30843;
	wire [4-1:0] node30844;
	wire [4-1:0] node30848;
	wire [4-1:0] node30849;
	wire [4-1:0] node30850;
	wire [4-1:0] node30851;
	wire [4-1:0] node30852;
	wire [4-1:0] node30853;
	wire [4-1:0] node30854;
	wire [4-1:0] node30855;
	wire [4-1:0] node30856;
	wire [4-1:0] node30858;
	wire [4-1:0] node30861;
	wire [4-1:0] node30864;
	wire [4-1:0] node30865;
	wire [4-1:0] node30868;
	wire [4-1:0] node30871;
	wire [4-1:0] node30872;
	wire [4-1:0] node30874;
	wire [4-1:0] node30875;
	wire [4-1:0] node30878;
	wire [4-1:0] node30881;
	wire [4-1:0] node30882;
	wire [4-1:0] node30885;
	wire [4-1:0] node30888;
	wire [4-1:0] node30889;
	wire [4-1:0] node30890;
	wire [4-1:0] node30893;
	wire [4-1:0] node30896;
	wire [4-1:0] node30897;
	wire [4-1:0] node30899;
	wire [4-1:0] node30900;
	wire [4-1:0] node30904;
	wire [4-1:0] node30907;
	wire [4-1:0] node30908;
	wire [4-1:0] node30909;
	wire [4-1:0] node30910;
	wire [4-1:0] node30911;
	wire [4-1:0] node30914;
	wire [4-1:0] node30917;
	wire [4-1:0] node30920;
	wire [4-1:0] node30921;
	wire [4-1:0] node30922;
	wire [4-1:0] node30925;
	wire [4-1:0] node30928;
	wire [4-1:0] node30929;
	wire [4-1:0] node30930;
	wire [4-1:0] node30932;
	wire [4-1:0] node30936;
	wire [4-1:0] node30937;
	wire [4-1:0] node30940;
	wire [4-1:0] node30943;
	wire [4-1:0] node30944;
	wire [4-1:0] node30945;
	wire [4-1:0] node30946;
	wire [4-1:0] node30949;
	wire [4-1:0] node30952;
	wire [4-1:0] node30953;
	wire [4-1:0] node30954;
	wire [4-1:0] node30957;
	wire [4-1:0] node30961;
	wire [4-1:0] node30962;
	wire [4-1:0] node30963;
	wire [4-1:0] node30966;
	wire [4-1:0] node30969;
	wire [4-1:0] node30971;
	wire [4-1:0] node30972;
	wire [4-1:0] node30975;
	wire [4-1:0] node30978;
	wire [4-1:0] node30979;
	wire [4-1:0] node30980;
	wire [4-1:0] node30981;
	wire [4-1:0] node30982;
	wire [4-1:0] node30983;
	wire [4-1:0] node30984;
	wire [4-1:0] node30986;
	wire [4-1:0] node30990;
	wire [4-1:0] node30991;
	wire [4-1:0] node30995;
	wire [4-1:0] node30996;
	wire [4-1:0] node30997;
	wire [4-1:0] node31001;
	wire [4-1:0] node31004;
	wire [4-1:0] node31005;
	wire [4-1:0] node31006;
	wire [4-1:0] node31010;
	wire [4-1:0] node31012;
	wire [4-1:0] node31014;
	wire [4-1:0] node31017;
	wire [4-1:0] node31018;
	wire [4-1:0] node31019;
	wire [4-1:0] node31020;
	wire [4-1:0] node31021;
	wire [4-1:0] node31026;
	wire [4-1:0] node31027;
	wire [4-1:0] node31031;
	wire [4-1:0] node31032;
	wire [4-1:0] node31034;
	wire [4-1:0] node31036;
	wire [4-1:0] node31039;
	wire [4-1:0] node31040;
	wire [4-1:0] node31041;
	wire [4-1:0] node31044;
	wire [4-1:0] node31046;
	wire [4-1:0] node31050;
	wire [4-1:0] node31051;
	wire [4-1:0] node31052;
	wire [4-1:0] node31054;
	wire [4-1:0] node31057;
	wire [4-1:0] node31058;
	wire [4-1:0] node31062;
	wire [4-1:0] node31065;
	wire [4-1:0] node31066;
	wire [4-1:0] node31067;
	wire [4-1:0] node31068;
	wire [4-1:0] node31069;
	wire [4-1:0] node31070;
	wire [4-1:0] node31071;
	wire [4-1:0] node31072;
	wire [4-1:0] node31075;
	wire [4-1:0] node31078;
	wire [4-1:0] node31080;
	wire [4-1:0] node31083;
	wire [4-1:0] node31085;
	wire [4-1:0] node31087;
	wire [4-1:0] node31090;
	wire [4-1:0] node31091;
	wire [4-1:0] node31092;
	wire [4-1:0] node31094;
	wire [4-1:0] node31098;
	wire [4-1:0] node31099;
	wire [4-1:0] node31100;
	wire [4-1:0] node31105;
	wire [4-1:0] node31106;
	wire [4-1:0] node31107;
	wire [4-1:0] node31109;
	wire [4-1:0] node31110;
	wire [4-1:0] node31113;
	wire [4-1:0] node31116;
	wire [4-1:0] node31117;
	wire [4-1:0] node31118;
	wire [4-1:0] node31119;
	wire [4-1:0] node31123;
	wire [4-1:0] node31125;
	wire [4-1:0] node31129;
	wire [4-1:0] node31130;
	wire [4-1:0] node31131;
	wire [4-1:0] node31134;
	wire [4-1:0] node31135;
	wire [4-1:0] node31139;
	wire [4-1:0] node31140;
	wire [4-1:0] node31141;
	wire [4-1:0] node31146;
	wire [4-1:0] node31147;
	wire [4-1:0] node31148;
	wire [4-1:0] node31149;
	wire [4-1:0] node31152;
	wire [4-1:0] node31153;
	wire [4-1:0] node31154;
	wire [4-1:0] node31157;
	wire [4-1:0] node31160;
	wire [4-1:0] node31163;
	wire [4-1:0] node31164;
	wire [4-1:0] node31165;
	wire [4-1:0] node31168;
	wire [4-1:0] node31170;
	wire [4-1:0] node31173;
	wire [4-1:0] node31174;
	wire [4-1:0] node31175;
	wire [4-1:0] node31180;
	wire [4-1:0] node31181;
	wire [4-1:0] node31182;
	wire [4-1:0] node31183;
	wire [4-1:0] node31185;
	wire [4-1:0] node31188;
	wire [4-1:0] node31189;
	wire [4-1:0] node31193;
	wire [4-1:0] node31195;
	wire [4-1:0] node31198;
	wire [4-1:0] node31199;
	wire [4-1:0] node31200;
	wire [4-1:0] node31201;
	wire [4-1:0] node31204;
	wire [4-1:0] node31207;
	wire [4-1:0] node31208;
	wire [4-1:0] node31211;
	wire [4-1:0] node31214;
	wire [4-1:0] node31215;
	wire [4-1:0] node31218;
	wire [4-1:0] node31220;
	wire [4-1:0] node31223;
	wire [4-1:0] node31224;
	wire [4-1:0] node31225;
	wire [4-1:0] node31226;
	wire [4-1:0] node31227;
	wire [4-1:0] node31231;
	wire [4-1:0] node31233;
	wire [4-1:0] node31236;
	wire [4-1:0] node31237;
	wire [4-1:0] node31238;
	wire [4-1:0] node31241;
	wire [4-1:0] node31244;
	wire [4-1:0] node31245;
	wire [4-1:0] node31246;
	wire [4-1:0] node31249;
	wire [4-1:0] node31252;
	wire [4-1:0] node31253;
	wire [4-1:0] node31256;
	wire [4-1:0] node31259;
	wire [4-1:0] node31260;
	wire [4-1:0] node31261;
	wire [4-1:0] node31263;
	wire [4-1:0] node31266;
	wire [4-1:0] node31267;
	wire [4-1:0] node31271;
	wire [4-1:0] node31274;
	wire [4-1:0] node31275;
	wire [4-1:0] node31276;
	wire [4-1:0] node31277;
	wire [4-1:0] node31278;
	wire [4-1:0] node31279;
	wire [4-1:0] node31281;
	wire [4-1:0] node31284;
	wire [4-1:0] node31285;
	wire [4-1:0] node31286;
	wire [4-1:0] node31290;
	wire [4-1:0] node31291;
	wire [4-1:0] node31294;
	wire [4-1:0] node31297;
	wire [4-1:0] node31298;
	wire [4-1:0] node31299;
	wire [4-1:0] node31301;
	wire [4-1:0] node31305;
	wire [4-1:0] node31306;
	wire [4-1:0] node31309;
	wire [4-1:0] node31312;
	wire [4-1:0] node31313;
	wire [4-1:0] node31314;
	wire [4-1:0] node31316;
	wire [4-1:0] node31319;
	wire [4-1:0] node31321;
	wire [4-1:0] node31322;
	wire [4-1:0] node31326;
	wire [4-1:0] node31327;
	wire [4-1:0] node31328;
	wire [4-1:0] node31329;
	wire [4-1:0] node31333;
	wire [4-1:0] node31335;
	wire [4-1:0] node31336;
	wire [4-1:0] node31339;
	wire [4-1:0] node31342;
	wire [4-1:0] node31343;
	wire [4-1:0] node31347;
	wire [4-1:0] node31348;
	wire [4-1:0] node31349;
	wire [4-1:0] node31350;
	wire [4-1:0] node31351;
	wire [4-1:0] node31355;
	wire [4-1:0] node31356;
	wire [4-1:0] node31360;
	wire [4-1:0] node31361;
	wire [4-1:0] node31362;
	wire [4-1:0] node31365;
	wire [4-1:0] node31368;
	wire [4-1:0] node31369;
	wire [4-1:0] node31370;
	wire [4-1:0] node31374;
	wire [4-1:0] node31375;
	wire [4-1:0] node31378;
	wire [4-1:0] node31381;
	wire [4-1:0] node31382;
	wire [4-1:0] node31383;
	wire [4-1:0] node31385;
	wire [4-1:0] node31388;
	wire [4-1:0] node31389;
	wire [4-1:0] node31393;
	wire [4-1:0] node31396;
	wire [4-1:0] node31397;
	wire [4-1:0] node31398;
	wire [4-1:0] node31399;
	wire [4-1:0] node31400;
	wire [4-1:0] node31403;
	wire [4-1:0] node31404;
	wire [4-1:0] node31406;
	wire [4-1:0] node31407;
	wire [4-1:0] node31410;
	wire [4-1:0] node31412;
	wire [4-1:0] node31415;
	wire [4-1:0] node31418;
	wire [4-1:0] node31419;
	wire [4-1:0] node31420;
	wire [4-1:0] node31423;
	wire [4-1:0] node31425;
	wire [4-1:0] node31428;
	wire [4-1:0] node31429;
	wire [4-1:0] node31430;
	wire [4-1:0] node31434;
	wire [4-1:0] node31437;
	wire [4-1:0] node31438;
	wire [4-1:0] node31439;
	wire [4-1:0] node31441;
	wire [4-1:0] node31444;
	wire [4-1:0] node31445;
	wire [4-1:0] node31446;
	wire [4-1:0] node31450;
	wire [4-1:0] node31452;
	wire [4-1:0] node31453;
	wire [4-1:0] node31456;
	wire [4-1:0] node31459;
	wire [4-1:0] node31460;
	wire [4-1:0] node31461;
	wire [4-1:0] node31463;
	wire [4-1:0] node31467;
	wire [4-1:0] node31468;
	wire [4-1:0] node31472;
	wire [4-1:0] node31473;
	wire [4-1:0] node31474;
	wire [4-1:0] node31475;
	wire [4-1:0] node31476;
	wire [4-1:0] node31480;
	wire [4-1:0] node31482;
	wire [4-1:0] node31485;
	wire [4-1:0] node31486;
	wire [4-1:0] node31487;
	wire [4-1:0] node31488;
	wire [4-1:0] node31491;
	wire [4-1:0] node31494;
	wire [4-1:0] node31495;
	wire [4-1:0] node31498;
	wire [4-1:0] node31501;
	wire [4-1:0] node31502;
	wire [4-1:0] node31503;
	wire [4-1:0] node31506;
	wire [4-1:0] node31509;
	wire [4-1:0] node31510;
	wire [4-1:0] node31514;
	wire [4-1:0] node31515;
	wire [4-1:0] node31516;
	wire [4-1:0] node31518;
	wire [4-1:0] node31521;
	wire [4-1:0] node31522;
	wire [4-1:0] node31526;
	wire [4-1:0] node31529;
	wire [4-1:0] node31530;
	wire [4-1:0] node31531;
	wire [4-1:0] node31532;
	wire [4-1:0] node31533;
	wire [4-1:0] node31534;
	wire [4-1:0] node31535;
	wire [4-1:0] node31536;
	wire [4-1:0] node31537;
	wire [4-1:0] node31538;
	wire [4-1:0] node31541;
	wire [4-1:0] node31543;
	wire [4-1:0] node31545;
	wire [4-1:0] node31548;
	wire [4-1:0] node31549;
	wire [4-1:0] node31552;
	wire [4-1:0] node31555;
	wire [4-1:0] node31556;
	wire [4-1:0] node31557;
	wire [4-1:0] node31558;
	wire [4-1:0] node31561;
	wire [4-1:0] node31564;
	wire [4-1:0] node31566;
	wire [4-1:0] node31569;
	wire [4-1:0] node31570;
	wire [4-1:0] node31573;
	wire [4-1:0] node31574;
	wire [4-1:0] node31575;
	wire [4-1:0] node31578;
	wire [4-1:0] node31581;
	wire [4-1:0] node31584;
	wire [4-1:0] node31585;
	wire [4-1:0] node31586;
	wire [4-1:0] node31588;
	wire [4-1:0] node31589;
	wire [4-1:0] node31592;
	wire [4-1:0] node31595;
	wire [4-1:0] node31596;
	wire [4-1:0] node31597;
	wire [4-1:0] node31600;
	wire [4-1:0] node31603;
	wire [4-1:0] node31606;
	wire [4-1:0] node31607;
	wire [4-1:0] node31608;
	wire [4-1:0] node31609;
	wire [4-1:0] node31612;
	wire [4-1:0] node31615;
	wire [4-1:0] node31617;
	wire [4-1:0] node31620;
	wire [4-1:0] node31621;
	wire [4-1:0] node31622;
	wire [4-1:0] node31625;
	wire [4-1:0] node31629;
	wire [4-1:0] node31630;
	wire [4-1:0] node31631;
	wire [4-1:0] node31632;
	wire [4-1:0] node31633;
	wire [4-1:0] node31636;
	wire [4-1:0] node31637;
	wire [4-1:0] node31638;
	wire [4-1:0] node31642;
	wire [4-1:0] node31645;
	wire [4-1:0] node31646;
	wire [4-1:0] node31647;
	wire [4-1:0] node31648;
	wire [4-1:0] node31651;
	wire [4-1:0] node31654;
	wire [4-1:0] node31657;
	wire [4-1:0] node31658;
	wire [4-1:0] node31661;
	wire [4-1:0] node31664;
	wire [4-1:0] node31665;
	wire [4-1:0] node31666;
	wire [4-1:0] node31667;
	wire [4-1:0] node31671;
	wire [4-1:0] node31672;
	wire [4-1:0] node31673;
	wire [4-1:0] node31676;
	wire [4-1:0] node31680;
	wire [4-1:0] node31682;
	wire [4-1:0] node31683;
	wire [4-1:0] node31684;
	wire [4-1:0] node31687;
	wire [4-1:0] node31690;
	wire [4-1:0] node31692;
	wire [4-1:0] node31695;
	wire [4-1:0] node31696;
	wire [4-1:0] node31697;
	wire [4-1:0] node31698;
	wire [4-1:0] node31700;
	wire [4-1:0] node31703;
	wire [4-1:0] node31704;
	wire [4-1:0] node31708;
	wire [4-1:0] node31710;
	wire [4-1:0] node31712;
	wire [4-1:0] node31714;
	wire [4-1:0] node31717;
	wire [4-1:0] node31718;
	wire [4-1:0] node31719;
	wire [4-1:0] node31722;
	wire [4-1:0] node31725;
	wire [4-1:0] node31726;
	wire [4-1:0] node31727;
	wire [4-1:0] node31730;
	wire [4-1:0] node31733;
	wire [4-1:0] node31736;
	wire [4-1:0] node31737;
	wire [4-1:0] node31738;
	wire [4-1:0] node31739;
	wire [4-1:0] node31740;
	wire [4-1:0] node31741;
	wire [4-1:0] node31743;
	wire [4-1:0] node31747;
	wire [4-1:0] node31748;
	wire [4-1:0] node31752;
	wire [4-1:0] node31753;
	wire [4-1:0] node31754;
	wire [4-1:0] node31755;
	wire [4-1:0] node31756;
	wire [4-1:0] node31759;
	wire [4-1:0] node31764;
	wire [4-1:0] node31766;
	wire [4-1:0] node31767;
	wire [4-1:0] node31768;
	wire [4-1:0] node31773;
	wire [4-1:0] node31774;
	wire [4-1:0] node31775;
	wire [4-1:0] node31776;
	wire [4-1:0] node31778;
	wire [4-1:0] node31781;
	wire [4-1:0] node31782;
	wire [4-1:0] node31785;
	wire [4-1:0] node31788;
	wire [4-1:0] node31789;
	wire [4-1:0] node31792;
	wire [4-1:0] node31793;
	wire [4-1:0] node31797;
	wire [4-1:0] node31798;
	wire [4-1:0] node31799;
	wire [4-1:0] node31800;
	wire [4-1:0] node31803;
	wire [4-1:0] node31804;
	wire [4-1:0] node31807;
	wire [4-1:0] node31811;
	wire [4-1:0] node31812;
	wire [4-1:0] node31814;
	wire [4-1:0] node31816;
	wire [4-1:0] node31820;
	wire [4-1:0] node31821;
	wire [4-1:0] node31822;
	wire [4-1:0] node31823;
	wire [4-1:0] node31825;
	wire [4-1:0] node31826;
	wire [4-1:0] node31829;
	wire [4-1:0] node31832;
	wire [4-1:0] node31833;
	wire [4-1:0] node31835;
	wire [4-1:0] node31836;
	wire [4-1:0] node31839;
	wire [4-1:0] node31843;
	wire [4-1:0] node31844;
	wire [4-1:0] node31846;
	wire [4-1:0] node31847;
	wire [4-1:0] node31851;
	wire [4-1:0] node31852;
	wire [4-1:0] node31853;
	wire [4-1:0] node31857;
	wire [4-1:0] node31860;
	wire [4-1:0] node31861;
	wire [4-1:0] node31862;
	wire [4-1:0] node31864;
	wire [4-1:0] node31867;
	wire [4-1:0] node31868;
	wire [4-1:0] node31869;
	wire [4-1:0] node31873;
	wire [4-1:0] node31875;
	wire [4-1:0] node31877;
	wire [4-1:0] node31880;
	wire [4-1:0] node31881;
	wire [4-1:0] node31882;
	wire [4-1:0] node31883;
	wire [4-1:0] node31888;
	wire [4-1:0] node31890;
	wire [4-1:0] node31893;
	wire [4-1:0] node31894;
	wire [4-1:0] node31895;
	wire [4-1:0] node31896;
	wire [4-1:0] node31897;
	wire [4-1:0] node31898;
	wire [4-1:0] node31899;
	wire [4-1:0] node31902;
	wire [4-1:0] node31905;
	wire [4-1:0] node31906;
	wire [4-1:0] node31909;
	wire [4-1:0] node31912;
	wire [4-1:0] node31913;
	wire [4-1:0] node31914;
	wire [4-1:0] node31917;
	wire [4-1:0] node31920;
	wire [4-1:0] node31921;
	wire [4-1:0] node31923;
	wire [4-1:0] node31924;
	wire [4-1:0] node31928;
	wire [4-1:0] node31929;
	wire [4-1:0] node31930;
	wire [4-1:0] node31934;
	wire [4-1:0] node31935;
	wire [4-1:0] node31939;
	wire [4-1:0] node31940;
	wire [4-1:0] node31941;
	wire [4-1:0] node31942;
	wire [4-1:0] node31945;
	wire [4-1:0] node31948;
	wire [4-1:0] node31951;
	wire [4-1:0] node31952;
	wire [4-1:0] node31953;
	wire [4-1:0] node31956;
	wire [4-1:0] node31959;
	wire [4-1:0] node31960;
	wire [4-1:0] node31962;
	wire [4-1:0] node31966;
	wire [4-1:0] node31967;
	wire [4-1:0] node31968;
	wire [4-1:0] node31969;
	wire [4-1:0] node31971;
	wire [4-1:0] node31973;
	wire [4-1:0] node31976;
	wire [4-1:0] node31977;
	wire [4-1:0] node31978;
	wire [4-1:0] node31982;
	wire [4-1:0] node31983;
	wire [4-1:0] node31987;
	wire [4-1:0] node31988;
	wire [4-1:0] node31991;
	wire [4-1:0] node31993;
	wire [4-1:0] node31995;
	wire [4-1:0] node31997;
	wire [4-1:0] node32000;
	wire [4-1:0] node32001;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32005;
	wire [4-1:0] node32009;
	wire [4-1:0] node32010;
	wire [4-1:0] node32012;
	wire [4-1:0] node32015;
	wire [4-1:0] node32018;
	wire [4-1:0] node32019;
	wire [4-1:0] node32020;
	wire [4-1:0] node32021;
	wire [4-1:0] node32024;
	wire [4-1:0] node32025;
	wire [4-1:0] node32029;
	wire [4-1:0] node32031;
	wire [4-1:0] node32034;
	wire [4-1:0] node32035;
	wire [4-1:0] node32036;
	wire [4-1:0] node32039;
	wire [4-1:0] node32043;
	wire [4-1:0] node32044;
	wire [4-1:0] node32045;
	wire [4-1:0] node32046;
	wire [4-1:0] node32047;
	wire [4-1:0] node32050;
	wire [4-1:0] node32053;
	wire [4-1:0] node32054;
	wire [4-1:0] node32056;
	wire [4-1:0] node32059;
	wire [4-1:0] node32062;
	wire [4-1:0] node32063;
	wire [4-1:0] node32064;
	wire [4-1:0] node32065;
	wire [4-1:0] node32066;
	wire [4-1:0] node32070;
	wire [4-1:0] node32072;
	wire [4-1:0] node32075;
	wire [4-1:0] node32076;
	wire [4-1:0] node32079;
	wire [4-1:0] node32082;
	wire [4-1:0] node32083;
	wire [4-1:0] node32084;
	wire [4-1:0] node32085;
	wire [4-1:0] node32089;
	wire [4-1:0] node32090;
	wire [4-1:0] node32091;
	wire [4-1:0] node32095;
	wire [4-1:0] node32096;
	wire [4-1:0] node32099;
	wire [4-1:0] node32102;
	wire [4-1:0] node32103;
	wire [4-1:0] node32104;
	wire [4-1:0] node32108;
	wire [4-1:0] node32109;
	wire [4-1:0] node32112;
	wire [4-1:0] node32115;
	wire [4-1:0] node32116;
	wire [4-1:0] node32117;
	wire [4-1:0] node32118;
	wire [4-1:0] node32121;
	wire [4-1:0] node32122;
	wire [4-1:0] node32125;
	wire [4-1:0] node32128;
	wire [4-1:0] node32129;
	wire [4-1:0] node32130;
	wire [4-1:0] node32131;
	wire [4-1:0] node32136;
	wire [4-1:0] node32137;
	wire [4-1:0] node32140;
	wire [4-1:0] node32143;
	wire [4-1:0] node32144;
	wire [4-1:0] node32145;
	wire [4-1:0] node32147;
	wire [4-1:0] node32149;
	wire [4-1:0] node32153;
	wire [4-1:0] node32154;
	wire [4-1:0] node32155;
	wire [4-1:0] node32156;
	wire [4-1:0] node32160;
	wire [4-1:0] node32163;
	wire [4-1:0] node32164;
	wire [4-1:0] node32167;
	wire [4-1:0] node32170;
	wire [4-1:0] node32171;
	wire [4-1:0] node32172;
	wire [4-1:0] node32173;
	wire [4-1:0] node32174;
	wire [4-1:0] node32175;
	wire [4-1:0] node32177;
	wire [4-1:0] node32180;
	wire [4-1:0] node32182;
	wire [4-1:0] node32185;
	wire [4-1:0] node32186;
	wire [4-1:0] node32188;
	wire [4-1:0] node32191;
	wire [4-1:0] node32193;
	wire [4-1:0] node32196;
	wire [4-1:0] node32197;
	wire [4-1:0] node32198;
	wire [4-1:0] node32201;
	wire [4-1:0] node32204;
	wire [4-1:0] node32205;
	wire [4-1:0] node32208;
	wire [4-1:0] node32211;
	wire [4-1:0] node32212;
	wire [4-1:0] node32213;
	wire [4-1:0] node32214;
	wire [4-1:0] node32216;
	wire [4-1:0] node32219;
	wire [4-1:0] node32220;
	wire [4-1:0] node32224;
	wire [4-1:0] node32225;
	wire [4-1:0] node32226;
	wire [4-1:0] node32230;
	wire [4-1:0] node32231;
	wire [4-1:0] node32235;
	wire [4-1:0] node32236;
	wire [4-1:0] node32237;
	wire [4-1:0] node32238;
	wire [4-1:0] node32239;
	wire [4-1:0] node32242;
	wire [4-1:0] node32245;
	wire [4-1:0] node32247;
	wire [4-1:0] node32248;
	wire [4-1:0] node32249;
	wire [4-1:0] node32252;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32259;
	wire [4-1:0] node32261;
	wire [4-1:0] node32264;
	wire [4-1:0] node32265;
	wire [4-1:0] node32268;
	wire [4-1:0] node32271;
	wire [4-1:0] node32272;
	wire [4-1:0] node32275;
	wire [4-1:0] node32278;
	wire [4-1:0] node32279;
	wire [4-1:0] node32280;
	wire [4-1:0] node32281;
	wire [4-1:0] node32282;
	wire [4-1:0] node32283;
	wire [4-1:0] node32284;
	wire [4-1:0] node32285;
	wire [4-1:0] node32289;
	wire [4-1:0] node32292;
	wire [4-1:0] node32293;
	wire [4-1:0] node32297;
	wire [4-1:0] node32298;
	wire [4-1:0] node32299;
	wire [4-1:0] node32302;
	wire [4-1:0] node32305;
	wire [4-1:0] node32307;
	wire [4-1:0] node32310;
	wire [4-1:0] node32311;
	wire [4-1:0] node32312;
	wire [4-1:0] node32313;
	wire [4-1:0] node32314;
	wire [4-1:0] node32315;
	wire [4-1:0] node32318;
	wire [4-1:0] node32321;
	wire [4-1:0] node32322;
	wire [4-1:0] node32326;
	wire [4-1:0] node32327;
	wire [4-1:0] node32330;
	wire [4-1:0] node32333;
	wire [4-1:0] node32335;
	wire [4-1:0] node32336;
	wire [4-1:0] node32340;
	wire [4-1:0] node32341;
	wire [4-1:0] node32342;
	wire [4-1:0] node32344;
	wire [4-1:0] node32348;
	wire [4-1:0] node32349;
	wire [4-1:0] node32350;
	wire [4-1:0] node32353;
	wire [4-1:0] node32356;
	wire [4-1:0] node32359;
	wire [4-1:0] node32360;
	wire [4-1:0] node32361;
	wire [4-1:0] node32362;
	wire [4-1:0] node32363;
	wire [4-1:0] node32364;
	wire [4-1:0] node32368;
	wire [4-1:0] node32371;
	wire [4-1:0] node32372;
	wire [4-1:0] node32376;
	wire [4-1:0] node32377;
	wire [4-1:0] node32378;
	wire [4-1:0] node32382;
	wire [4-1:0] node32383;
	wire [4-1:0] node32384;
	wire [4-1:0] node32385;
	wire [4-1:0] node32389;
	wire [4-1:0] node32391;
	wire [4-1:0] node32394;
	wire [4-1:0] node32396;
	wire [4-1:0] node32399;
	wire [4-1:0] node32400;
	wire [4-1:0] node32401;
	wire [4-1:0] node32405;
	wire [4-1:0] node32406;
	wire [4-1:0] node32409;
	wire [4-1:0] node32412;
	wire [4-1:0] node32413;
	wire [4-1:0] node32414;
	wire [4-1:0] node32415;
	wire [4-1:0] node32416;
	wire [4-1:0] node32417;
	wire [4-1:0] node32421;
	wire [4-1:0] node32422;
	wire [4-1:0] node32425;
	wire [4-1:0] node32428;
	wire [4-1:0] node32429;
	wire [4-1:0] node32431;
	wire [4-1:0] node32434;
	wire [4-1:0] node32435;
	wire [4-1:0] node32438;
	wire [4-1:0] node32441;
	wire [4-1:0] node32442;
	wire [4-1:0] node32443;
	wire [4-1:0] node32445;
	wire [4-1:0] node32446;
	wire [4-1:0] node32450;
	wire [4-1:0] node32451;
	wire [4-1:0] node32454;
	wire [4-1:0] node32457;
	wire [4-1:0] node32458;
	wire [4-1:0] node32459;
	wire [4-1:0] node32462;
	wire [4-1:0] node32465;
	wire [4-1:0] node32467;
	wire [4-1:0] node32470;
	wire [4-1:0] node32471;
	wire [4-1:0] node32472;
	wire [4-1:0] node32473;
	wire [4-1:0] node32476;
	wire [4-1:0] node32477;
	wire [4-1:0] node32478;
	wire [4-1:0] node32481;
	wire [4-1:0] node32484;
	wire [4-1:0] node32485;
	wire [4-1:0] node32489;
	wire [4-1:0] node32490;
	wire [4-1:0] node32494;
	wire [4-1:0] node32495;
	wire [4-1:0] node32496;
	wire [4-1:0] node32497;
	wire [4-1:0] node32500;
	wire [4-1:0] node32503;
	wire [4-1:0] node32506;
	wire [4-1:0] node32507;
	wire [4-1:0] node32511;
	wire [4-1:0] node32512;
	wire [4-1:0] node32513;
	wire [4-1:0] node32514;
	wire [4-1:0] node32515;
	wire [4-1:0] node32516;
	wire [4-1:0] node32517;
	wire [4-1:0] node32518;
	wire [4-1:0] node32519;
	wire [4-1:0] node32521;
	wire [4-1:0] node32523;
	wire [4-1:0] node32527;
	wire [4-1:0] node32528;
	wire [4-1:0] node32529;
	wire [4-1:0] node32532;
	wire [4-1:0] node32536;
	wire [4-1:0] node32537;
	wire [4-1:0] node32538;
	wire [4-1:0] node32539;
	wire [4-1:0] node32540;
	wire [4-1:0] node32544;
	wire [4-1:0] node32548;
	wire [4-1:0] node32549;
	wire [4-1:0] node32550;
	wire [4-1:0] node32554;
	wire [4-1:0] node32555;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32562;
	wire [4-1:0] node32564;
	wire [4-1:0] node32567;
	wire [4-1:0] node32568;
	wire [4-1:0] node32570;
	wire [4-1:0] node32573;
	wire [4-1:0] node32575;
	wire [4-1:0] node32578;
	wire [4-1:0] node32579;
	wire [4-1:0] node32580;
	wire [4-1:0] node32581;
	wire [4-1:0] node32583;
	wire [4-1:0] node32586;
	wire [4-1:0] node32588;
	wire [4-1:0] node32591;
	wire [4-1:0] node32592;
	wire [4-1:0] node32594;
	wire [4-1:0] node32597;
	wire [4-1:0] node32599;
	wire [4-1:0] node32602;
	wire [4-1:0] node32603;
	wire [4-1:0] node32604;
	wire [4-1:0] node32606;
	wire [4-1:0] node32610;
	wire [4-1:0] node32611;
	wire [4-1:0] node32613;
	wire [4-1:0] node32616;
	wire [4-1:0] node32618;
	wire [4-1:0] node32621;
	wire [4-1:0] node32622;
	wire [4-1:0] node32623;
	wire [4-1:0] node32624;
	wire [4-1:0] node32625;
	wire [4-1:0] node32626;
	wire [4-1:0] node32631;
	wire [4-1:0] node32632;
	wire [4-1:0] node32633;
	wire [4-1:0] node32634;
	wire [4-1:0] node32635;
	wire [4-1:0] node32638;
	wire [4-1:0] node32643;
	wire [4-1:0] node32644;
	wire [4-1:0] node32647;
	wire [4-1:0] node32648;
	wire [4-1:0] node32652;
	wire [4-1:0] node32653;
	wire [4-1:0] node32654;
	wire [4-1:0] node32655;
	wire [4-1:0] node32656;
	wire [4-1:0] node32660;
	wire [4-1:0] node32661;
	wire [4-1:0] node32665;
	wire [4-1:0] node32666;
	wire [4-1:0] node32669;
	wire [4-1:0] node32670;
	wire [4-1:0] node32674;
	wire [4-1:0] node32675;
	wire [4-1:0] node32676;
	wire [4-1:0] node32677;
	wire [4-1:0] node32678;
	wire [4-1:0] node32682;
	wire [4-1:0] node32683;
	wire [4-1:0] node32686;
	wire [4-1:0] node32690;
	wire [4-1:0] node32691;
	wire [4-1:0] node32692;
	wire [4-1:0] node32695;
	wire [4-1:0] node32699;
	wire [4-1:0] node32700;
	wire [4-1:0] node32701;
	wire [4-1:0] node32703;
	wire [4-1:0] node32704;
	wire [4-1:0] node32707;
	wire [4-1:0] node32708;
	wire [4-1:0] node32712;
	wire [4-1:0] node32713;
	wire [4-1:0] node32714;
	wire [4-1:0] node32715;
	wire [4-1:0] node32719;
	wire [4-1:0] node32720;
	wire [4-1:0] node32724;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32730;
	wire [4-1:0] node32731;
	wire [4-1:0] node32735;
	wire [4-1:0] node32736;
	wire [4-1:0] node32737;
	wire [4-1:0] node32738;
	wire [4-1:0] node32741;
	wire [4-1:0] node32742;
	wire [4-1:0] node32744;
	wire [4-1:0] node32747;
	wire [4-1:0] node32750;
	wire [4-1:0] node32751;
	wire [4-1:0] node32752;
	wire [4-1:0] node32756;
	wire [4-1:0] node32757;
	wire [4-1:0] node32761;
	wire [4-1:0] node32762;
	wire [4-1:0] node32764;
	wire [4-1:0] node32767;
	wire [4-1:0] node32768;
	wire [4-1:0] node32771;
	wire [4-1:0] node32772;
	wire [4-1:0] node32776;
	wire [4-1:0] node32777;
	wire [4-1:0] node32778;
	wire [4-1:0] node32779;
	wire [4-1:0] node32781;
	wire [4-1:0] node32782;
	wire [4-1:0] node32786;
	wire [4-1:0] node32787;
	wire [4-1:0] node32789;
	wire [4-1:0] node32792;
	wire [4-1:0] node32793;
	wire [4-1:0] node32797;
	wire [4-1:0] node32798;
	wire [4-1:0] node32799;
	wire [4-1:0] node32800;
	wire [4-1:0] node32802;
	wire [4-1:0] node32803;
	wire [4-1:0] node32804;
	wire [4-1:0] node32809;
	wire [4-1:0] node32810;
	wire [4-1:0] node32813;
	wire [4-1:0] node32816;
	wire [4-1:0] node32817;
	wire [4-1:0] node32818;
	wire [4-1:0] node32819;
	wire [4-1:0] node32822;
	wire [4-1:0] node32826;
	wire [4-1:0] node32827;
	wire [4-1:0] node32829;
	wire [4-1:0] node32830;
	wire [4-1:0] node32833;
	wire [4-1:0] node32836;
	wire [4-1:0] node32837;
	wire [4-1:0] node32841;
	wire [4-1:0] node32842;
	wire [4-1:0] node32843;
	wire [4-1:0] node32846;
	wire [4-1:0] node32849;
	wire [4-1:0] node32850;
	wire [4-1:0] node32851;
	wire [4-1:0] node32854;
	wire [4-1:0] node32857;
	wire [4-1:0] node32859;
	wire [4-1:0] node32861;
	wire [4-1:0] node32864;
	wire [4-1:0] node32865;
	wire [4-1:0] node32866;
	wire [4-1:0] node32867;
	wire [4-1:0] node32868;
	wire [4-1:0] node32869;
	wire [4-1:0] node32873;
	wire [4-1:0] node32874;
	wire [4-1:0] node32875;
	wire [4-1:0] node32880;
	wire [4-1:0] node32881;
	wire [4-1:0] node32882;
	wire [4-1:0] node32883;
	wire [4-1:0] node32888;
	wire [4-1:0] node32889;
	wire [4-1:0] node32890;
	wire [4-1:0] node32895;
	wire [4-1:0] node32896;
	wire [4-1:0] node32897;
	wire [4-1:0] node32900;
	wire [4-1:0] node32901;
	wire [4-1:0] node32903;
	wire [4-1:0] node32907;
	wire [4-1:0] node32908;
	wire [4-1:0] node32909;
	wire [4-1:0] node32913;
	wire [4-1:0] node32914;
	wire [4-1:0] node32918;
	wire [4-1:0] node32919;
	wire [4-1:0] node32920;
	wire [4-1:0] node32921;
	wire [4-1:0] node32922;
	wire [4-1:0] node32923;
	wire [4-1:0] node32924;
	wire [4-1:0] node32930;
	wire [4-1:0] node32932;
	wire [4-1:0] node32933;
	wire [4-1:0] node32934;
	wire [4-1:0] node32937;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32943;
	wire [4-1:0] node32944;
	wire [4-1:0] node32945;
	wire [4-1:0] node32949;
	wire [4-1:0] node32951;
	wire [4-1:0] node32954;
	wire [4-1:0] node32955;
	wire [4-1:0] node32958;
	wire [4-1:0] node32960;
	wire [4-1:0] node32963;
	wire [4-1:0] node32964;
	wire [4-1:0] node32968;
	wire [4-1:0] node32969;
	wire [4-1:0] node32970;
	wire [4-1:0] node32971;
	wire [4-1:0] node32973;
	wire [4-1:0] node32974;
	wire [4-1:0] node32977;
	wire [4-1:0] node32980;
	wire [4-1:0] node32981;
	wire [4-1:0] node32982;
	wire [4-1:0] node32985;
	wire [4-1:0] node32988;
	wire [4-1:0] node32990;
	wire [4-1:0] node32993;
	wire [4-1:0] node32994;
	wire [4-1:0] node32998;
	wire [4-1:0] node33000;
	wire [4-1:0] node33002;
	wire [4-1:0] node33005;
	wire [4-1:0] node33006;
	wire [4-1:0] node33007;
	wire [4-1:0] node33008;
	wire [4-1:0] node33009;
	wire [4-1:0] node33010;
	wire [4-1:0] node33011;
	wire [4-1:0] node33013;
	wire [4-1:0] node33014;
	wire [4-1:0] node33018;
	wire [4-1:0] node33019;
	wire [4-1:0] node33020;
	wire [4-1:0] node33021;
	wire [4-1:0] node33025;
	wire [4-1:0] node33027;
	wire [4-1:0] node33030;
	wire [4-1:0] node33032;
	wire [4-1:0] node33035;
	wire [4-1:0] node33036;
	wire [4-1:0] node33037;
	wire [4-1:0] node33038;
	wire [4-1:0] node33041;
	wire [4-1:0] node33045;
	wire [4-1:0] node33046;
	wire [4-1:0] node33047;
	wire [4-1:0] node33051;
	wire [4-1:0] node33052;
	wire [4-1:0] node33053;
	wire [4-1:0] node33056;
	wire [4-1:0] node33060;
	wire [4-1:0] node33061;
	wire [4-1:0] node33062;
	wire [4-1:0] node33063;
	wire [4-1:0] node33064;
	wire [4-1:0] node33066;
	wire [4-1:0] node33070;
	wire [4-1:0] node33071;
	wire [4-1:0] node33074;
	wire [4-1:0] node33076;
	wire [4-1:0] node33079;
	wire [4-1:0] node33082;
	wire [4-1:0] node33083;
	wire [4-1:0] node33086;
	wire [4-1:0] node33089;
	wire [4-1:0] node33090;
	wire [4-1:0] node33091;
	wire [4-1:0] node33092;
	wire [4-1:0] node33093;
	wire [4-1:0] node33094;
	wire [4-1:0] node33098;
	wire [4-1:0] node33100;
	wire [4-1:0] node33104;
	wire [4-1:0] node33105;
	wire [4-1:0] node33107;
	wire [4-1:0] node33108;
	wire [4-1:0] node33111;
	wire [4-1:0] node33114;
	wire [4-1:0] node33116;
	wire [4-1:0] node33118;
	wire [4-1:0] node33121;
	wire [4-1:0] node33122;
	wire [4-1:0] node33123;
	wire [4-1:0] node33124;
	wire [4-1:0] node33127;
	wire [4-1:0] node33130;
	wire [4-1:0] node33131;
	wire [4-1:0] node33133;
	wire [4-1:0] node33137;
	wire [4-1:0] node33138;
	wire [4-1:0] node33141;
	wire [4-1:0] node33144;
	wire [4-1:0] node33145;
	wire [4-1:0] node33146;
	wire [4-1:0] node33147;
	wire [4-1:0] node33148;
	wire [4-1:0] node33149;
	wire [4-1:0] node33152;
	wire [4-1:0] node33155;
	wire [4-1:0] node33156;
	wire [4-1:0] node33159;
	wire [4-1:0] node33162;
	wire [4-1:0] node33163;
	wire [4-1:0] node33164;
	wire [4-1:0] node33168;
	wire [4-1:0] node33169;
	wire [4-1:0] node33170;
	wire [4-1:0] node33172;
	wire [4-1:0] node33175;
	wire [4-1:0] node33177;
	wire [4-1:0] node33180;
	wire [4-1:0] node33181;
	wire [4-1:0] node33185;
	wire [4-1:0] node33186;
	wire [4-1:0] node33187;
	wire [4-1:0] node33188;
	wire [4-1:0] node33189;
	wire [4-1:0] node33191;
	wire [4-1:0] node33194;
	wire [4-1:0] node33195;
	wire [4-1:0] node33199;
	wire [4-1:0] node33201;
	wire [4-1:0] node33202;
	wire [4-1:0] node33206;
	wire [4-1:0] node33207;
	wire [4-1:0] node33208;
	wire [4-1:0] node33211;
	wire [4-1:0] node33215;
	wire [4-1:0] node33216;
	wire [4-1:0] node33220;
	wire [4-1:0] node33221;
	wire [4-1:0] node33222;
	wire [4-1:0] node33223;
	wire [4-1:0] node33224;
	wire [4-1:0] node33226;
	wire [4-1:0] node33227;
	wire [4-1:0] node33230;
	wire [4-1:0] node33233;
	wire [4-1:0] node33234;
	wire [4-1:0] node33235;
	wire [4-1:0] node33238;
	wire [4-1:0] node33242;
	wire [4-1:0] node33243;
	wire [4-1:0] node33244;
	wire [4-1:0] node33247;
	wire [4-1:0] node33250;
	wire [4-1:0] node33251;
	wire [4-1:0] node33254;
	wire [4-1:0] node33257;
	wire [4-1:0] node33258;
	wire [4-1:0] node33260;
	wire [4-1:0] node33261;
	wire [4-1:0] node33262;
	wire [4-1:0] node33266;
	wire [4-1:0] node33267;
	wire [4-1:0] node33270;
	wire [4-1:0] node33273;
	wire [4-1:0] node33274;
	wire [4-1:0] node33275;
	wire [4-1:0] node33279;
	wire [4-1:0] node33280;
	wire [4-1:0] node33283;
	wire [4-1:0] node33286;
	wire [4-1:0] node33287;
	wire [4-1:0] node33288;
	wire [4-1:0] node33291;
	wire [4-1:0] node33294;
	wire [4-1:0] node33295;
	wire [4-1:0] node33296;
	wire [4-1:0] node33297;
	wire [4-1:0] node33301;
	wire [4-1:0] node33302;
	wire [4-1:0] node33303;
	wire [4-1:0] node33306;
	wire [4-1:0] node33309;
	wire [4-1:0] node33311;
	wire [4-1:0] node33314;
	wire [4-1:0] node33315;
	wire [4-1:0] node33318;
	wire [4-1:0] node33321;
	wire [4-1:0] node33322;
	wire [4-1:0] node33323;
	wire [4-1:0] node33324;
	wire [4-1:0] node33325;
	wire [4-1:0] node33329;
	wire [4-1:0] node33330;
	wire [4-1:0] node33335;
	wire [4-1:0] node33336;
	wire [4-1:0] node33337;
	wire [4-1:0] node33338;
	wire [4-1:0] node33342;
	wire [4-1:0] node33343;
	wire [4-1:0] node33348;
	wire [4-1:0] node33349;
	wire [4-1:0] node33350;
	wire [4-1:0] node33351;
	wire [4-1:0] node33352;
	wire [4-1:0] node33353;
	wire [4-1:0] node33354;
	wire [4-1:0] node33355;
	wire [4-1:0] node33356;
	wire [4-1:0] node33357;
	wire [4-1:0] node33359;
	wire [4-1:0] node33363;
	wire [4-1:0] node33364;
	wire [4-1:0] node33365;
	wire [4-1:0] node33366;
	wire [4-1:0] node33370;
	wire [4-1:0] node33373;
	wire [4-1:0] node33375;
	wire [4-1:0] node33378;
	wire [4-1:0] node33379;
	wire [4-1:0] node33381;
	wire [4-1:0] node33384;
	wire [4-1:0] node33385;
	wire [4-1:0] node33387;
	wire [4-1:0] node33388;
	wire [4-1:0] node33391;
	wire [4-1:0] node33394;
	wire [4-1:0] node33395;
	wire [4-1:0] node33399;
	wire [4-1:0] node33400;
	wire [4-1:0] node33402;
	wire [4-1:0] node33403;
	wire [4-1:0] node33404;
	wire [4-1:0] node33406;
	wire [4-1:0] node33410;
	wire [4-1:0] node33413;
	wire [4-1:0] node33414;
	wire [4-1:0] node33416;
	wire [4-1:0] node33417;
	wire [4-1:0] node33421;
	wire [4-1:0] node33422;
	wire [4-1:0] node33425;
	wire [4-1:0] node33426;
	wire [4-1:0] node33428;
	wire [4-1:0] node33432;
	wire [4-1:0] node33433;
	wire [4-1:0] node33434;
	wire [4-1:0] node33435;
	wire [4-1:0] node33437;
	wire [4-1:0] node33438;
	wire [4-1:0] node33442;
	wire [4-1:0] node33443;
	wire [4-1:0] node33444;
	wire [4-1:0] node33445;
	wire [4-1:0] node33449;
	wire [4-1:0] node33450;
	wire [4-1:0] node33453;
	wire [4-1:0] node33454;
	wire [4-1:0] node33458;
	wire [4-1:0] node33461;
	wire [4-1:0] node33462;
	wire [4-1:0] node33464;
	wire [4-1:0] node33466;
	wire [4-1:0] node33469;
	wire [4-1:0] node33470;
	wire [4-1:0] node33471;
	wire [4-1:0] node33474;
	wire [4-1:0] node33477;
	wire [4-1:0] node33478;
	wire [4-1:0] node33482;
	wire [4-1:0] node33483;
	wire [4-1:0] node33484;
	wire [4-1:0] node33486;
	wire [4-1:0] node33487;
	wire [4-1:0] node33489;
	wire [4-1:0] node33492;
	wire [4-1:0] node33494;
	wire [4-1:0] node33497;
	wire [4-1:0] node33498;
	wire [4-1:0] node33499;
	wire [4-1:0] node33504;
	wire [4-1:0] node33505;
	wire [4-1:0] node33506;
	wire [4-1:0] node33508;
	wire [4-1:0] node33509;
	wire [4-1:0] node33514;
	wire [4-1:0] node33515;
	wire [4-1:0] node33516;
	wire [4-1:0] node33517;
	wire [4-1:0] node33519;
	wire [4-1:0] node33524;
	wire [4-1:0] node33525;
	wire [4-1:0] node33529;
	wire [4-1:0] node33530;
	wire [4-1:0] node33531;
	wire [4-1:0] node33532;
	wire [4-1:0] node33533;
	wire [4-1:0] node33534;
	wire [4-1:0] node33536;
	wire [4-1:0] node33539;
	wire [4-1:0] node33540;
	wire [4-1:0] node33543;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33549;
	wire [4-1:0] node33552;
	wire [4-1:0] node33553;
	wire [4-1:0] node33556;
	wire [4-1:0] node33559;
	wire [4-1:0] node33560;
	wire [4-1:0] node33561;
	wire [4-1:0] node33563;
	wire [4-1:0] node33566;
	wire [4-1:0] node33567;
	wire [4-1:0] node33570;
	wire [4-1:0] node33573;
	wire [4-1:0] node33574;
	wire [4-1:0] node33576;
	wire [4-1:0] node33579;
	wire [4-1:0] node33581;
	wire [4-1:0] node33584;
	wire [4-1:0] node33585;
	wire [4-1:0] node33586;
	wire [4-1:0] node33588;
	wire [4-1:0] node33590;
	wire [4-1:0] node33591;
	wire [4-1:0] node33595;
	wire [4-1:0] node33596;
	wire [4-1:0] node33597;
	wire [4-1:0] node33601;
	wire [4-1:0] node33603;
	wire [4-1:0] node33606;
	wire [4-1:0] node33607;
	wire [4-1:0] node33609;
	wire [4-1:0] node33612;
	wire [4-1:0] node33613;
	wire [4-1:0] node33614;
	wire [4-1:0] node33618;
	wire [4-1:0] node33620;
	wire [4-1:0] node33623;
	wire [4-1:0] node33624;
	wire [4-1:0] node33625;
	wire [4-1:0] node33626;
	wire [4-1:0] node33627;
	wire [4-1:0] node33628;
	wire [4-1:0] node33629;
	wire [4-1:0] node33632;
	wire [4-1:0] node33636;
	wire [4-1:0] node33637;
	wire [4-1:0] node33638;
	wire [4-1:0] node33641;
	wire [4-1:0] node33644;
	wire [4-1:0] node33646;
	wire [4-1:0] node33649;
	wire [4-1:0] node33650;
	wire [4-1:0] node33652;
	wire [4-1:0] node33655;
	wire [4-1:0] node33657;
	wire [4-1:0] node33658;
	wire [4-1:0] node33662;
	wire [4-1:0] node33663;
	wire [4-1:0] node33664;
	wire [4-1:0] node33665;
	wire [4-1:0] node33667;
	wire [4-1:0] node33671;
	wire [4-1:0] node33672;
	wire [4-1:0] node33673;
	wire [4-1:0] node33675;
	wire [4-1:0] node33679;
	wire [4-1:0] node33681;
	wire [4-1:0] node33682;
	wire [4-1:0] node33686;
	wire [4-1:0] node33687;
	wire [4-1:0] node33688;
	wire [4-1:0] node33689;
	wire [4-1:0] node33693;
	wire [4-1:0] node33694;
	wire [4-1:0] node33697;
	wire [4-1:0] node33700;
	wire [4-1:0] node33701;
	wire [4-1:0] node33702;
	wire [4-1:0] node33706;
	wire [4-1:0] node33708;
	wire [4-1:0] node33711;
	wire [4-1:0] node33712;
	wire [4-1:0] node33713;
	wire [4-1:0] node33714;
	wire [4-1:0] node33715;
	wire [4-1:0] node33719;
	wire [4-1:0] node33721;
	wire [4-1:0] node33724;
	wire [4-1:0] node33725;
	wire [4-1:0] node33726;
	wire [4-1:0] node33730;
	wire [4-1:0] node33732;
	wire [4-1:0] node33735;
	wire [4-1:0] node33736;
	wire [4-1:0] node33739;
	wire [4-1:0] node33742;
	wire [4-1:0] node33743;
	wire [4-1:0] node33744;
	wire [4-1:0] node33745;
	wire [4-1:0] node33746;
	wire [4-1:0] node33747;
	wire [4-1:0] node33748;
	wire [4-1:0] node33749;
	wire [4-1:0] node33753;
	wire [4-1:0] node33755;
	wire [4-1:0] node33757;
	wire [4-1:0] node33760;
	wire [4-1:0] node33761;
	wire [4-1:0] node33764;
	wire [4-1:0] node33765;
	wire [4-1:0] node33769;
	wire [4-1:0] node33770;
	wire [4-1:0] node33771;
	wire [4-1:0] node33772;
	wire [4-1:0] node33774;
	wire [4-1:0] node33777;
	wire [4-1:0] node33779;
	wire [4-1:0] node33782;
	wire [4-1:0] node33783;
	wire [4-1:0] node33784;
	wire [4-1:0] node33787;
	wire [4-1:0] node33789;
	wire [4-1:0] node33792;
	wire [4-1:0] node33793;
	wire [4-1:0] node33797;
	wire [4-1:0] node33798;
	wire [4-1:0] node33799;
	wire [4-1:0] node33802;
	wire [4-1:0] node33803;
	wire [4-1:0] node33806;
	wire [4-1:0] node33809;
	wire [4-1:0] node33811;
	wire [4-1:0] node33812;
	wire [4-1:0] node33816;
	wire [4-1:0] node33817;
	wire [4-1:0] node33818;
	wire [4-1:0] node33819;
	wire [4-1:0] node33820;
	wire [4-1:0] node33821;
	wire [4-1:0] node33824;
	wire [4-1:0] node33828;
	wire [4-1:0] node33829;
	wire [4-1:0] node33832;
	wire [4-1:0] node33835;
	wire [4-1:0] node33836;
	wire [4-1:0] node33839;
	wire [4-1:0] node33842;
	wire [4-1:0] node33843;
	wire [4-1:0] node33844;
	wire [4-1:0] node33846;
	wire [4-1:0] node33849;
	wire [4-1:0] node33850;
	wire [4-1:0] node33854;
	wire [4-1:0] node33855;
	wire [4-1:0] node33857;
	wire [4-1:0] node33858;
	wire [4-1:0] node33862;
	wire [4-1:0] node33863;
	wire [4-1:0] node33866;
	wire [4-1:0] node33869;
	wire [4-1:0] node33870;
	wire [4-1:0] node33871;
	wire [4-1:0] node33872;
	wire [4-1:0] node33874;
	wire [4-1:0] node33876;
	wire [4-1:0] node33879;
	wire [4-1:0] node33881;
	wire [4-1:0] node33883;
	wire [4-1:0] node33886;
	wire [4-1:0] node33887;
	wire [4-1:0] node33888;
	wire [4-1:0] node33890;
	wire [4-1:0] node33893;
	wire [4-1:0] node33894;
	wire [4-1:0] node33897;
	wire [4-1:0] node33900;
	wire [4-1:0] node33901;
	wire [4-1:0] node33902;
	wire [4-1:0] node33905;
	wire [4-1:0] node33908;
	wire [4-1:0] node33909;
	wire [4-1:0] node33913;
	wire [4-1:0] node33914;
	wire [4-1:0] node33915;
	wire [4-1:0] node33917;
	wire [4-1:0] node33920;
	wire [4-1:0] node33921;
	wire [4-1:0] node33923;
	wire [4-1:0] node33926;
	wire [4-1:0] node33927;
	wire [4-1:0] node33930;
	wire [4-1:0] node33933;
	wire [4-1:0] node33934;
	wire [4-1:0] node33936;
	wire [4-1:0] node33937;
	wire [4-1:0] node33941;
	wire [4-1:0] node33942;
	wire [4-1:0] node33943;
	wire [4-1:0] node33944;
	wire [4-1:0] node33947;
	wire [4-1:0] node33950;
	wire [4-1:0] node33951;
	wire [4-1:0] node33955;
	wire [4-1:0] node33956;
	wire [4-1:0] node33960;
	wire [4-1:0] node33961;
	wire [4-1:0] node33962;
	wire [4-1:0] node33963;
	wire [4-1:0] node33964;
	wire [4-1:0] node33965;
	wire [4-1:0] node33968;
	wire [4-1:0] node33970;
	wire [4-1:0] node33971;
	wire [4-1:0] node33975;
	wire [4-1:0] node33976;
	wire [4-1:0] node33977;
	wire [4-1:0] node33978;
	wire [4-1:0] node33981;
	wire [4-1:0] node33985;
	wire [4-1:0] node33986;
	wire [4-1:0] node33990;
	wire [4-1:0] node33991;
	wire [4-1:0] node33993;
	wire [4-1:0] node33994;
	wire [4-1:0] node33998;
	wire [4-1:0] node33999;
	wire [4-1:0] node34001;
	wire [4-1:0] node34005;
	wire [4-1:0] node34006;
	wire [4-1:0] node34007;
	wire [4-1:0] node34008;
	wire [4-1:0] node34009;
	wire [4-1:0] node34012;
	wire [4-1:0] node34015;
	wire [4-1:0] node34016;
	wire [4-1:0] node34017;
	wire [4-1:0] node34021;
	wire [4-1:0] node34022;
	wire [4-1:0] node34026;
	wire [4-1:0] node34027;
	wire [4-1:0] node34028;
	wire [4-1:0] node34032;
	wire [4-1:0] node34034;
	wire [4-1:0] node34037;
	wire [4-1:0] node34038;
	wire [4-1:0] node34039;
	wire [4-1:0] node34041;
	wire [4-1:0] node34044;
	wire [4-1:0] node34045;
	wire [4-1:0] node34049;
	wire [4-1:0] node34052;
	wire [4-1:0] node34053;
	wire [4-1:0] node34054;
	wire [4-1:0] node34055;
	wire [4-1:0] node34056;
	wire [4-1:0] node34057;
	wire [4-1:0] node34059;
	wire [4-1:0] node34060;
	wire [4-1:0] node34065;
	wire [4-1:0] node34067;
	wire [4-1:0] node34068;
	wire [4-1:0] node34072;
	wire [4-1:0] node34073;
	wire [4-1:0] node34074;
	wire [4-1:0] node34077;
	wire [4-1:0] node34080;
	wire [4-1:0] node34082;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34089;
	wire [4-1:0] node34092;
	wire [4-1:0] node34095;
	wire [4-1:0] node34098;
	wire [4-1:0] node34099;
	wire [4-1:0] node34100;
	wire [4-1:0] node34101;
	wire [4-1:0] node34102;
	wire [4-1:0] node34105;
	wire [4-1:0] node34108;
	wire [4-1:0] node34109;
	wire [4-1:0] node34113;
	wire [4-1:0] node34114;
	wire [4-1:0] node34115;
	wire [4-1:0] node34118;
	wire [4-1:0] node34121;
	wire [4-1:0] node34124;
	wire [4-1:0] node34125;
	wire [4-1:0] node34126;
	wire [4-1:0] node34128;
	wire [4-1:0] node34131;
	wire [4-1:0] node34132;
	wire [4-1:0] node34136;
	wire [4-1:0] node34139;
	wire [4-1:0] node34140;
	wire [4-1:0] node34141;
	wire [4-1:0] node34142;
	wire [4-1:0] node34143;
	wire [4-1:0] node34144;
	wire [4-1:0] node34145;
	wire [4-1:0] node34147;
	wire [4-1:0] node34150;
	wire [4-1:0] node34152;
	wire [4-1:0] node34155;
	wire [4-1:0] node34156;
	wire [4-1:0] node34158;
	wire [4-1:0] node34161;
	wire [4-1:0] node34163;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34168;
	wire [4-1:0] node34170;
	wire [4-1:0] node34173;
	wire [4-1:0] node34175;
	wire [4-1:0] node34178;
	wire [4-1:0] node34179;
	wire [4-1:0] node34181;
	wire [4-1:0] node34184;
	wire [4-1:0] node34186;
	wire [4-1:0] node34189;
	wire [4-1:0] node34190;
	wire [4-1:0] node34191;
	wire [4-1:0] node34192;
	wire [4-1:0] node34193;
	wire [4-1:0] node34194;
	wire [4-1:0] node34197;
	wire [4-1:0] node34200;
	wire [4-1:0] node34202;
	wire [4-1:0] node34205;
	wire [4-1:0] node34206;
	wire [4-1:0] node34207;
	wire [4-1:0] node34208;
	wire [4-1:0] node34211;
	wire [4-1:0] node34215;
	wire [4-1:0] node34217;
	wire [4-1:0] node34220;
	wire [4-1:0] node34221;
	wire [4-1:0] node34222;
	wire [4-1:0] node34224;
	wire [4-1:0] node34225;
	wire [4-1:0] node34228;
	wire [4-1:0] node34231;
	wire [4-1:0] node34232;
	wire [4-1:0] node34233;
	wire [4-1:0] node34237;
	wire [4-1:0] node34238;
	wire [4-1:0] node34242;
	wire [4-1:0] node34243;
	wire [4-1:0] node34247;
	wire [4-1:0] node34248;
	wire [4-1:0] node34251;
	wire [4-1:0] node34254;
	wire [4-1:0] node34255;
	wire [4-1:0] node34256;
	wire [4-1:0] node34257;
	wire [4-1:0] node34258;
	wire [4-1:0] node34259;
	wire [4-1:0] node34260;
	wire [4-1:0] node34264;
	wire [4-1:0] node34265;
	wire [4-1:0] node34267;
	wire [4-1:0] node34270;
	wire [4-1:0] node34271;
	wire [4-1:0] node34274;
	wire [4-1:0] node34278;
	wire [4-1:0] node34279;
	wire [4-1:0] node34281;
	wire [4-1:0] node34282;
	wire [4-1:0] node34284;
	wire [4-1:0] node34287;
	wire [4-1:0] node34289;
	wire [4-1:0] node34293;
	wire [4-1:0] node34294;
	wire [4-1:0] node34295;
	wire [4-1:0] node34299;
	wire [4-1:0] node34300;
	wire [4-1:0] node34304;
	wire [4-1:0] node34305;
	wire [4-1:0] node34306;
	wire [4-1:0] node34307;
	wire [4-1:0] node34309;
	wire [4-1:0] node34312;
	wire [4-1:0] node34315;
	wire [4-1:0] node34316;
	wire [4-1:0] node34317;
	wire [4-1:0] node34321;
	wire [4-1:0] node34324;
	wire [4-1:0] node34325;
	wire [4-1:0] node34326;
	wire [4-1:0] node34327;
	wire [4-1:0] node34332;
	wire [4-1:0] node34333;
	wire [4-1:0] node34334;
	wire [4-1:0] node34339;
	wire [4-1:0] node34340;
	wire [4-1:0] node34341;
	wire [4-1:0] node34342;
	wire [4-1:0] node34343;
	wire [4-1:0] node34344;
	wire [4-1:0] node34348;
	wire [4-1:0] node34349;
	wire [4-1:0] node34353;
	wire [4-1:0] node34354;
	wire [4-1:0] node34355;
	wire [4-1:0] node34359;
	wire [4-1:0] node34361;
	wire [4-1:0] node34364;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34367;
	wire [4-1:0] node34368;
	wire [4-1:0] node34370;
	wire [4-1:0] node34373;
	wire [4-1:0] node34374;
	wire [4-1:0] node34377;
	wire [4-1:0] node34380;
	wire [4-1:0] node34381;
	wire [4-1:0] node34382;
	wire [4-1:0] node34386;
	wire [4-1:0] node34387;
	wire [4-1:0] node34391;
	wire [4-1:0] node34392;
	wire [4-1:0] node34393;
	wire [4-1:0] node34394;
	wire [4-1:0] node34397;
	wire [4-1:0] node34400;
	wire [4-1:0] node34402;
	wire [4-1:0] node34405;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34411;
	wire [4-1:0] node34412;
	wire [4-1:0] node34415;
	wire [4-1:0] node34418;
	wire [4-1:0] node34419;
	wire [4-1:0] node34420;
	wire [4-1:0] node34423;
	wire [4-1:0] node34426;
	wire [4-1:0] node34427;
	wire [4-1:0] node34430;
	wire [4-1:0] node34433;
	wire [4-1:0] node34434;
	wire [4-1:0] node34435;
	wire [4-1:0] node34436;
	wire [4-1:0] node34437;
	wire [4-1:0] node34441;
	wire [4-1:0] node34442;
	wire [4-1:0] node34447;
	wire [4-1:0] node34448;
	wire [4-1:0] node34449;
	wire [4-1:0] node34450;
	wire [4-1:0] node34454;
	wire [4-1:0] node34455;
	wire [4-1:0] node34460;
	wire [4-1:0] node34461;
	wire [4-1:0] node34462;
	wire [4-1:0] node34463;
	wire [4-1:0] node34464;
	wire [4-1:0] node34465;
	wire [4-1:0] node34466;
	wire [4-1:0] node34467;
	wire [4-1:0] node34468;
	wire [4-1:0] node34470;
	wire [4-1:0] node34471;
	wire [4-1:0] node34472;
	wire [4-1:0] node34476;
	wire [4-1:0] node34478;
	wire [4-1:0] node34481;
	wire [4-1:0] node34482;
	wire [4-1:0] node34485;
	wire [4-1:0] node34488;
	wire [4-1:0] node34489;
	wire [4-1:0] node34490;
	wire [4-1:0] node34494;
	wire [4-1:0] node34496;
	wire [4-1:0] node34499;
	wire [4-1:0] node34500;
	wire [4-1:0] node34501;
	wire [4-1:0] node34502;
	wire [4-1:0] node34504;
	wire [4-1:0] node34505;
	wire [4-1:0] node34508;
	wire [4-1:0] node34511;
	wire [4-1:0] node34512;
	wire [4-1:0] node34514;
	wire [4-1:0] node34518;
	wire [4-1:0] node34519;
	wire [4-1:0] node34520;
	wire [4-1:0] node34523;
	wire [4-1:0] node34526;
	wire [4-1:0] node34527;
	wire [4-1:0] node34530;
	wire [4-1:0] node34533;
	wire [4-1:0] node34534;
	wire [4-1:0] node34535;
	wire [4-1:0] node34537;
	wire [4-1:0] node34541;
	wire [4-1:0] node34542;
	wire [4-1:0] node34545;
	wire [4-1:0] node34548;
	wire [4-1:0] node34549;
	wire [4-1:0] node34550;
	wire [4-1:0] node34551;
	wire [4-1:0] node34552;
	wire [4-1:0] node34554;
	wire [4-1:0] node34555;
	wire [4-1:0] node34558;
	wire [4-1:0] node34561;
	wire [4-1:0] node34563;
	wire [4-1:0] node34567;
	wire [4-1:0] node34568;
	wire [4-1:0] node34571;
	wire [4-1:0] node34574;
	wire [4-1:0] node34575;
	wire [4-1:0] node34576;
	wire [4-1:0] node34577;
	wire [4-1:0] node34578;
	wire [4-1:0] node34581;
	wire [4-1:0] node34584;
	wire [4-1:0] node34585;
	wire [4-1:0] node34589;
	wire [4-1:0] node34591;
	wire [4-1:0] node34593;
	wire [4-1:0] node34594;
	wire [4-1:0] node34597;
	wire [4-1:0] node34600;
	wire [4-1:0] node34601;
	wire [4-1:0] node34602;
	wire [4-1:0] node34605;
	wire [4-1:0] node34608;
	wire [4-1:0] node34609;
	wire [4-1:0] node34613;
	wire [4-1:0] node34614;
	wire [4-1:0] node34615;
	wire [4-1:0] node34616;
	wire [4-1:0] node34617;
	wire [4-1:0] node34620;
	wire [4-1:0] node34623;
	wire [4-1:0] node34625;
	wire [4-1:0] node34626;
	wire [4-1:0] node34627;
	wire [4-1:0] node34630;
	wire [4-1:0] node34633;
	wire [4-1:0] node34634;
	wire [4-1:0] node34638;
	wire [4-1:0] node34639;
	wire [4-1:0] node34640;
	wire [4-1:0] node34641;
	wire [4-1:0] node34644;
	wire [4-1:0] node34647;
	wire [4-1:0] node34648;
	wire [4-1:0] node34651;
	wire [4-1:0] node34654;
	wire [4-1:0] node34655;
	wire [4-1:0] node34658;
	wire [4-1:0] node34661;
	wire [4-1:0] node34662;
	wire [4-1:0] node34663;
	wire [4-1:0] node34664;
	wire [4-1:0] node34666;
	wire [4-1:0] node34667;
	wire [4-1:0] node34669;
	wire [4-1:0] node34672;
	wire [4-1:0] node34675;
	wire [4-1:0] node34676;
	wire [4-1:0] node34677;
	wire [4-1:0] node34681;
	wire [4-1:0] node34683;
	wire [4-1:0] node34684;
	wire [4-1:0] node34687;
	wire [4-1:0] node34690;
	wire [4-1:0] node34691;
	wire [4-1:0] node34692;
	wire [4-1:0] node34696;
	wire [4-1:0] node34697;
	wire [4-1:0] node34700;
	wire [4-1:0] node34703;
	wire [4-1:0] node34704;
	wire [4-1:0] node34705;
	wire [4-1:0] node34708;
	wire [4-1:0] node34711;
	wire [4-1:0] node34712;
	wire [4-1:0] node34714;
	wire [4-1:0] node34716;
	wire [4-1:0] node34719;
	wire [4-1:0] node34721;
	wire [4-1:0] node34722;
	wire [4-1:0] node34723;
	wire [4-1:0] node34727;
	wire [4-1:0] node34729;
	wire [4-1:0] node34732;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34735;
	wire [4-1:0] node34736;
	wire [4-1:0] node34737;
	wire [4-1:0] node34738;
	wire [4-1:0] node34741;
	wire [4-1:0] node34744;
	wire [4-1:0] node34745;
	wire [4-1:0] node34746;
	wire [4-1:0] node34750;
	wire [4-1:0] node34751;
	wire [4-1:0] node34752;
	wire [4-1:0] node34755;
	wire [4-1:0] node34760;
	wire [4-1:0] node34761;
	wire [4-1:0] node34765;
	wire [4-1:0] node34766;
	wire [4-1:0] node34767;
	wire [4-1:0] node34768;
	wire [4-1:0] node34769;
	wire [4-1:0] node34772;
	wire [4-1:0] node34775;
	wire [4-1:0] node34776;
	wire [4-1:0] node34777;
	wire [4-1:0] node34778;
	wire [4-1:0] node34782;
	wire [4-1:0] node34784;
	wire [4-1:0] node34787;
	wire [4-1:0] node34788;
	wire [4-1:0] node34791;
	wire [4-1:0] node34795;
	wire [4-1:0] node34796;
	wire [4-1:0] node34800;
	wire [4-1:0] node34801;
	wire [4-1:0] node34802;
	wire [4-1:0] node34803;
	wire [4-1:0] node34804;
	wire [4-1:0] node34808;
	wire [4-1:0] node34809;
	wire [4-1:0] node34813;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34816;
	wire [4-1:0] node34819;
	wire [4-1:0] node34823;
	wire [4-1:0] node34824;
	wire [4-1:0] node34825;
	wire [4-1:0] node34828;
	wire [4-1:0] node34831;
	wire [4-1:0] node34832;
	wire [4-1:0] node34835;
	wire [4-1:0] node34838;
	wire [4-1:0] node34839;
	wire [4-1:0] node34840;
	wire [4-1:0] node34841;
	wire [4-1:0] node34846;
	wire [4-1:0] node34847;
	wire [4-1:0] node34848;
	wire [4-1:0] node34853;
	wire [4-1:0] node34854;
	wire [4-1:0] node34855;
	wire [4-1:0] node34856;
	wire [4-1:0] node34857;
	wire [4-1:0] node34860;
	wire [4-1:0] node34863;
	wire [4-1:0] node34864;
	wire [4-1:0] node34867;
	wire [4-1:0] node34870;
	wire [4-1:0] node34871;
	wire [4-1:0] node34872;
	wire [4-1:0] node34873;
	wire [4-1:0] node34874;
	wire [4-1:0] node34875;
	wire [4-1:0] node34879;
	wire [4-1:0] node34880;
	wire [4-1:0] node34883;
	wire [4-1:0] node34886;
	wire [4-1:0] node34887;
	wire [4-1:0] node34888;
	wire [4-1:0] node34890;
	wire [4-1:0] node34893;
	wire [4-1:0] node34895;
	wire [4-1:0] node34899;
	wire [4-1:0] node34900;
	wire [4-1:0] node34901;
	wire [4-1:0] node34902;
	wire [4-1:0] node34905;
	wire [4-1:0] node34908;
	wire [4-1:0] node34910;
	wire [4-1:0] node34912;
	wire [4-1:0] node34915;
	wire [4-1:0] node34916;
	wire [4-1:0] node34917;
	wire [4-1:0] node34918;
	wire [4-1:0] node34922;
	wire [4-1:0] node34924;
	wire [4-1:0] node34927;
	wire [4-1:0] node34929;
	wire [4-1:0] node34932;
	wire [4-1:0] node34933;
	wire [4-1:0] node34934;
	wire [4-1:0] node34935;
	wire [4-1:0] node34938;
	wire [4-1:0] node34941;
	wire [4-1:0] node34942;
	wire [4-1:0] node34944;
	wire [4-1:0] node34947;
	wire [4-1:0] node34948;
	wire [4-1:0] node34951;
	wire [4-1:0] node34954;
	wire [4-1:0] node34955;
	wire [4-1:0] node34958;
	wire [4-1:0] node34961;
	wire [4-1:0] node34962;
	wire [4-1:0] node34963;
	wire [4-1:0] node34967;
	wire [4-1:0] node34968;
	wire [4-1:0] node34972;
	wire [4-1:0] node34973;
	wire [4-1:0] node34974;
	wire [4-1:0] node34975;
	wire [4-1:0] node34976;
	wire [4-1:0] node34977;
	wire [4-1:0] node34978;
	wire [4-1:0] node34979;
	wire [4-1:0] node34983;
	wire [4-1:0] node34985;
	wire [4-1:0] node34988;
	wire [4-1:0] node34989;
	wire [4-1:0] node34990;
	wire [4-1:0] node34994;
	wire [4-1:0] node34995;
	wire [4-1:0] node34999;
	wire [4-1:0] node35000;
	wire [4-1:0] node35001;
	wire [4-1:0] node35002;
	wire [4-1:0] node35003;
	wire [4-1:0] node35006;
	wire [4-1:0] node35009;
	wire [4-1:0] node35011;
	wire [4-1:0] node35014;
	wire [4-1:0] node35015;
	wire [4-1:0] node35016;
	wire [4-1:0] node35018;
	wire [4-1:0] node35021;
	wire [4-1:0] node35022;
	wire [4-1:0] node35025;
	wire [4-1:0] node35028;
	wire [4-1:0] node35029;
	wire [4-1:0] node35032;
	wire [4-1:0] node35035;
	wire [4-1:0] node35036;
	wire [4-1:0] node35037;
	wire [4-1:0] node35038;
	wire [4-1:0] node35039;
	wire [4-1:0] node35040;
	wire [4-1:0] node35044;
	wire [4-1:0] node35046;
	wire [4-1:0] node35050;
	wire [4-1:0] node35052;
	wire [4-1:0] node35053;
	wire [4-1:0] node35054;
	wire [4-1:0] node35057;
	wire [4-1:0] node35061;
	wire [4-1:0] node35062;
	wire [4-1:0] node35063;
	wire [4-1:0] node35064;
	wire [4-1:0] node35067;
	wire [4-1:0] node35071;
	wire [4-1:0] node35073;
	wire [4-1:0] node35076;
	wire [4-1:0] node35077;
	wire [4-1:0] node35078;
	wire [4-1:0] node35079;
	wire [4-1:0] node35080;
	wire [4-1:0] node35083;
	wire [4-1:0] node35086;
	wire [4-1:0] node35087;
	wire [4-1:0] node35089;
	wire [4-1:0] node35092;
	wire [4-1:0] node35093;
	wire [4-1:0] node35097;
	wire [4-1:0] node35098;
	wire [4-1:0] node35101;
	wire [4-1:0] node35104;
	wire [4-1:0] node35105;
	wire [4-1:0] node35106;
	wire [4-1:0] node35109;
	wire [4-1:0] node35112;
	wire [4-1:0] node35113;
	wire [4-1:0] node35116;
	wire [4-1:0] node35119;
	wire [4-1:0] node35120;
	wire [4-1:0] node35121;
	wire [4-1:0] node35122;
	wire [4-1:0] node35123;
	wire [4-1:0] node35127;
	wire [4-1:0] node35128;
	wire [4-1:0] node35133;
	wire [4-1:0] node35134;
	wire [4-1:0] node35135;
	wire [4-1:0] node35136;
	wire [4-1:0] node35140;
	wire [4-1:0] node35141;
	wire [4-1:0] node35146;
	wire [4-1:0] node35147;
	wire [4-1:0] node35148;
	wire [4-1:0] node35149;
	wire [4-1:0] node35153;
	wire [4-1:0] node35154;
	wire [4-1:0] node35158;
	wire [4-1:0] node35159;

	assign outp = (inp[3]) ? node19848 : node1;
		assign node1 = (inp[6]) ? node12083 : node2;
			assign node2 = (inp[14]) ? node5980 : node3;
				assign node3 = (inp[8]) ? node2949 : node4;
					assign node4 = (inp[2]) ? node1460 : node5;
						assign node5 = (inp[13]) ? node733 : node6;
							assign node6 = (inp[1]) ? node366 : node7;
								assign node7 = (inp[12]) ? node195 : node8;
									assign node8 = (inp[7]) ? node96 : node9;
										assign node9 = (inp[4]) ? node45 : node10;
											assign node10 = (inp[11]) ? node24 : node11;
												assign node11 = (inp[15]) ? node19 : node12;
													assign node12 = (inp[10]) ? node16 : node13;
														assign node13 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node16 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node19 = (inp[10]) ? node21 : 4'b0001;
														assign node21 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node24 = (inp[5]) ? node38 : node25;
													assign node25 = (inp[9]) ? node31 : node26;
														assign node26 = (inp[15]) ? node28 : 4'b0001;
															assign node28 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node31 = (inp[10]) ? node35 : node32;
															assign node32 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node35 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node38 = (inp[10]) ? node40 : 4'b0000;
														assign node40 = (inp[9]) ? node42 : 4'b0000;
															assign node42 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node45 = (inp[15]) ? node61 : node46;
												assign node46 = (inp[11]) ? 4'b0001 : node47;
													assign node47 = (inp[10]) ? node53 : node48;
														assign node48 = (inp[9]) ? 4'b0001 : node49;
															assign node49 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node53 = (inp[9]) ? 4'b0000 : node54;
															assign node54 = (inp[0]) ? node56 : 4'b0001;
																assign node56 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node61 = (inp[5]) ? node83 : node62;
													assign node62 = (inp[11]) ? node70 : node63;
														assign node63 = (inp[0]) ? 4'b0010 : node64;
															assign node64 = (inp[10]) ? 4'b0010 : node65;
																assign node65 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node70 = (inp[9]) ? node76 : node71;
															assign node71 = (inp[10]) ? 4'b0011 : node72;
																assign node72 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node76 = (inp[0]) ? node80 : node77;
																assign node77 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node80 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node83 = (inp[0]) ? node91 : node84;
														assign node84 = (inp[11]) ? 4'b0111 : node85;
															assign node85 = (inp[10]) ? 4'b0110 : node86;
																assign node86 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node91 = (inp[11]) ? node93 : 4'b0111;
															assign node93 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node96 = (inp[15]) ? node154 : node97;
											assign node97 = (inp[11]) ? node127 : node98;
												assign node98 = (inp[0]) ? node116 : node99;
													assign node99 = (inp[10]) ? 4'b0011 : node100;
														assign node100 = (inp[4]) ? node108 : node101;
															assign node101 = (inp[5]) ? node105 : node102;
																assign node102 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node105 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node108 = (inp[9]) ? node112 : node109;
																assign node109 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node112 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node116 = (inp[9]) ? node120 : node117;
														assign node117 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node120 = (inp[10]) ? 4'b0010 : node121;
															assign node121 = (inp[4]) ? 4'b0011 : node122;
																assign node122 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node127 = (inp[10]) ? node137 : node128;
													assign node128 = (inp[0]) ? 4'b0011 : node129;
														assign node129 = (inp[9]) ? node131 : 4'b0010;
															assign node131 = (inp[4]) ? 4'b0011 : node132;
																assign node132 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node137 = (inp[5]) ? node145 : node138;
														assign node138 = (inp[4]) ? 4'b0010 : node139;
															assign node139 = (inp[9]) ? 4'b0011 : node140;
																assign node140 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node145 = (inp[0]) ? 4'b0011 : node146;
															assign node146 = (inp[4]) ? node150 : node147;
																assign node147 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node150 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node154 = (inp[4]) ? node172 : node155;
												assign node155 = (inp[9]) ? node165 : node156;
													assign node156 = (inp[5]) ? 4'b0111 : node157;
														assign node157 = (inp[10]) ? node159 : 4'b0110;
															assign node159 = (inp[0]) ? node161 : 4'b0111;
																assign node161 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node165 = (inp[5]) ? 4'b0110 : node166;
														assign node166 = (inp[10]) ? node168 : 4'b0111;
															assign node168 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node172 = (inp[9]) ? node182 : node173;
													assign node173 = (inp[11]) ? 4'b0001 : node174;
														assign node174 = (inp[10]) ? node178 : node175;
															assign node175 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node178 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node182 = (inp[0]) ? node190 : node183;
														assign node183 = (inp[5]) ? 4'b0001 : node184;
															assign node184 = (inp[11]) ? 4'b0000 : node185;
																assign node185 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node190 = (inp[10]) ? node192 : 4'b0000;
															assign node192 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node195 = (inp[7]) ? node261 : node196;
										assign node196 = (inp[4]) ? node216 : node197;
											assign node197 = (inp[9]) ? node205 : node198;
												assign node198 = (inp[10]) ? 4'b0011 : node199;
													assign node199 = (inp[0]) ? node201 : 4'b0010;
														assign node201 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node205 = (inp[10]) ? node211 : node206;
													assign node206 = (inp[11]) ? node208 : 4'b0011;
														assign node208 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node211 = (inp[11]) ? node213 : 4'b0010;
														assign node213 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node216 = (inp[15]) ? node234 : node217;
												assign node217 = (inp[9]) ? node227 : node218;
													assign node218 = (inp[11]) ? 4'b0110 : node219;
														assign node219 = (inp[5]) ? node221 : 4'b0111;
															assign node221 = (inp[10]) ? 4'b0110 : node222;
																assign node222 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node227 = (inp[0]) ? 4'b0111 : node228;
														assign node228 = (inp[10]) ? 4'b0110 : node229;
															assign node229 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node234 = (inp[11]) ? node244 : node235;
													assign node235 = (inp[5]) ? 4'b0000 : node236;
														assign node236 = (inp[9]) ? 4'b0001 : node237;
															assign node237 = (inp[10]) ? 4'b0000 : node238;
																assign node238 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node244 = (inp[10]) ? node256 : node245;
														assign node245 = (inp[9]) ? node251 : node246;
															assign node246 = (inp[5]) ? node248 : 4'b0001;
																assign node248 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node251 = (inp[5]) ? node253 : 4'b0000;
																assign node253 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node256 = (inp[0]) ? node258 : 4'b0001;
															assign node258 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node261 = (inp[15]) ? node313 : node262;
											assign node262 = (inp[11]) ? node284 : node263;
												assign node263 = (inp[4]) ? node275 : node264;
													assign node264 = (inp[5]) ? 4'b0101 : node265;
														assign node265 = (inp[9]) ? 4'b0001 : node266;
															assign node266 = (inp[0]) ? node270 : node267;
																assign node267 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node270 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node275 = (inp[5]) ? node279 : node276;
														assign node276 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node279 = (inp[9]) ? node281 : 4'b0000;
															assign node281 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node284 = (inp[0]) ? node304 : node285;
													assign node285 = (inp[5]) ? node293 : node286;
														assign node286 = (inp[4]) ? node288 : 4'b0001;
															assign node288 = (inp[9]) ? node290 : 4'b0101;
																assign node290 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node293 = (inp[4]) ? node299 : node294;
															assign node294 = (inp[9]) ? 4'b0101 : node295;
																assign node295 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node299 = (inp[9]) ? 4'b0001 : node300;
																assign node300 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node304 = (inp[9]) ? 4'b0001 : node305;
														assign node305 = (inp[5]) ? node309 : node306;
															assign node306 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node309 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node313 = (inp[4]) ? node339 : node314;
												assign node314 = (inp[5]) ? node328 : node315;
													assign node315 = (inp[0]) ? node323 : node316;
														assign node316 = (inp[9]) ? node318 : 4'b0101;
															assign node318 = (inp[10]) ? node320 : 4'b0101;
																assign node320 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node323 = (inp[10]) ? node325 : 4'b0100;
															assign node325 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node328 = (inp[9]) ? node330 : 4'b0000;
														assign node330 = (inp[0]) ? node332 : 4'b0001;
															assign node332 = (inp[11]) ? node336 : node333;
																assign node333 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node336 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node339 = (inp[5]) ? node357 : node340;
													assign node340 = (inp[10]) ? node346 : node341;
														assign node341 = (inp[0]) ? 4'b0111 : node342;
															assign node342 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node346 = (inp[9]) ? node352 : node347;
															assign node347 = (inp[0]) ? node349 : 4'b0110;
																assign node349 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node352 = (inp[11]) ? node354 : 4'b0111;
																assign node354 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node357 = (inp[0]) ? node359 : 4'b0111;
														assign node359 = (inp[10]) ? node363 : node360;
															assign node360 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node363 = (inp[9]) ? 4'b0111 : 4'b0110;
								assign node366 = (inp[5]) ? node560 : node367;
									assign node367 = (inp[12]) ? node449 : node368;
										assign node368 = (inp[15]) ? node404 : node369;
											assign node369 = (inp[7]) ? node387 : node370;
												assign node370 = (inp[10]) ? node382 : node371;
													assign node371 = (inp[9]) ? node377 : node372;
														assign node372 = (inp[11]) ? node374 : 4'b0000;
															assign node374 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node377 = (inp[0]) ? node379 : 4'b0001;
															assign node379 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node382 = (inp[9]) ? node384 : 4'b0001;
														assign node384 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node387 = (inp[0]) ? node395 : node388;
													assign node388 = (inp[10]) ? node392 : node389;
														assign node389 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node392 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node395 = (inp[9]) ? 4'b0010 : node396;
														assign node396 = (inp[11]) ? node400 : node397;
															assign node397 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node400 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node404 = (inp[7]) ? node422 : node405;
												assign node405 = (inp[4]) ? node413 : node406;
													assign node406 = (inp[9]) ? node408 : 4'b0001;
														assign node408 = (inp[0]) ? node410 : 4'b0000;
															assign node410 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node413 = (inp[9]) ? node417 : node414;
														assign node414 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node417 = (inp[10]) ? node419 : 4'b0110;
															assign node419 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node422 = (inp[4]) ? node432 : node423;
													assign node423 = (inp[11]) ? node425 : 4'b0111;
														assign node425 = (inp[0]) ? node427 : 4'b0110;
															assign node427 = (inp[10]) ? 4'b0111 : node428;
																assign node428 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node432 = (inp[9]) ? node442 : node433;
														assign node433 = (inp[10]) ? node437 : node434;
															assign node434 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node437 = (inp[0]) ? node439 : 4'b0000;
																assign node439 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node442 = (inp[10]) ? 4'b0001 : node443;
															assign node443 = (inp[11]) ? node445 : 4'b0000;
																assign node445 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node449 = (inp[7]) ? node503 : node450;
											assign node450 = (inp[15]) ? node476 : node451;
												assign node451 = (inp[4]) ? node465 : node452;
													assign node452 = (inp[11]) ? node460 : node453;
														assign node453 = (inp[9]) ? node457 : node454;
															assign node454 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node457 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node460 = (inp[9]) ? node462 : 4'b0010;
															assign node462 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node465 = (inp[9]) ? node471 : node466;
														assign node466 = (inp[11]) ? 4'b0111 : node467;
															assign node467 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node471 = (inp[10]) ? 4'b0111 : node472;
															assign node472 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node476 = (inp[4]) ? node492 : node477;
													assign node477 = (inp[0]) ? node485 : node478;
														assign node478 = (inp[9]) ? node480 : 4'b0011;
															assign node480 = (inp[10]) ? node482 : 4'b0011;
																assign node482 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node485 = (inp[10]) ? node489 : node486;
															assign node486 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node489 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node492 = (inp[11]) ? node498 : node493;
														assign node493 = (inp[10]) ? node495 : 4'b0001;
															assign node495 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node498 = (inp[0]) ? 4'b0000 : node499;
															assign node499 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node503 = (inp[15]) ? node529 : node504;
												assign node504 = (inp[4]) ? node518 : node505;
													assign node505 = (inp[10]) ? 4'b0101 : node506;
														assign node506 = (inp[9]) ? node512 : node507;
															assign node507 = (inp[11]) ? 4'b0100 : node508;
																assign node508 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node512 = (inp[11]) ? 4'b0101 : node513;
																assign node513 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node518 = (inp[9]) ? 4'b0000 : node519;
														assign node519 = (inp[10]) ? node523 : node520;
															assign node520 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node523 = (inp[11]) ? node525 : 4'b0001;
																assign node525 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node529 = (inp[4]) ? node543 : node530;
													assign node530 = (inp[9]) ? node536 : node531;
														assign node531 = (inp[11]) ? 4'b0000 : node532;
															assign node532 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node536 = (inp[11]) ? node540 : node537;
															assign node537 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node540 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node543 = (inp[10]) ? node553 : node544;
														assign node544 = (inp[9]) ? node548 : node545;
															assign node545 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node548 = (inp[0]) ? 4'b0110 : node549;
																assign node549 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node553 = (inp[9]) ? 4'b0111 : node554;
															assign node554 = (inp[11]) ? 4'b0110 : node555;
																assign node555 = (inp[0]) ? 4'b0110 : 4'b0111;
									assign node560 = (inp[12]) ? node636 : node561;
										assign node561 = (inp[7]) ? node599 : node562;
											assign node562 = (inp[15]) ? node584 : node563;
												assign node563 = (inp[9]) ? node575 : node564;
													assign node564 = (inp[0]) ? node566 : 4'b0100;
														assign node566 = (inp[10]) ? node570 : node567;
															assign node567 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node570 = (inp[4]) ? 4'b0100 : node571;
																assign node571 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node575 = (inp[11]) ? node581 : node576;
														assign node576 = (inp[0]) ? 4'b0101 : node577;
															assign node577 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node581 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node584 = (inp[4]) ? node594 : node585;
													assign node585 = (inp[10]) ? node587 : 4'b0101;
														assign node587 = (inp[11]) ? 4'b0100 : node588;
															assign node588 = (inp[0]) ? 4'b0101 : node589;
																assign node589 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node594 = (inp[10]) ? node596 : 4'b0110;
														assign node596 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node599 = (inp[15]) ? node613 : node600;
												assign node600 = (inp[9]) ? node602 : 4'b0110;
													assign node602 = (inp[11]) ? node608 : node603;
														assign node603 = (inp[10]) ? node605 : 4'b0110;
															assign node605 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node608 = (inp[10]) ? node610 : 4'b0111;
															assign node610 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node613 = (inp[4]) ? node623 : node614;
													assign node614 = (inp[10]) ? node618 : node615;
														assign node615 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node618 = (inp[9]) ? node620 : 4'b0011;
															assign node620 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node623 = (inp[11]) ? node625 : 4'b0101;
														assign node625 = (inp[0]) ? node631 : node626;
															assign node626 = (inp[9]) ? node628 : 4'b0101;
																assign node628 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node631 = (inp[9]) ? 4'b0101 : node632;
																assign node632 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node636 = (inp[7]) ? node700 : node637;
											assign node637 = (inp[15]) ? node669 : node638;
												assign node638 = (inp[4]) ? node652 : node639;
													assign node639 = (inp[9]) ? node647 : node640;
														assign node640 = (inp[10]) ? node642 : 4'b0111;
															assign node642 = (inp[11]) ? node644 : 4'b0110;
																assign node644 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node647 = (inp[10]) ? node649 : 4'b0110;
															assign node649 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node652 = (inp[0]) ? node660 : node653;
														assign node653 = (inp[9]) ? node657 : node654;
															assign node654 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node657 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node660 = (inp[9]) ? node662 : 4'b0011;
															assign node662 = (inp[11]) ? node666 : node663;
																assign node663 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node666 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node669 = (inp[4]) ? node685 : node670;
													assign node670 = (inp[0]) ? node676 : node671;
														assign node671 = (inp[9]) ? node673 : 4'b0110;
															assign node673 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node676 = (inp[11]) ? node678 : 4'b0111;
															assign node678 = (inp[9]) ? node682 : node679;
																assign node679 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node682 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node685 = (inp[10]) ? node691 : node686;
														assign node686 = (inp[9]) ? node688 : 4'b0101;
															assign node688 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node691 = (inp[9]) ? node697 : node692;
															assign node692 = (inp[0]) ? 4'b0100 : node693;
																assign node693 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node697 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node700 = (inp[4]) ? node722 : node701;
												assign node701 = (inp[15]) ? node703 : 4'b0100;
													assign node703 = (inp[0]) ? node709 : node704;
														assign node704 = (inp[11]) ? node706 : 4'b0001;
															assign node706 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node709 = (inp[11]) ? node717 : node710;
															assign node710 = (inp[9]) ? node714 : node711;
																assign node711 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node714 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node717 = (inp[9]) ? 4'b0000 : node718;
																assign node718 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node722 = (inp[15]) ? 4'b0010 : node723;
													assign node723 = (inp[0]) ? node725 : 4'b0000;
														assign node725 = (inp[9]) ? node729 : node726;
															assign node726 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node729 = (inp[10]) ? 4'b0000 : 4'b0001;
							assign node733 = (inp[1]) ? node1093 : node734;
								assign node734 = (inp[7]) ? node900 : node735;
									assign node735 = (inp[12]) ? node817 : node736;
										assign node736 = (inp[4]) ? node776 : node737;
											assign node737 = (inp[15]) ? node753 : node738;
												assign node738 = (inp[10]) ? node748 : node739;
													assign node739 = (inp[0]) ? node743 : node740;
														assign node740 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node743 = (inp[11]) ? node745 : 4'b0101;
															assign node745 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node748 = (inp[9]) ? 4'b0100 : node749;
														assign node749 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node753 = (inp[0]) ? node765 : node754;
													assign node754 = (inp[11]) ? node760 : node755;
														assign node755 = (inp[10]) ? node757 : 4'b0101;
															assign node757 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node760 = (inp[9]) ? 4'b0100 : node761;
															assign node761 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node765 = (inp[10]) ? node773 : node766;
														assign node766 = (inp[11]) ? node770 : node767;
															assign node767 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node770 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node773 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node776 = (inp[15]) ? node798 : node777;
												assign node777 = (inp[11]) ? node787 : node778;
													assign node778 = (inp[5]) ? 4'b0101 : node779;
														assign node779 = (inp[10]) ? node783 : node780;
															assign node780 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node783 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node787 = (inp[0]) ? node793 : node788;
														assign node788 = (inp[10]) ? node790 : 4'b0101;
															assign node790 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node793 = (inp[10]) ? 4'b0100 : node794;
															assign node794 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node798 = (inp[5]) ? node808 : node799;
													assign node799 = (inp[10]) ? node801 : 4'b0111;
														assign node801 = (inp[0]) ? node803 : 4'b0110;
															assign node803 = (inp[11]) ? node805 : 4'b0110;
																assign node805 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node808 = (inp[0]) ? 4'b0010 : node809;
														assign node809 = (inp[10]) ? node813 : node810;
															assign node810 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node813 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node817 = (inp[4]) ? node859 : node818;
											assign node818 = (inp[10]) ? node838 : node819;
												assign node819 = (inp[0]) ? node827 : node820;
													assign node820 = (inp[9]) ? node824 : node821;
														assign node821 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node824 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node827 = (inp[9]) ? node833 : node828;
														assign node828 = (inp[5]) ? 4'b0110 : node829;
															assign node829 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node833 = (inp[15]) ? node835 : 4'b0111;
															assign node835 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node838 = (inp[15]) ? node850 : node839;
													assign node839 = (inp[5]) ? 4'b0110 : node840;
														assign node840 = (inp[0]) ? node842 : 4'b0110;
															assign node842 = (inp[11]) ? node846 : node843;
																assign node843 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node846 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node850 = (inp[9]) ? node854 : node851;
														assign node851 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node854 = (inp[0]) ? node856 : 4'b0111;
															assign node856 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node859 = (inp[15]) ? node885 : node860;
												assign node860 = (inp[11]) ? node876 : node861;
													assign node861 = (inp[5]) ? 4'b0010 : node862;
														assign node862 = (inp[9]) ? node870 : node863;
															assign node863 = (inp[10]) ? node867 : node864;
																assign node864 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node867 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node870 = (inp[10]) ? 4'b0011 : node871;
																assign node871 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node876 = (inp[5]) ? 4'b0011 : node877;
														assign node877 = (inp[9]) ? node881 : node878;
															assign node878 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node881 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node885 = (inp[10]) ? node893 : node886;
													assign node886 = (inp[9]) ? node888 : 4'b0100;
														assign node888 = (inp[0]) ? 4'b0101 : node889;
															assign node889 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node893 = (inp[9]) ? node895 : 4'b0101;
														assign node895 = (inp[11]) ? 4'b0100 : node896;
															assign node896 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node900 = (inp[12]) ? node994 : node901;
										assign node901 = (inp[15]) ? node955 : node902;
											assign node902 = (inp[11]) ? node936 : node903;
												assign node903 = (inp[5]) ? node921 : node904;
													assign node904 = (inp[0]) ? node916 : node905;
														assign node905 = (inp[4]) ? node911 : node906;
															assign node906 = (inp[9]) ? node908 : 4'b0110;
																assign node908 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node911 = (inp[9]) ? 4'b0111 : node912;
																assign node912 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node916 = (inp[10]) ? node918 : 4'b0110;
															assign node918 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node921 = (inp[10]) ? node929 : node922;
														assign node922 = (inp[9]) ? node926 : node923;
															assign node923 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node926 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node929 = (inp[9]) ? 4'b0111 : node930;
															assign node930 = (inp[0]) ? node932 : 4'b0110;
																assign node932 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node936 = (inp[10]) ? node944 : node937;
													assign node937 = (inp[9]) ? 4'b0111 : node938;
														assign node938 = (inp[4]) ? node940 : 4'b0111;
															assign node940 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node944 = (inp[9]) ? node950 : node945;
														assign node945 = (inp[5]) ? 4'b0111 : node946;
															assign node946 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node950 = (inp[0]) ? node952 : 4'b0110;
															assign node952 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node955 = (inp[4]) ? node981 : node956;
												assign node956 = (inp[10]) ? node966 : node957;
													assign node957 = (inp[11]) ? node961 : node958;
														assign node958 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node961 = (inp[5]) ? node963 : 4'b0011;
															assign node963 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node966 = (inp[5]) ? node976 : node967;
														assign node967 = (inp[0]) ? node973 : node968;
															assign node968 = (inp[11]) ? 4'b0010 : node969;
																assign node969 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node973 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node976 = (inp[9]) ? node978 : 4'b0010;
															assign node978 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node981 = (inp[10]) ? node991 : node982;
													assign node982 = (inp[11]) ? node984 : 4'b0100;
														assign node984 = (inp[9]) ? 4'b0101 : node985;
															assign node985 = (inp[5]) ? node987 : 4'b0100;
																assign node987 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node991 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node994 = (inp[4]) ? node1056 : node995;
											assign node995 = (inp[0]) ? node1019 : node996;
												assign node996 = (inp[11]) ? node1008 : node997;
													assign node997 = (inp[15]) ? 4'b0000 : node998;
														assign node998 = (inp[5]) ? node1002 : node999;
															assign node999 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node1002 = (inp[9]) ? 4'b0001 : node1003;
																assign node1003 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node1008 = (inp[5]) ? node1012 : node1009;
														assign node1009 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node1012 = (inp[15]) ? node1016 : node1013;
															assign node1013 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node1016 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node1019 = (inp[5]) ? node1039 : node1020;
													assign node1020 = (inp[15]) ? node1026 : node1021;
														assign node1021 = (inp[9]) ? node1023 : 4'b0100;
															assign node1023 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node1026 = (inp[10]) ? node1032 : node1027;
															assign node1027 = (inp[9]) ? 4'b0001 : node1028;
																assign node1028 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node1032 = (inp[11]) ? node1036 : node1033;
																assign node1033 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node1036 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node1039 = (inp[15]) ? node1043 : node1040;
														assign node1040 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1043 = (inp[10]) ? node1049 : node1044;
															assign node1044 = (inp[9]) ? 4'b0100 : node1045;
																assign node1045 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node1049 = (inp[11]) ? node1053 : node1050;
																assign node1050 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node1053 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node1056 = (inp[15]) ? node1074 : node1057;
												assign node1057 = (inp[5]) ? node1065 : node1058;
													assign node1058 = (inp[9]) ? node1060 : 4'b0000;
														assign node1060 = (inp[10]) ? 4'b0001 : node1061;
															assign node1061 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node1065 = (inp[10]) ? node1069 : node1066;
														assign node1066 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node1069 = (inp[11]) ? 4'b0101 : node1070;
															assign node1070 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node1074 = (inp[5]) ? node1088 : node1075;
													assign node1075 = (inp[9]) ? node1083 : node1076;
														assign node1076 = (inp[10]) ? 4'b0010 : node1077;
															assign node1077 = (inp[0]) ? 4'b0011 : node1078;
																assign node1078 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1083 = (inp[10]) ? node1085 : 4'b0010;
															assign node1085 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1088 = (inp[10]) ? 4'b0011 : node1089;
														assign node1089 = (inp[9]) ? 4'b0011 : 4'b0010;
								assign node1093 = (inp[5]) ? node1283 : node1094;
									assign node1094 = (inp[12]) ? node1172 : node1095;
										assign node1095 = (inp[7]) ? node1135 : node1096;
											assign node1096 = (inp[4]) ? node1118 : node1097;
												assign node1097 = (inp[9]) ? node1103 : node1098;
													assign node1098 = (inp[0]) ? 4'b0101 : node1099;
														assign node1099 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node1103 = (inp[10]) ? node1109 : node1104;
														assign node1104 = (inp[0]) ? node1106 : 4'b0101;
															assign node1106 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node1109 = (inp[11]) ? node1113 : node1110;
															assign node1110 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1113 = (inp[15]) ? 4'b0100 : node1114;
																assign node1114 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node1118 = (inp[15]) ? node1126 : node1119;
													assign node1119 = (inp[0]) ? 4'b0101 : node1120;
														assign node1120 = (inp[9]) ? node1122 : 4'b0100;
															assign node1122 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1126 = (inp[9]) ? node1130 : node1127;
														assign node1127 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1130 = (inp[10]) ? node1132 : 4'b0011;
															assign node1132 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node1135 = (inp[15]) ? node1153 : node1136;
												assign node1136 = (inp[9]) ? node1146 : node1137;
													assign node1137 = (inp[10]) ? node1141 : node1138;
														assign node1138 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1141 = (inp[11]) ? node1143 : 4'b0111;
															assign node1143 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1146 = (inp[10]) ? 4'b0110 : node1147;
														assign node1147 = (inp[0]) ? node1149 : 4'b0111;
															assign node1149 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node1153 = (inp[4]) ? node1167 : node1154;
													assign node1154 = (inp[10]) ? node1158 : node1155;
														assign node1155 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1158 = (inp[11]) ? node1160 : 4'b0010;
															assign node1160 = (inp[0]) ? node1164 : node1161;
																assign node1161 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node1164 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node1167 = (inp[0]) ? node1169 : 4'b0101;
														assign node1169 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node1172 = (inp[7]) ? node1220 : node1173;
											assign node1173 = (inp[15]) ? node1199 : node1174;
												assign node1174 = (inp[4]) ? node1184 : node1175;
													assign node1175 = (inp[9]) ? node1177 : 4'b0110;
														assign node1177 = (inp[10]) ? node1179 : 4'b0110;
															assign node1179 = (inp[11]) ? node1181 : 4'b0111;
																assign node1181 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1184 = (inp[11]) ? node1194 : node1185;
														assign node1185 = (inp[0]) ? 4'b0010 : node1186;
															assign node1186 = (inp[10]) ? node1190 : node1187;
																assign node1187 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node1190 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node1194 = (inp[10]) ? node1196 : 4'b0011;
															assign node1196 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node1199 = (inp[4]) ? node1211 : node1200;
													assign node1200 = (inp[9]) ? node1206 : node1201;
														assign node1201 = (inp[10]) ? 4'b0110 : node1202;
															assign node1202 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1206 = (inp[0]) ? node1208 : 4'b0111;
															assign node1208 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node1211 = (inp[10]) ? node1213 : 4'b0100;
														assign node1213 = (inp[9]) ? node1217 : node1214;
															assign node1214 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node1217 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node1220 = (inp[15]) ? node1252 : node1221;
												assign node1221 = (inp[4]) ? node1237 : node1222;
													assign node1222 = (inp[0]) ? node1230 : node1223;
														assign node1223 = (inp[10]) ? node1227 : node1224;
															assign node1224 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node1227 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node1230 = (inp[11]) ? 4'b0001 : node1231;
															assign node1231 = (inp[10]) ? 4'b0001 : node1232;
																assign node1232 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node1237 = (inp[9]) ? node1243 : node1238;
														assign node1238 = (inp[10]) ? 4'b0101 : node1239;
															assign node1239 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node1243 = (inp[10]) ? node1247 : node1244;
															assign node1244 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node1247 = (inp[0]) ? node1249 : 4'b0100;
																assign node1249 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1252 = (inp[4]) ? node1268 : node1253;
													assign node1253 = (inp[11]) ? node1259 : node1254;
														assign node1254 = (inp[0]) ? 4'b0100 : node1255;
															assign node1255 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node1259 = (inp[0]) ? node1261 : 4'b0101;
															assign node1261 = (inp[9]) ? node1265 : node1262;
																assign node1262 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node1265 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1268 = (inp[10]) ? node1274 : node1269;
														assign node1269 = (inp[9]) ? node1271 : 4'b0010;
															assign node1271 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1274 = (inp[11]) ? node1276 : 4'b0011;
															assign node1276 = (inp[0]) ? node1280 : node1277;
																assign node1277 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node1280 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node1283 = (inp[7]) ? node1375 : node1284;
										assign node1284 = (inp[12]) ? node1322 : node1285;
											assign node1285 = (inp[0]) ? node1305 : node1286;
												assign node1286 = (inp[10]) ? node1294 : node1287;
													assign node1287 = (inp[9]) ? node1291 : node1288;
														assign node1288 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node1291 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node1294 = (inp[4]) ? 4'b0001 : node1295;
														assign node1295 = (inp[9]) ? node1301 : node1296;
															assign node1296 = (inp[15]) ? 4'b0001 : node1297;
																assign node1297 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node1301 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node1305 = (inp[15]) ? node1317 : node1306;
													assign node1306 = (inp[9]) ? 4'b0001 : node1307;
														assign node1307 = (inp[11]) ? node1311 : node1308;
															assign node1308 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node1311 = (inp[4]) ? node1313 : 4'b0000;
																assign node1313 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node1317 = (inp[10]) ? 4'b0010 : node1318;
														assign node1318 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node1322 = (inp[4]) ? node1354 : node1323;
												assign node1323 = (inp[0]) ? node1339 : node1324;
													assign node1324 = (inp[10]) ? node1334 : node1325;
														assign node1325 = (inp[9]) ? node1331 : node1326;
															assign node1326 = (inp[15]) ? 4'b0011 : node1327;
																assign node1327 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node1331 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node1334 = (inp[15]) ? 4'b0011 : node1335;
															assign node1335 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1339 = (inp[11]) ? node1347 : node1340;
														assign node1340 = (inp[10]) ? node1342 : 4'b0010;
															assign node1342 = (inp[9]) ? 4'b0011 : node1343;
																assign node1343 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node1347 = (inp[15]) ? 4'b0010 : node1348;
															assign node1348 = (inp[9]) ? node1350 : 4'b0010;
																assign node1350 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node1354 = (inp[15]) ? node1366 : node1355;
													assign node1355 = (inp[9]) ? node1361 : node1356;
														assign node1356 = (inp[0]) ? 4'b0111 : node1357;
															assign node1357 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node1361 = (inp[11]) ? node1363 : 4'b0110;
															assign node1363 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node1366 = (inp[9]) ? 4'b0001 : node1367;
														assign node1367 = (inp[10]) ? node1369 : 4'b0000;
															assign node1369 = (inp[0]) ? node1371 : 4'b0001;
																assign node1371 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node1375 = (inp[12]) ? node1423 : node1376;
											assign node1376 = (inp[15]) ? node1404 : node1377;
												assign node1377 = (inp[4]) ? node1391 : node1378;
													assign node1378 = (inp[11]) ? 4'b0011 : node1379;
														assign node1379 = (inp[0]) ? node1385 : node1380;
															assign node1380 = (inp[9]) ? node1382 : 4'b0010;
																assign node1382 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node1385 = (inp[10]) ? node1387 : 4'b0011;
																assign node1387 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node1391 = (inp[9]) ? node1399 : node1392;
														assign node1392 = (inp[0]) ? node1394 : 4'b0010;
															assign node1394 = (inp[11]) ? node1396 : 4'b0011;
																assign node1396 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node1399 = (inp[10]) ? 4'b0010 : node1400;
															assign node1400 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node1404 = (inp[4]) ? node1412 : node1405;
													assign node1405 = (inp[10]) ? node1407 : 4'b0110;
														assign node1407 = (inp[9]) ? 4'b0111 : node1408;
															assign node1408 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node1412 = (inp[0]) ? node1418 : node1413;
														assign node1413 = (inp[10]) ? 4'b0000 : node1414;
															assign node1414 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1418 = (inp[10]) ? node1420 : 4'b0001;
															assign node1420 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1423 = (inp[4]) ? node1443 : node1424;
												assign node1424 = (inp[15]) ? node1436 : node1425;
													assign node1425 = (inp[0]) ? 4'b0000 : node1426;
														assign node1426 = (inp[11]) ? node1432 : node1427;
															assign node1427 = (inp[10]) ? 4'b0001 : node1428;
																assign node1428 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node1432 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node1436 = (inp[10]) ? node1438 : 4'b0101;
														assign node1438 = (inp[11]) ? node1440 : 4'b0100;
															assign node1440 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node1443 = (inp[15]) ? node1451 : node1444;
													assign node1444 = (inp[9]) ? 4'b0100 : node1445;
														assign node1445 = (inp[10]) ? node1447 : 4'b0100;
															assign node1447 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node1451 = (inp[10]) ? node1453 : 4'b0110;
														assign node1453 = (inp[9]) ? node1457 : node1454;
															assign node1454 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1457 = (inp[11]) ? 4'b0110 : 4'b0111;
						assign node1460 = (inp[13]) ? node2182 : node1461;
							assign node1461 = (inp[1]) ? node1813 : node1462;
								assign node1462 = (inp[12]) ? node1634 : node1463;
									assign node1463 = (inp[7]) ? node1539 : node1464;
										assign node1464 = (inp[15]) ? node1512 : node1465;
											assign node1465 = (inp[10]) ? node1481 : node1466;
												assign node1466 = (inp[11]) ? node1476 : node1467;
													assign node1467 = (inp[5]) ? 4'b0101 : node1468;
														assign node1468 = (inp[4]) ? node1472 : node1469;
															assign node1469 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node1472 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1476 = (inp[4]) ? 4'b0101 : node1477;
														assign node1477 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node1481 = (inp[9]) ? node1497 : node1482;
													assign node1482 = (inp[5]) ? node1488 : node1483;
														assign node1483 = (inp[11]) ? node1485 : 4'b0100;
															assign node1485 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node1488 = (inp[0]) ? node1492 : node1489;
															assign node1489 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node1492 = (inp[4]) ? 4'b0101 : node1493;
																assign node1493 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node1497 = (inp[5]) ? node1505 : node1498;
														assign node1498 = (inp[11]) ? node1500 : 4'b0100;
															assign node1500 = (inp[4]) ? node1502 : 4'b0101;
																assign node1502 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1505 = (inp[11]) ? 4'b0100 : node1506;
															assign node1506 = (inp[0]) ? 4'b0100 : node1507;
																assign node1507 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node1512 = (inp[4]) ? node1528 : node1513;
												assign node1513 = (inp[0]) ? node1521 : node1514;
													assign node1514 = (inp[10]) ? node1518 : node1515;
														assign node1515 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node1518 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1521 = (inp[9]) ? node1523 : 4'b0101;
														assign node1523 = (inp[11]) ? node1525 : 4'b0100;
															assign node1525 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node1528 = (inp[5]) ? node1532 : node1529;
													assign node1529 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node1532 = (inp[10]) ? 4'b0011 : node1533;
														assign node1533 = (inp[9]) ? 4'b0011 : node1534;
															assign node1534 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node1539 = (inp[15]) ? node1597 : node1540;
											assign node1540 = (inp[5]) ? node1572 : node1541;
												assign node1541 = (inp[11]) ? node1553 : node1542;
													assign node1542 = (inp[0]) ? node1544 : 4'b0110;
														assign node1544 = (inp[4]) ? node1546 : 4'b0111;
															assign node1546 = (inp[10]) ? node1550 : node1547;
																assign node1547 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node1550 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node1553 = (inp[0]) ? node1563 : node1554;
														assign node1554 = (inp[9]) ? node1556 : 4'b0111;
															assign node1556 = (inp[10]) ? node1560 : node1557;
																assign node1557 = (inp[4]) ? 4'b0110 : 4'b0111;
																assign node1560 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node1563 = (inp[4]) ? node1565 : 4'b0110;
															assign node1565 = (inp[10]) ? node1569 : node1566;
																assign node1566 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node1569 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node1572 = (inp[0]) ? node1588 : node1573;
													assign node1573 = (inp[9]) ? node1579 : node1574;
														assign node1574 = (inp[10]) ? node1576 : 4'b0111;
															assign node1576 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node1579 = (inp[11]) ? 4'b0110 : node1580;
															assign node1580 = (inp[4]) ? node1584 : node1581;
																assign node1581 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node1584 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node1588 = (inp[10]) ? 4'b0111 : node1589;
														assign node1589 = (inp[9]) ? node1591 : 4'b0111;
															assign node1591 = (inp[11]) ? node1593 : 4'b0110;
																assign node1593 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node1597 = (inp[4]) ? node1613 : node1598;
												assign node1598 = (inp[11]) ? node1600 : 4'b0011;
													assign node1600 = (inp[0]) ? node1602 : 4'b0010;
														assign node1602 = (inp[5]) ? node1608 : node1603;
															assign node1603 = (inp[10]) ? 4'b0011 : node1604;
																assign node1604 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node1608 = (inp[10]) ? 4'b0010 : node1609;
																assign node1609 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node1613 = (inp[9]) ? node1619 : node1614;
													assign node1614 = (inp[10]) ? node1616 : 4'b0100;
														assign node1616 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node1619 = (inp[5]) ? node1631 : node1620;
														assign node1620 = (inp[10]) ? node1626 : node1621;
															assign node1621 = (inp[11]) ? 4'b0101 : node1622;
																assign node1622 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1626 = (inp[0]) ? 4'b0100 : node1627;
																assign node1627 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node1631 = (inp[11]) ? 4'b0101 : 4'b0100;
									assign node1634 = (inp[7]) ? node1724 : node1635;
										assign node1635 = (inp[15]) ? node1681 : node1636;
											assign node1636 = (inp[4]) ? node1652 : node1637;
												assign node1637 = (inp[0]) ? node1643 : node1638;
													assign node1638 = (inp[10]) ? node1640 : 4'b0110;
														assign node1640 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node1643 = (inp[5]) ? 4'b0111 : node1644;
														assign node1644 = (inp[9]) ? node1648 : node1645;
															assign node1645 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1648 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node1652 = (inp[11]) ? node1664 : node1653;
													assign node1653 = (inp[0]) ? node1661 : node1654;
														assign node1654 = (inp[9]) ? 4'b0011 : node1655;
															assign node1655 = (inp[5]) ? node1657 : 4'b0010;
																assign node1657 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1661 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node1664 = (inp[5]) ? node1674 : node1665;
														assign node1665 = (inp[0]) ? node1667 : 4'b0011;
															assign node1667 = (inp[10]) ? node1671 : node1668;
																assign node1668 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node1671 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node1674 = (inp[0]) ? 4'b0011 : node1675;
															assign node1675 = (inp[10]) ? node1677 : 4'b0010;
																assign node1677 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node1681 = (inp[4]) ? node1701 : node1682;
												assign node1682 = (inp[9]) ? node1692 : node1683;
													assign node1683 = (inp[10]) ? node1687 : node1684;
														assign node1684 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1687 = (inp[11]) ? node1689 : 4'b0111;
															assign node1689 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1692 = (inp[10]) ? node1696 : node1693;
														assign node1693 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1696 = (inp[0]) ? node1698 : 4'b0110;
															assign node1698 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node1701 = (inp[11]) ? node1713 : node1702;
													assign node1702 = (inp[5]) ? 4'b0100 : node1703;
														assign node1703 = (inp[0]) ? 4'b0100 : node1704;
															assign node1704 = (inp[10]) ? node1708 : node1705;
																assign node1705 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node1708 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node1713 = (inp[9]) ? node1717 : node1714;
														assign node1714 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node1717 = (inp[10]) ? node1721 : node1718;
															assign node1718 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1721 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node1724 = (inp[15]) ? node1770 : node1725;
											assign node1725 = (inp[10]) ? node1745 : node1726;
												assign node1726 = (inp[4]) ? node1736 : node1727;
													assign node1727 = (inp[5]) ? 4'b0001 : node1728;
														assign node1728 = (inp[9]) ? node1732 : node1729;
															assign node1729 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1732 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node1736 = (inp[5]) ? node1740 : node1737;
														assign node1737 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node1740 = (inp[9]) ? node1742 : 4'b0100;
															assign node1742 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1745 = (inp[5]) ? node1763 : node1746;
													assign node1746 = (inp[4]) ? node1756 : node1747;
														assign node1747 = (inp[11]) ? 4'b0101 : node1748;
															assign node1748 = (inp[9]) ? node1752 : node1749;
																assign node1749 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node1752 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node1756 = (inp[11]) ? node1760 : node1757;
															assign node1757 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node1760 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node1763 = (inp[4]) ? 4'b0100 : node1764;
														assign node1764 = (inp[9]) ? 4'b0000 : node1765;
															assign node1765 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1770 = (inp[4]) ? node1798 : node1771;
												assign node1771 = (inp[5]) ? node1787 : node1772;
													assign node1772 = (inp[11]) ? node1778 : node1773;
														assign node1773 = (inp[10]) ? node1775 : 4'b0000;
															assign node1775 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1778 = (inp[9]) ? node1780 : 4'b0001;
															assign node1780 = (inp[10]) ? node1784 : node1781;
																assign node1781 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node1784 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node1787 = (inp[11]) ? node1793 : node1788;
														assign node1788 = (inp[9]) ? 4'b0100 : node1789;
															assign node1789 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node1793 = (inp[10]) ? 4'b0101 : node1794;
															assign node1794 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node1798 = (inp[5]) ? node1806 : node1799;
													assign node1799 = (inp[9]) ? 4'b0011 : node1800;
														assign node1800 = (inp[10]) ? 4'b0010 : node1801;
															assign node1801 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1806 = (inp[9]) ? node1808 : 4'b0011;
														assign node1808 = (inp[0]) ? node1810 : 4'b0010;
															assign node1810 = (inp[11]) ? 4'b0011 : 4'b0010;
								assign node1813 = (inp[5]) ? node1997 : node1814;
									assign node1814 = (inp[4]) ? node1906 : node1815;
										assign node1815 = (inp[7]) ? node1857 : node1816;
											assign node1816 = (inp[12]) ? node1830 : node1817;
												assign node1817 = (inp[15]) ? node1823 : node1818;
													assign node1818 = (inp[9]) ? node1820 : 4'b0100;
														assign node1820 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1823 = (inp[9]) ? node1825 : 4'b0101;
														assign node1825 = (inp[10]) ? node1827 : 4'b0100;
															assign node1827 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1830 = (inp[11]) ? node1846 : node1831;
													assign node1831 = (inp[15]) ? node1833 : 4'b0110;
														assign node1833 = (inp[0]) ? node1839 : node1834;
															assign node1834 = (inp[9]) ? node1836 : 4'b0110;
																assign node1836 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node1839 = (inp[10]) ? node1843 : node1840;
																assign node1840 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node1843 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node1846 = (inp[9]) ? 4'b0111 : node1847;
														assign node1847 = (inp[0]) ? 4'b0111 : node1848;
															assign node1848 = (inp[10]) ? node1852 : node1849;
																assign node1849 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node1852 = (inp[15]) ? 4'b0111 : 4'b0110;
											assign node1857 = (inp[12]) ? node1885 : node1858;
												assign node1858 = (inp[15]) ? node1866 : node1859;
													assign node1859 = (inp[0]) ? 4'b0110 : node1860;
														assign node1860 = (inp[9]) ? 4'b0110 : node1861;
															assign node1861 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node1866 = (inp[11]) ? node1872 : node1867;
														assign node1867 = (inp[0]) ? node1869 : 4'b0010;
															assign node1869 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1872 = (inp[9]) ? node1880 : node1873;
															assign node1873 = (inp[0]) ? node1877 : node1874;
																assign node1874 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node1877 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node1880 = (inp[0]) ? 4'b0011 : node1881;
																assign node1881 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node1885 = (inp[15]) ? node1895 : node1886;
													assign node1886 = (inp[0]) ? node1888 : 4'b0001;
														assign node1888 = (inp[11]) ? node1892 : node1889;
															assign node1889 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node1892 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node1895 = (inp[9]) ? node1901 : node1896;
														assign node1896 = (inp[10]) ? node1898 : 4'b0101;
															assign node1898 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node1901 = (inp[10]) ? node1903 : 4'b0100;
															assign node1903 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node1906 = (inp[15]) ? node1952 : node1907;
											assign node1907 = (inp[12]) ? node1933 : node1908;
												assign node1908 = (inp[7]) ? node1922 : node1909;
													assign node1909 = (inp[10]) ? node1919 : node1910;
														assign node1910 = (inp[0]) ? node1912 : 4'b0100;
															assign node1912 = (inp[11]) ? node1916 : node1913;
																assign node1913 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node1916 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node1919 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node1922 = (inp[10]) ? node1924 : 4'b0111;
														assign node1924 = (inp[0]) ? node1926 : 4'b0111;
															assign node1926 = (inp[11]) ? node1930 : node1927;
																assign node1927 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node1930 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node1933 = (inp[7]) ? node1943 : node1934;
													assign node1934 = (inp[10]) ? 4'b0011 : node1935;
														assign node1935 = (inp[0]) ? 4'b0010 : node1936;
															assign node1936 = (inp[9]) ? node1938 : 4'b0011;
																assign node1938 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1943 = (inp[10]) ? node1945 : 4'b0101;
														assign node1945 = (inp[11]) ? node1947 : 4'b0101;
															assign node1947 = (inp[9]) ? node1949 : 4'b0100;
																assign node1949 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node1952 = (inp[9]) ? node1976 : node1953;
												assign node1953 = (inp[0]) ? node1965 : node1954;
													assign node1954 = (inp[10]) ? node1960 : node1955;
														assign node1955 = (inp[7]) ? 4'b0010 : node1956;
															assign node1956 = (inp[12]) ? 4'b0101 : 4'b0010;
														assign node1960 = (inp[7]) ? node1962 : 4'b0011;
															assign node1962 = (inp[12]) ? 4'b0011 : 4'b0101;
													assign node1965 = (inp[12]) ? node1971 : node1966;
														assign node1966 = (inp[10]) ? node1968 : 4'b0010;
															assign node1968 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1971 = (inp[7]) ? node1973 : 4'b0101;
															assign node1973 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node1976 = (inp[10]) ? node1984 : node1977;
													assign node1977 = (inp[12]) ? node1981 : node1978;
														assign node1978 = (inp[7]) ? 4'b0101 : 4'b0011;
														assign node1981 = (inp[7]) ? 4'b0011 : 4'b0100;
													assign node1984 = (inp[0]) ? node1990 : node1985;
														assign node1985 = (inp[7]) ? node1987 : 4'b0010;
															assign node1987 = (inp[12]) ? 4'b0010 : 4'b0100;
														assign node1990 = (inp[7]) ? node1994 : node1991;
															assign node1991 = (inp[11]) ? 4'b0011 : 4'b0101;
															assign node1994 = (inp[12]) ? 4'b0010 : 4'b0101;
									assign node1997 = (inp[12]) ? node2075 : node1998;
										assign node1998 = (inp[7]) ? node2024 : node1999;
											assign node1999 = (inp[4]) ? node2011 : node2000;
												assign node2000 = (inp[11]) ? node2006 : node2001;
													assign node2001 = (inp[10]) ? node2003 : 4'b0000;
														assign node2003 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node2006 = (inp[10]) ? node2008 : 4'b0001;
														assign node2008 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node2011 = (inp[15]) ? node2017 : node2012;
													assign node2012 = (inp[0]) ? node2014 : 4'b0000;
														assign node2014 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node2017 = (inp[9]) ? node2021 : node2018;
														assign node2018 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node2021 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node2024 = (inp[15]) ? node2056 : node2025;
												assign node2025 = (inp[4]) ? node2045 : node2026;
													assign node2026 = (inp[0]) ? node2032 : node2027;
														assign node2027 = (inp[10]) ? node2029 : 4'b0011;
															assign node2029 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node2032 = (inp[11]) ? node2038 : node2033;
															assign node2033 = (inp[10]) ? node2035 : 4'b0010;
																assign node2035 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node2038 = (inp[9]) ? node2042 : node2039;
																assign node2039 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node2042 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2045 = (inp[11]) ? node2049 : node2046;
														assign node2046 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node2049 = (inp[9]) ? 4'b0010 : node2050;
															assign node2050 = (inp[0]) ? 4'b0010 : node2051;
																assign node2051 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node2056 = (inp[4]) ? node2066 : node2057;
													assign node2057 = (inp[11]) ? node2059 : 4'b0110;
														assign node2059 = (inp[0]) ? 4'b0111 : node2060;
															assign node2060 = (inp[9]) ? node2062 : 4'b0110;
																assign node2062 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2066 = (inp[11]) ? node2068 : 4'b0001;
														assign node2068 = (inp[10]) ? node2070 : 4'b0000;
															assign node2070 = (inp[0]) ? node2072 : 4'b0001;
																assign node2072 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node2075 = (inp[7]) ? node2135 : node2076;
											assign node2076 = (inp[15]) ? node2106 : node2077;
												assign node2077 = (inp[4]) ? node2093 : node2078;
													assign node2078 = (inp[0]) ? node2088 : node2079;
														assign node2079 = (inp[9]) ? 4'b0011 : node2080;
															assign node2080 = (inp[11]) ? node2084 : node2081;
																assign node2081 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node2084 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node2088 = (inp[9]) ? 4'b0010 : node2089;
															assign node2089 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node2093 = (inp[11]) ? node2099 : node2094;
														assign node2094 = (inp[9]) ? 4'b0110 : node2095;
															assign node2095 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node2099 = (inp[10]) ? 4'b0111 : node2100;
															assign node2100 = (inp[9]) ? 4'b0110 : node2101;
																assign node2101 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node2106 = (inp[4]) ? node2120 : node2107;
													assign node2107 = (inp[11]) ? node2115 : node2108;
														assign node2108 = (inp[9]) ? node2112 : node2109;
															assign node2109 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2112 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node2115 = (inp[0]) ? 4'b0011 : node2116;
															assign node2116 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node2120 = (inp[9]) ? node2126 : node2121;
														assign node2121 = (inp[10]) ? 4'b0001 : node2122;
															assign node2122 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node2126 = (inp[10]) ? node2132 : node2127;
															assign node2127 = (inp[11]) ? node2129 : 4'b0001;
																assign node2129 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node2132 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node2135 = (inp[15]) ? node2161 : node2136;
												assign node2136 = (inp[4]) ? node2154 : node2137;
													assign node2137 = (inp[11]) ? node2143 : node2138;
														assign node2138 = (inp[0]) ? 4'b0000 : node2139;
															assign node2139 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node2143 = (inp[0]) ? node2149 : node2144;
															assign node2144 = (inp[10]) ? node2146 : 4'b0000;
																assign node2146 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node2149 = (inp[10]) ? 4'b0001 : node2150;
																assign node2150 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node2154 = (inp[11]) ? node2156 : 4'b0100;
														assign node2156 = (inp[10]) ? 4'b0101 : node2157;
															assign node2157 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node2161 = (inp[4]) ? node2175 : node2162;
													assign node2162 = (inp[9]) ? node2170 : node2163;
														assign node2163 = (inp[10]) ? node2167 : node2164;
															assign node2164 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node2167 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node2170 = (inp[10]) ? 4'b0100 : node2171;
															assign node2171 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node2175 = (inp[10]) ? node2179 : node2176;
														assign node2176 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node2179 = (inp[9]) ? 4'b0110 : 4'b0111;
							assign node2182 = (inp[5]) ? node2564 : node2183;
								assign node2183 = (inp[7]) ? node2373 : node2184;
									assign node2184 = (inp[12]) ? node2284 : node2185;
										assign node2185 = (inp[15]) ? node2223 : node2186;
											assign node2186 = (inp[0]) ? node2208 : node2187;
												assign node2187 = (inp[9]) ? node2201 : node2188;
													assign node2188 = (inp[11]) ? node2196 : node2189;
														assign node2189 = (inp[4]) ? node2193 : node2190;
															assign node2190 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node2193 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2196 = (inp[10]) ? node2198 : 4'b0000;
															assign node2198 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node2201 = (inp[11]) ? 4'b0001 : node2202;
														assign node2202 = (inp[1]) ? 4'b0000 : node2203;
															assign node2203 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node2208 = (inp[10]) ? node2216 : node2209;
													assign node2209 = (inp[9]) ? node2213 : node2210;
														assign node2210 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node2213 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node2216 = (inp[4]) ? node2220 : node2217;
														assign node2217 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node2220 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node2223 = (inp[4]) ? node2247 : node2224;
												assign node2224 = (inp[0]) ? node2236 : node2225;
													assign node2225 = (inp[9]) ? 4'b0000 : node2226;
														assign node2226 = (inp[1]) ? node2232 : node2227;
															assign node2227 = (inp[11]) ? 4'b0000 : node2228;
																assign node2228 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node2232 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2236 = (inp[11]) ? node2242 : node2237;
														assign node2237 = (inp[9]) ? node2239 : 4'b0001;
															assign node2239 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2242 = (inp[10]) ? node2244 : 4'b0000;
															assign node2244 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node2247 = (inp[1]) ? node2267 : node2248;
													assign node2248 = (inp[10]) ? node2258 : node2249;
														assign node2249 = (inp[11]) ? node2255 : node2250;
															assign node2250 = (inp[9]) ? 4'b0011 : node2251;
																assign node2251 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node2255 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node2258 = (inp[9]) ? node2264 : node2259;
															assign node2259 = (inp[0]) ? 4'b0010 : node2260;
																assign node2260 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node2264 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node2267 = (inp[9]) ? node2275 : node2268;
														assign node2268 = (inp[11]) ? node2270 : 4'b0111;
															assign node2270 = (inp[10]) ? 4'b0111 : node2271;
																assign node2271 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node2275 = (inp[0]) ? node2277 : 4'b0110;
															assign node2277 = (inp[10]) ? node2281 : node2278;
																assign node2278 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node2281 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node2284 = (inp[4]) ? node2328 : node2285;
											assign node2285 = (inp[11]) ? node2303 : node2286;
												assign node2286 = (inp[15]) ? node2298 : node2287;
													assign node2287 = (inp[10]) ? node2289 : 4'b0011;
														assign node2289 = (inp[0]) ? 4'b0010 : node2290;
															assign node2290 = (inp[9]) ? node2294 : node2291;
																assign node2291 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node2294 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node2298 = (inp[0]) ? node2300 : 4'b0011;
														assign node2300 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node2303 = (inp[15]) ? node2321 : node2304;
													assign node2304 = (inp[9]) ? node2314 : node2305;
														assign node2305 = (inp[0]) ? node2311 : node2306;
															assign node2306 = (inp[10]) ? node2308 : 4'b0010;
																assign node2308 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node2311 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node2314 = (inp[1]) ? node2318 : node2315;
															assign node2315 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2318 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2321 = (inp[10]) ? node2323 : 4'b0010;
														assign node2323 = (inp[0]) ? 4'b0010 : node2324;
															assign node2324 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node2328 = (inp[15]) ? node2350 : node2329;
												assign node2329 = (inp[1]) ? node2343 : node2330;
													assign node2330 = (inp[11]) ? 4'b0110 : node2331;
														assign node2331 = (inp[0]) ? node2337 : node2332;
															assign node2332 = (inp[9]) ? node2334 : 4'b0111;
																assign node2334 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2337 = (inp[9]) ? node2339 : 4'b0110;
																assign node2339 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2343 = (inp[10]) ? node2345 : 4'b0110;
														assign node2345 = (inp[0]) ? 4'b0110 : node2346;
															assign node2346 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node2350 = (inp[9]) ? node2362 : node2351;
													assign node2351 = (inp[11]) ? node2353 : 4'b0000;
														assign node2353 = (inp[1]) ? 4'b0000 : node2354;
															assign node2354 = (inp[0]) ? node2358 : node2355;
																assign node2355 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node2358 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2362 = (inp[0]) ? node2368 : node2363;
														assign node2363 = (inp[1]) ? node2365 : 4'b0001;
															assign node2365 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2368 = (inp[10]) ? node2370 : 4'b0000;
															assign node2370 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node2373 = (inp[12]) ? node2453 : node2374;
										assign node2374 = (inp[4]) ? node2414 : node2375;
											assign node2375 = (inp[15]) ? node2393 : node2376;
												assign node2376 = (inp[10]) ? node2384 : node2377;
													assign node2377 = (inp[0]) ? 4'b0010 : node2378;
														assign node2378 = (inp[11]) ? 4'b0011 : node2379;
															assign node2379 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node2384 = (inp[9]) ? node2390 : node2385;
														assign node2385 = (inp[0]) ? 4'b0010 : node2386;
															assign node2386 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node2390 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node2393 = (inp[11]) ? node2399 : node2394;
													assign node2394 = (inp[9]) ? 4'b0111 : node2395;
														assign node2395 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node2399 = (inp[0]) ? node2405 : node2400;
														assign node2400 = (inp[10]) ? node2402 : 4'b0110;
															assign node2402 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node2405 = (inp[10]) ? node2407 : 4'b0111;
															assign node2407 = (inp[1]) ? node2411 : node2408;
																assign node2408 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node2411 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node2414 = (inp[15]) ? node2436 : node2415;
												assign node2415 = (inp[0]) ? node2427 : node2416;
													assign node2416 = (inp[9]) ? node2422 : node2417;
														assign node2417 = (inp[10]) ? 4'b0011 : node2418;
															assign node2418 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node2422 = (inp[11]) ? node2424 : 4'b0010;
															assign node2424 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2427 = (inp[1]) ? 4'b0010 : node2428;
														assign node2428 = (inp[11]) ? 4'b0010 : node2429;
															assign node2429 = (inp[9]) ? node2431 : 4'b0011;
																assign node2431 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node2436 = (inp[10]) ? node2448 : node2437;
													assign node2437 = (inp[0]) ? node2441 : node2438;
														assign node2438 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node2441 = (inp[11]) ? 4'b0000 : node2442;
															assign node2442 = (inp[1]) ? 4'b0001 : node2443;
																assign node2443 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node2448 = (inp[0]) ? 4'b0001 : node2449;
														assign node2449 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node2453 = (inp[4]) ? node2515 : node2454;
											assign node2454 = (inp[10]) ? node2490 : node2455;
												assign node2455 = (inp[0]) ? node2471 : node2456;
													assign node2456 = (inp[9]) ? node2464 : node2457;
														assign node2457 = (inp[15]) ? node2461 : node2458;
															assign node2458 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node2461 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node2464 = (inp[1]) ? node2468 : node2465;
															assign node2465 = (inp[15]) ? 4'b0101 : 4'b0000;
															assign node2468 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2471 = (inp[9]) ? node2483 : node2472;
														assign node2472 = (inp[11]) ? node2478 : node2473;
															assign node2473 = (inp[1]) ? 4'b0100 : node2474;
																assign node2474 = (inp[15]) ? 4'b0100 : 4'b0001;
															assign node2478 = (inp[1]) ? node2480 : 4'b0000;
																assign node2480 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node2483 = (inp[11]) ? node2485 : 4'b0000;
															assign node2485 = (inp[15]) ? node2487 : 4'b0100;
																assign node2487 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node2490 = (inp[9]) ? node2502 : node2491;
													assign node2491 = (inp[1]) ? node2499 : node2492;
														assign node2492 = (inp[15]) ? node2494 : 4'b0000;
															assign node2494 = (inp[0]) ? node2496 : 4'b0101;
																assign node2496 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2499 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2502 = (inp[1]) ? node2508 : node2503;
														assign node2503 = (inp[11]) ? node2505 : 4'b0001;
															assign node2505 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node2508 = (inp[15]) ? node2512 : node2509;
															assign node2509 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node2512 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node2515 = (inp[15]) ? node2533 : node2516;
												assign node2516 = (inp[1]) ? node2522 : node2517;
													assign node2517 = (inp[10]) ? 4'b0100 : node2518;
														assign node2518 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node2522 = (inp[9]) ? node2526 : node2523;
														assign node2523 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node2526 = (inp[10]) ? node2528 : 4'b0001;
															assign node2528 = (inp[0]) ? 4'b0000 : node2529;
																assign node2529 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node2533 = (inp[9]) ? node2551 : node2534;
													assign node2534 = (inp[11]) ? node2542 : node2535;
														assign node2535 = (inp[10]) ? node2539 : node2536;
															assign node2536 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node2539 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node2542 = (inp[10]) ? node2548 : node2543;
															assign node2543 = (inp[1]) ? node2545 : 4'b0110;
																assign node2545 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node2548 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node2551 = (inp[11]) ? node2561 : node2552;
														assign node2552 = (inp[10]) ? node2556 : node2553;
															assign node2553 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node2556 = (inp[1]) ? 4'b0111 : node2557;
																assign node2557 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node2561 = (inp[10]) ? 4'b0110 : 4'b0111;
								assign node2564 = (inp[1]) ? node2740 : node2565;
									assign node2565 = (inp[7]) ? node2647 : node2566;
										assign node2566 = (inp[12]) ? node2602 : node2567;
											assign node2567 = (inp[15]) ? node2585 : node2568;
												assign node2568 = (inp[0]) ? node2570 : 4'b0000;
													assign node2570 = (inp[10]) ? node2576 : node2571;
														assign node2571 = (inp[9]) ? node2573 : 4'b0001;
															assign node2573 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node2576 = (inp[11]) ? node2582 : node2577;
															assign node2577 = (inp[4]) ? node2579 : 4'b0001;
																assign node2579 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node2582 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node2585 = (inp[4]) ? node2595 : node2586;
													assign node2586 = (inp[10]) ? node2590 : node2587;
														assign node2587 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node2590 = (inp[9]) ? node2592 : 4'b0001;
															assign node2592 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node2595 = (inp[0]) ? 4'b0111 : node2596;
														assign node2596 = (inp[10]) ? node2598 : 4'b0110;
															assign node2598 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node2602 = (inp[15]) ? node2624 : node2603;
												assign node2603 = (inp[4]) ? node2611 : node2604;
													assign node2604 = (inp[9]) ? node2606 : 4'b0010;
														assign node2606 = (inp[0]) ? 4'b0011 : node2607;
															assign node2607 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2611 = (inp[10]) ? node2617 : node2612;
														assign node2612 = (inp[9]) ? 4'b0111 : node2613;
															assign node2613 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node2617 = (inp[9]) ? node2619 : 4'b0111;
															assign node2619 = (inp[0]) ? node2621 : 4'b0110;
																assign node2621 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node2624 = (inp[4]) ? node2630 : node2625;
													assign node2625 = (inp[10]) ? node2627 : 4'b0011;
														assign node2627 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node2630 = (inp[11]) ? node2640 : node2631;
														assign node2631 = (inp[0]) ? node2633 : 4'b0001;
															assign node2633 = (inp[10]) ? node2637 : node2634;
																assign node2634 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node2637 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node2640 = (inp[10]) ? node2644 : node2641;
															assign node2641 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node2644 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node2647 = (inp[12]) ? node2687 : node2648;
											assign node2648 = (inp[15]) ? node2666 : node2649;
												assign node2649 = (inp[4]) ? node2661 : node2650;
													assign node2650 = (inp[9]) ? 4'b0010 : node2651;
														assign node2651 = (inp[10]) ? node2657 : node2652;
															assign node2652 = (inp[11]) ? 4'b0010 : node2653;
																assign node2653 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node2657 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node2661 = (inp[10]) ? node2663 : 4'b0011;
														assign node2663 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node2666 = (inp[4]) ? node2676 : node2667;
													assign node2667 = (inp[10]) ? node2669 : 4'b0111;
														assign node2669 = (inp[9]) ? 4'b0111 : node2670;
															assign node2670 = (inp[11]) ? 4'b0110 : node2671;
																assign node2671 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node2676 = (inp[10]) ? 4'b0001 : node2677;
														assign node2677 = (inp[11]) ? 4'b0000 : node2678;
															assign node2678 = (inp[0]) ? node2682 : node2679;
																assign node2679 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node2682 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node2687 = (inp[15]) ? node2713 : node2688;
												assign node2688 = (inp[4]) ? node2702 : node2689;
													assign node2689 = (inp[0]) ? node2697 : node2690;
														assign node2690 = (inp[10]) ? node2694 : node2691;
															assign node2691 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node2694 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node2697 = (inp[9]) ? node2699 : 4'b0101;
															assign node2699 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node2702 = (inp[10]) ? node2704 : 4'b0001;
														assign node2704 = (inp[9]) ? node2710 : node2705;
															assign node2705 = (inp[11]) ? node2707 : 4'b0001;
																assign node2707 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node2710 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node2713 = (inp[4]) ? node2721 : node2714;
													assign node2714 = (inp[10]) ? node2716 : 4'b0001;
														assign node2716 = (inp[9]) ? 4'b0000 : node2717;
															assign node2717 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node2721 = (inp[0]) ? node2727 : node2722;
														assign node2722 = (inp[11]) ? 4'b0110 : node2723;
															assign node2723 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node2727 = (inp[11]) ? node2733 : node2728;
															assign node2728 = (inp[9]) ? 4'b0110 : node2729;
																assign node2729 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node2733 = (inp[10]) ? node2737 : node2734;
																assign node2734 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node2737 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node2740 = (inp[12]) ? node2840 : node2741;
										assign node2741 = (inp[7]) ? node2789 : node2742;
											assign node2742 = (inp[15]) ? node2764 : node2743;
												assign node2743 = (inp[9]) ? node2753 : node2744;
													assign node2744 = (inp[4]) ? 4'b0101 : node2745;
														assign node2745 = (inp[11]) ? 4'b0100 : node2746;
															assign node2746 = (inp[0]) ? 4'b0101 : node2747;
																assign node2747 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node2753 = (inp[4]) ? node2755 : 4'b0100;
														assign node2755 = (inp[10]) ? node2759 : node2756;
															assign node2756 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node2759 = (inp[0]) ? node2761 : 4'b0100;
																assign node2761 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node2764 = (inp[4]) ? node2774 : node2765;
													assign node2765 = (inp[0]) ? 4'b0100 : node2766;
														assign node2766 = (inp[11]) ? node2768 : 4'b0101;
															assign node2768 = (inp[10]) ? 4'b0100 : node2769;
																assign node2769 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node2774 = (inp[11]) ? node2784 : node2775;
														assign node2775 = (inp[10]) ? 4'b0111 : node2776;
															assign node2776 = (inp[0]) ? node2780 : node2777;
																assign node2777 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node2780 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node2784 = (inp[10]) ? node2786 : 4'b0110;
															assign node2786 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node2789 = (inp[15]) ? node2817 : node2790;
												assign node2790 = (inp[9]) ? node2798 : node2791;
													assign node2791 = (inp[10]) ? node2795 : node2792;
														assign node2792 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node2795 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node2798 = (inp[4]) ? node2806 : node2799;
														assign node2799 = (inp[0]) ? 4'b0110 : node2800;
															assign node2800 = (inp[11]) ? 4'b0110 : node2801;
																assign node2801 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node2806 = (inp[10]) ? node2812 : node2807;
															assign node2807 = (inp[11]) ? node2809 : 4'b0110;
																assign node2809 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node2812 = (inp[0]) ? node2814 : 4'b0111;
																assign node2814 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node2817 = (inp[4]) ? node2823 : node2818;
													assign node2818 = (inp[9]) ? node2820 : 4'b0011;
														assign node2820 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2823 = (inp[11]) ? node2829 : node2824;
														assign node2824 = (inp[10]) ? node2826 : 4'b0101;
															assign node2826 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node2829 = (inp[0]) ? node2835 : node2830;
															assign node2830 = (inp[10]) ? node2832 : 4'b0101;
																assign node2832 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node2835 = (inp[9]) ? 4'b0100 : node2836;
																assign node2836 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node2840 = (inp[7]) ? node2888 : node2841;
											assign node2841 = (inp[15]) ? node2869 : node2842;
												assign node2842 = (inp[4]) ? node2854 : node2843;
													assign node2843 = (inp[10]) ? node2849 : node2844;
														assign node2844 = (inp[9]) ? node2846 : 4'b0110;
															assign node2846 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node2849 = (inp[11]) ? node2851 : 4'b0111;
															assign node2851 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node2854 = (inp[9]) ? node2862 : node2855;
														assign node2855 = (inp[10]) ? node2857 : 4'b0010;
															assign node2857 = (inp[11]) ? 4'b0011 : node2858;
																assign node2858 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node2862 = (inp[10]) ? node2864 : 4'b0011;
															assign node2864 = (inp[0]) ? 4'b0010 : node2865;
																assign node2865 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node2869 = (inp[4]) ? node2875 : node2870;
													assign node2870 = (inp[0]) ? 4'b0110 : node2871;
														assign node2871 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node2875 = (inp[11]) ? node2877 : 4'b0101;
														assign node2877 = (inp[0]) ? node2883 : node2878;
															assign node2878 = (inp[9]) ? node2880 : 4'b0101;
																assign node2880 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node2883 = (inp[9]) ? 4'b0100 : node2884;
																assign node2884 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node2888 = (inp[4]) ? node2920 : node2889;
												assign node2889 = (inp[15]) ? node2907 : node2890;
													assign node2890 = (inp[0]) ? node2898 : node2891;
														assign node2891 = (inp[9]) ? node2895 : node2892;
															assign node2892 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2895 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node2898 = (inp[11]) ? node2900 : 4'b0101;
															assign node2900 = (inp[9]) ? node2904 : node2901;
																assign node2901 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node2904 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node2907 = (inp[0]) ? node2915 : node2908;
														assign node2908 = (inp[9]) ? node2912 : node2909;
															assign node2909 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node2912 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2915 = (inp[10]) ? 4'b0000 : node2916;
															assign node2916 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node2920 = (inp[15]) ? node2936 : node2921;
													assign node2921 = (inp[0]) ? node2927 : node2922;
														assign node2922 = (inp[10]) ? node2924 : 4'b0000;
															assign node2924 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node2927 = (inp[11]) ? 4'b0001 : node2928;
															assign node2928 = (inp[9]) ? node2932 : node2929;
																assign node2929 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node2932 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2936 = (inp[10]) ? node2942 : node2937;
														assign node2937 = (inp[11]) ? node2939 : 4'b0010;
															assign node2939 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node2942 = (inp[9]) ? 4'b0011 : node2943;
															assign node2943 = (inp[0]) ? node2945 : 4'b0010;
																assign node2945 = (inp[11]) ? 4'b0011 : 4'b0010;
					assign node2949 = (inp[9]) ? node4473 : node2950;
						assign node2950 = (inp[13]) ? node3674 : node2951;
							assign node2951 = (inp[5]) ? node3289 : node2952;
								assign node2952 = (inp[10]) ? node3118 : node2953;
									assign node2953 = (inp[0]) ? node3041 : node2954;
										assign node2954 = (inp[2]) ? node2994 : node2955;
											assign node2955 = (inp[1]) ? node2977 : node2956;
												assign node2956 = (inp[7]) ? node2964 : node2957;
													assign node2957 = (inp[12]) ? node2961 : node2958;
														assign node2958 = (inp[4]) ? 4'b1010 : 4'b1000;
														assign node2961 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node2964 = (inp[11]) ? node2966 : 4'b1010;
														assign node2966 = (inp[15]) ? node2972 : node2967;
															assign node2967 = (inp[12]) ? node2969 : 4'b1000;
																assign node2969 = (inp[4]) ? 4'b1001 : 4'b1011;
															assign node2972 = (inp[12]) ? node2974 : 4'b1011;
																assign node2974 = (inp[4]) ? 4'b1101 : 4'b1111;
												assign node2977 = (inp[4]) ? node2991 : node2978;
													assign node2978 = (inp[12]) ? node2984 : node2979;
														assign node2979 = (inp[11]) ? node2981 : 4'b1100;
															assign node2981 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node2984 = (inp[7]) ? 4'b1011 : node2985;
															assign node2985 = (inp[11]) ? node2987 : 4'b1111;
																assign node2987 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node2991 = (inp[12]) ? 4'b1100 : 4'b1110;
											assign node2994 = (inp[7]) ? node3012 : node2995;
												assign node2995 = (inp[4]) ? node2999 : node2996;
													assign node2996 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node2999 = (inp[12]) ? node3001 : 4'b1111;
														assign node3001 = (inp[11]) ? node3009 : node3002;
															assign node3002 = (inp[1]) ? node3006 : node3003;
																assign node3003 = (inp[15]) ? 4'b1101 : 4'b1001;
																assign node3006 = (inp[15]) ? 4'b1001 : 4'b1100;
															assign node3009 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node3012 = (inp[1]) ? node3028 : node3013;
													assign node3013 = (inp[15]) ? node3021 : node3014;
														assign node3014 = (inp[4]) ? node3018 : node3015;
															assign node3015 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node3018 = (inp[12]) ? 4'b1100 : 4'b1111;
														assign node3021 = (inp[4]) ? node3025 : node3022;
															assign node3022 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node3025 = (inp[12]) ? 4'b1000 : 4'b1110;
													assign node3028 = (inp[15]) ? node3036 : node3029;
														assign node3029 = (inp[12]) ? 4'b1010 : node3030;
															assign node3030 = (inp[4]) ? node3032 : 4'b1001;
																assign node3032 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node3036 = (inp[4]) ? node3038 : 4'b1101;
															assign node3038 = (inp[12]) ? 4'b1100 : 4'b1010;
										assign node3041 = (inp[15]) ? node3081 : node3042;
											assign node3042 = (inp[4]) ? node3056 : node3043;
												assign node3043 = (inp[12]) ? node3053 : node3044;
													assign node3044 = (inp[2]) ? node3048 : node3045;
														assign node3045 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node3048 = (inp[1]) ? node3050 : 4'b1101;
															assign node3050 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3053 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node3056 = (inp[12]) ? node3066 : node3057;
													assign node3057 = (inp[2]) ? node3061 : node3058;
														assign node3058 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node3061 = (inp[1]) ? node3063 : 4'b1110;
															assign node3063 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node3066 = (inp[7]) ? node3076 : node3067;
														assign node3067 = (inp[11]) ? 4'b1001 : node3068;
															assign node3068 = (inp[2]) ? node3072 : node3069;
																assign node3069 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node3072 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node3076 = (inp[2]) ? node3078 : 4'b1101;
															assign node3078 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node3081 = (inp[11]) ? node3099 : node3082;
												assign node3082 = (inp[4]) ? node3090 : node3083;
													assign node3083 = (inp[12]) ? 4'b1011 : node3084;
														assign node3084 = (inp[2]) ? node3086 : 4'b1101;
															assign node3086 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3090 = (inp[12]) ? node3096 : node3091;
														assign node3091 = (inp[1]) ? node3093 : 4'b1110;
															assign node3093 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node3096 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node3099 = (inp[1]) ? node3109 : node3100;
													assign node3100 = (inp[7]) ? node3104 : node3101;
														assign node3101 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node3104 = (inp[2]) ? 4'b1000 : node3105;
															assign node3105 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node3109 = (inp[7]) ? node3113 : node3110;
														assign node3110 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node3113 = (inp[2]) ? 4'b1110 : node3114;
															assign node3114 = (inp[4]) ? 4'b1000 : 4'b1010;
									assign node3118 = (inp[0]) ? node3206 : node3119;
										assign node3119 = (inp[4]) ? node3165 : node3120;
											assign node3120 = (inp[12]) ? node3144 : node3121;
												assign node3121 = (inp[1]) ? node3133 : node3122;
													assign node3122 = (inp[2]) ? node3128 : node3123;
														assign node3123 = (inp[7]) ? node3125 : 4'b1001;
															assign node3125 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node3128 = (inp[15]) ? node3130 : 4'b1101;
															assign node3130 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3133 = (inp[15]) ? node3139 : node3134;
														assign node3134 = (inp[2]) ? node3136 : 4'b1101;
															assign node3136 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node3139 = (inp[2]) ? node3141 : 4'b1000;
															assign node3141 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node3144 = (inp[7]) ? node3156 : node3145;
													assign node3145 = (inp[15]) ? node3147 : 4'b1011;
														assign node3147 = (inp[11]) ? node3149 : 4'b1011;
															assign node3149 = (inp[1]) ? node3153 : node3150;
																assign node3150 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node3153 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node3156 = (inp[11]) ? node3158 : 4'b1011;
														assign node3158 = (inp[2]) ? 4'b1011 : node3159;
															assign node3159 = (inp[1]) ? 4'b1010 : node3160;
																assign node3160 = (inp[15]) ? 4'b1110 : 4'b1010;
											assign node3165 = (inp[12]) ? node3183 : node3166;
												assign node3166 = (inp[2]) ? node3172 : node3167;
													assign node3167 = (inp[1]) ? node3169 : 4'b1011;
														assign node3169 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node3172 = (inp[1]) ? node3174 : 4'b1110;
														assign node3174 = (inp[7]) ? node3178 : node3175;
															assign node3175 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node3178 = (inp[15]) ? node3180 : 4'b1010;
																assign node3180 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node3183 = (inp[7]) ? node3199 : node3184;
													assign node3184 = (inp[1]) ? 4'b1101 : node3185;
														assign node3185 = (inp[11]) ? node3193 : node3186;
															assign node3186 = (inp[2]) ? node3190 : node3187;
																assign node3187 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node3190 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node3193 = (inp[2]) ? node3195 : 4'b1101;
																assign node3195 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node3199 = (inp[2]) ? node3203 : node3200;
														assign node3200 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node3203 = (inp[1]) ? 4'b1101 : 4'b1000;
										assign node3206 = (inp[4]) ? node3248 : node3207;
											assign node3207 = (inp[12]) ? node3227 : node3208;
												assign node3208 = (inp[1]) ? node3216 : node3209;
													assign node3209 = (inp[2]) ? 4'b1100 : node3210;
														assign node3210 = (inp[7]) ? node3212 : 4'b1000;
															assign node3212 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node3216 = (inp[2]) ? node3222 : node3217;
														assign node3217 = (inp[11]) ? node3219 : 4'b1100;
															assign node3219 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node3222 = (inp[7]) ? node3224 : 4'b1001;
															assign node3224 = (inp[15]) ? 4'b1101 : 4'b1000;
												assign node3227 = (inp[15]) ? node3235 : node3228;
													assign node3228 = (inp[11]) ? 4'b1110 : node3229;
														assign node3229 = (inp[7]) ? 4'b1010 : node3230;
															assign node3230 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node3235 = (inp[2]) ? node3245 : node3236;
														assign node3236 = (inp[7]) ? node3240 : node3237;
															assign node3237 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node3240 = (inp[1]) ? 4'b1010 : node3241;
																assign node3241 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node3245 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node3248 = (inp[12]) ? node3268 : node3249;
												assign node3249 = (inp[1]) ? node3255 : node3250;
													assign node3250 = (inp[2]) ? node3252 : 4'b1010;
														assign node3252 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node3255 = (inp[2]) ? node3259 : node3256;
														assign node3256 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node3259 = (inp[11]) ? node3263 : node3260;
															assign node3260 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node3263 = (inp[15]) ? node3265 : 4'b1010;
																assign node3265 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node3268 = (inp[11]) ? node3276 : node3269;
													assign node3269 = (inp[15]) ? node3271 : 4'b1001;
														assign node3271 = (inp[7]) ? 4'b1001 : node3272;
															assign node3272 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node3276 = (inp[2]) ? node3282 : node3277;
														assign node3277 = (inp[1]) ? node3279 : 4'b1001;
															assign node3279 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node3282 = (inp[15]) ? node3286 : node3283;
															assign node3283 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node3286 = (inp[7]) ? 4'b1001 : 4'b1100;
								assign node3289 = (inp[0]) ? node3465 : node3290;
									assign node3290 = (inp[10]) ? node3396 : node3291;
										assign node3291 = (inp[11]) ? node3347 : node3292;
											assign node3292 = (inp[15]) ? node3320 : node3293;
												assign node3293 = (inp[7]) ? node3305 : node3294;
													assign node3294 = (inp[12]) ? node3302 : node3295;
														assign node3295 = (inp[4]) ? node3299 : node3296;
															assign node3296 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node3299 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node3302 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node3305 = (inp[2]) ? node3307 : 4'b1111;
														assign node3307 = (inp[1]) ? node3313 : node3308;
															assign node3308 = (inp[4]) ? 4'b1101 : node3309;
																assign node3309 = (inp[12]) ? 4'b1010 : 4'b1001;
															assign node3313 = (inp[4]) ? node3317 : node3314;
																assign node3314 = (inp[12]) ? 4'b1111 : 4'b1101;
																assign node3317 = (inp[12]) ? 4'b1001 : 4'b1111;
												assign node3320 = (inp[12]) ? node3334 : node3321;
													assign node3321 = (inp[4]) ? node3327 : node3322;
														assign node3322 = (inp[1]) ? node3324 : 4'b1001;
															assign node3324 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node3327 = (inp[2]) ? node3329 : 4'b1011;
															assign node3329 = (inp[7]) ? node3331 : 4'b1010;
																assign node3331 = (inp[1]) ? 4'b1010 : 4'b1111;
													assign node3334 = (inp[4]) ? node3340 : node3335;
														assign node3335 = (inp[1]) ? 4'b1111 : node3336;
															assign node3336 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node3340 = (inp[1]) ? node3344 : node3341;
															assign node3341 = (inp[7]) ? 4'b1001 : 4'b1100;
															assign node3344 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node3347 = (inp[7]) ? node3367 : node3348;
												assign node3348 = (inp[2]) ? node3358 : node3349;
													assign node3349 = (inp[1]) ? node3355 : node3350;
														assign node3350 = (inp[4]) ? 4'b1001 : node3351;
															assign node3351 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node3355 = (inp[15]) ? 4'b1010 : 4'b1100;
													assign node3358 = (inp[1]) ? node3360 : 4'b1110;
														assign node3360 = (inp[12]) ? node3364 : node3361;
															assign node3361 = (inp[4]) ? 4'b1010 : 4'b1001;
															assign node3364 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node3367 = (inp[15]) ? node3389 : node3368;
													assign node3368 = (inp[1]) ? node3376 : node3369;
														assign node3369 = (inp[12]) ? node3371 : 4'b1101;
															assign node3371 = (inp[4]) ? 4'b1100 : node3372;
																assign node3372 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node3376 = (inp[2]) ? node3384 : node3377;
															assign node3377 = (inp[4]) ? node3381 : node3378;
																assign node3378 = (inp[12]) ? 4'b1011 : 4'b1000;
																assign node3381 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node3384 = (inp[12]) ? 4'b1001 : node3385;
																assign node3385 = (inp[4]) ? 4'b1111 : 4'b1100;
													assign node3389 = (inp[1]) ? node3393 : node3390;
														assign node3390 = (inp[4]) ? 4'b1010 : 4'b1000;
														assign node3393 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node3396 = (inp[4]) ? node3442 : node3397;
											assign node3397 = (inp[12]) ? node3419 : node3398;
												assign node3398 = (inp[15]) ? node3408 : node3399;
													assign node3399 = (inp[1]) ? node3401 : 4'b1001;
														assign node3401 = (inp[2]) ? node3405 : node3402;
															assign node3402 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node3405 = (inp[11]) ? 4'b1101 : 4'b1001;
													assign node3408 = (inp[2]) ? node3414 : node3409;
														assign node3409 = (inp[7]) ? node3411 : 4'b1001;
															assign node3411 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node3414 = (inp[1]) ? 4'b1000 : node3415;
															assign node3415 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node3419 = (inp[1]) ? node3427 : node3420;
													assign node3420 = (inp[2]) ? node3422 : 4'b1011;
														assign node3422 = (inp[15]) ? 4'b1111 : node3423;
															assign node3423 = (inp[7]) ? 4'b1011 : 4'b1111;
													assign node3427 = (inp[11]) ? node3435 : node3428;
														assign node3428 = (inp[15]) ? 4'b1110 : node3429;
															assign node3429 = (inp[7]) ? node3431 : 4'b1010;
																assign node3431 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node3435 = (inp[2]) ? 4'b1011 : node3436;
															assign node3436 = (inp[15]) ? 4'b1111 : node3437;
																assign node3437 = (inp[7]) ? 4'b1010 : 4'b1110;
											assign node3442 = (inp[12]) ? node3452 : node3443;
												assign node3443 = (inp[11]) ? 4'b1110 : node3444;
													assign node3444 = (inp[15]) ? node3448 : node3445;
														assign node3445 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node3448 = (inp[7]) ? 4'b1011 : 4'b1111;
												assign node3452 = (inp[2]) ? node3460 : node3453;
													assign node3453 = (inp[1]) ? node3455 : 4'b1000;
														assign node3455 = (inp[11]) ? node3457 : 4'b1101;
															assign node3457 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node3460 = (inp[1]) ? node3462 : 4'b1101;
														assign node3462 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node3465 = (inp[10]) ? node3561 : node3466;
										assign node3466 = (inp[2]) ? node3512 : node3467;
											assign node3467 = (inp[1]) ? node3485 : node3468;
												assign node3468 = (inp[4]) ? node3476 : node3469;
													assign node3469 = (inp[12]) ? node3473 : node3470;
														assign node3470 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node3473 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node3476 = (inp[12]) ? 4'b1000 : node3477;
														assign node3477 = (inp[7]) ? 4'b1111 : node3478;
															assign node3478 = (inp[15]) ? node3480 : 4'b1010;
																assign node3480 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node3485 = (inp[4]) ? node3501 : node3486;
													assign node3486 = (inp[12]) ? node3492 : node3487;
														assign node3487 = (inp[7]) ? 4'b1101 : node3488;
															assign node3488 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node3492 = (inp[7]) ? node3498 : node3493;
															assign node3493 = (inp[15]) ? node3495 : 4'b1110;
																assign node3495 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node3498 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node3501 = (inp[12]) ? node3503 : 4'b1110;
														assign node3503 = (inp[7]) ? node3509 : node3504;
															assign node3504 = (inp[15]) ? node3506 : 4'b1101;
																assign node3506 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node3509 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node3512 = (inp[1]) ? node3534 : node3513;
												assign node3513 = (inp[7]) ? node3523 : node3514;
													assign node3514 = (inp[4]) ? node3518 : node3515;
														assign node3515 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node3518 = (inp[12]) ? 4'b1101 : node3519;
															assign node3519 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node3523 = (inp[12]) ? node3527 : node3524;
														assign node3524 = (inp[4]) ? 4'b1010 : 4'b1000;
														assign node3527 = (inp[4]) ? node3531 : node3528;
															assign node3528 = (inp[11]) ? 4'b1111 : 4'b1011;
															assign node3531 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node3534 = (inp[11]) ? node3550 : node3535;
													assign node3535 = (inp[15]) ? node3547 : node3536;
														assign node3536 = (inp[7]) ? node3542 : node3537;
															assign node3537 = (inp[12]) ? node3539 : 4'b1011;
																assign node3539 = (inp[4]) ? 4'b1000 : 4'b1010;
															assign node3542 = (inp[12]) ? node3544 : 4'b1110;
																assign node3544 = (inp[4]) ? 4'b1000 : 4'b1110;
														assign node3547 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node3550 = (inp[4]) ? node3558 : node3551;
														assign node3551 = (inp[12]) ? 4'b1011 : node3552;
															assign node3552 = (inp[7]) ? node3554 : 4'b1000;
																assign node3554 = (inp[15]) ? 4'b1000 : 4'b1101;
														assign node3558 = (inp[7]) ? 4'b1011 : 4'b1001;
										assign node3561 = (inp[7]) ? node3615 : node3562;
											assign node3562 = (inp[1]) ? node3584 : node3563;
												assign node3563 = (inp[2]) ? node3573 : node3564;
													assign node3564 = (inp[4]) ? node3568 : node3565;
														assign node3565 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node3568 = (inp[12]) ? 4'b1001 : node3569;
															assign node3569 = (inp[11]) ? 4'b1111 : 4'b1010;
													assign node3573 = (inp[4]) ? node3577 : node3574;
														assign node3574 = (inp[12]) ? 4'b1110 : 4'b1100;
														assign node3577 = (inp[12]) ? 4'b1100 : node3578;
															assign node3578 = (inp[15]) ? 4'b1010 : node3579;
																assign node3579 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node3584 = (inp[2]) ? node3602 : node3585;
													assign node3585 = (inp[15]) ? node3595 : node3586;
														assign node3586 = (inp[11]) ? 4'b1111 : node3587;
															assign node3587 = (inp[4]) ? node3591 : node3588;
																assign node3588 = (inp[12]) ? 4'b1111 : 4'b1100;
																assign node3591 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node3595 = (inp[4]) ? node3599 : node3596;
															assign node3596 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node3599 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node3602 = (inp[12]) ? node3608 : node3603;
														assign node3603 = (inp[4]) ? 4'b1111 : node3604;
															assign node3604 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node3608 = (inp[4]) ? 4'b1000 : node3609;
															assign node3609 = (inp[15]) ? 4'b1010 : node3610;
																assign node3610 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node3615 = (inp[15]) ? node3651 : node3616;
												assign node3616 = (inp[11]) ? node3634 : node3617;
													assign node3617 = (inp[4]) ? node3627 : node3618;
														assign node3618 = (inp[12]) ? 4'b1011 : node3619;
															assign node3619 = (inp[1]) ? node3623 : node3620;
																assign node3620 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node3623 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node3627 = (inp[12]) ? 4'b1101 : node3628;
															assign node3628 = (inp[1]) ? 4'b1111 : node3629;
																assign node3629 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node3634 = (inp[1]) ? node3646 : node3635;
														assign node3635 = (inp[12]) ? node3641 : node3636;
															assign node3636 = (inp[2]) ? 4'b1011 : node3637;
																assign node3637 = (inp[4]) ? 4'b1110 : 4'b1101;
															assign node3641 = (inp[4]) ? node3643 : 4'b1010;
																assign node3643 = (inp[2]) ? 4'b1100 : 4'b1001;
														assign node3646 = (inp[4]) ? 4'b1001 : node3647;
															assign node3647 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node3651 = (inp[12]) ? node3661 : node3652;
													assign node3652 = (inp[4]) ? node3656 : node3653;
														assign node3653 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node3656 = (inp[11]) ? 4'b1111 : node3657;
															assign node3657 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node3661 = (inp[4]) ? node3667 : node3662;
														assign node3662 = (inp[1]) ? 4'b1111 : node3663;
															assign node3663 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node3667 = (inp[2]) ? node3671 : node3668;
															assign node3668 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node3671 = (inp[1]) ? 4'b1000 : 4'b1100;
							assign node3674 = (inp[1]) ? node4066 : node3675;
								assign node3675 = (inp[2]) ? node3855 : node3676;
									assign node3676 = (inp[7]) ? node3760 : node3677;
										assign node3677 = (inp[4]) ? node3717 : node3678;
											assign node3678 = (inp[12]) ? node3700 : node3679;
												assign node3679 = (inp[5]) ? node3685 : node3680;
													assign node3680 = (inp[15]) ? node3682 : 4'b1001;
														assign node3682 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node3685 = (inp[0]) ? node3693 : node3686;
														assign node3686 = (inp[11]) ? node3688 : 4'b1000;
															assign node3688 = (inp[10]) ? node3690 : 4'b1001;
																assign node3690 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node3693 = (inp[11]) ? 4'b1000 : node3694;
															assign node3694 = (inp[10]) ? node3696 : 4'b1000;
																assign node3696 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node3700 = (inp[15]) ? node3710 : node3701;
													assign node3701 = (inp[5]) ? node3703 : 4'b1010;
														assign node3703 = (inp[0]) ? node3705 : 4'b1011;
															assign node3705 = (inp[10]) ? node3707 : 4'b1010;
																assign node3707 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node3710 = (inp[10]) ? node3712 : 4'b1011;
														assign node3712 = (inp[11]) ? 4'b1011 : node3713;
															assign node3713 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node3717 = (inp[12]) ? node3735 : node3718;
												assign node3718 = (inp[5]) ? node3724 : node3719;
													assign node3719 = (inp[11]) ? 4'b1011 : node3720;
														assign node3720 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node3724 = (inp[15]) ? node3728 : node3725;
														assign node3725 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node3728 = (inp[0]) ? node3732 : node3729;
															assign node3729 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node3732 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node3735 = (inp[5]) ? node3745 : node3736;
													assign node3736 = (inp[15]) ? 4'b1001 : node3737;
														assign node3737 = (inp[10]) ? 4'b1101 : node3738;
															assign node3738 = (inp[11]) ? node3740 : 4'b1100;
																assign node3740 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node3745 = (inp[0]) ? node3751 : node3746;
														assign node3746 = (inp[15]) ? 4'b1000 : node3747;
															assign node3747 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node3751 = (inp[15]) ? node3753 : 4'b1000;
															assign node3753 = (inp[10]) ? node3757 : node3754;
																assign node3754 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node3757 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node3760 = (inp[5]) ? node3816 : node3761;
											assign node3761 = (inp[15]) ? node3787 : node3762;
												assign node3762 = (inp[12]) ? node3774 : node3763;
													assign node3763 = (inp[4]) ? node3765 : 4'b1000;
														assign node3765 = (inp[11]) ? 4'b1011 : node3766;
															assign node3766 = (inp[0]) ? node3770 : node3767;
																assign node3767 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node3770 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node3774 = (inp[4]) ? node3780 : node3775;
														assign node3775 = (inp[0]) ? node3777 : 4'b1011;
															assign node3777 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node3780 = (inp[11]) ? 4'b1000 : node3781;
															assign node3781 = (inp[0]) ? 4'b1001 : node3782;
																assign node3782 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node3787 = (inp[10]) ? node3805 : node3788;
													assign node3788 = (inp[0]) ? node3794 : node3789;
														assign node3789 = (inp[12]) ? node3791 : 4'b1100;
															assign node3791 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node3794 = (inp[11]) ? node3802 : node3795;
															assign node3795 = (inp[4]) ? node3799 : node3796;
																assign node3796 = (inp[12]) ? 4'b1111 : 4'b1100;
																assign node3799 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node3802 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node3805 = (inp[11]) ? node3811 : node3806;
														assign node3806 = (inp[0]) ? node3808 : 4'b1101;
															assign node3808 = (inp[12]) ? 4'b1110 : 4'b1101;
														assign node3811 = (inp[4]) ? 4'b1011 : node3812;
															assign node3812 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node3816 = (inp[15]) ? node3836 : node3817;
												assign node3817 = (inp[11]) ? node3827 : node3818;
													assign node3818 = (inp[10]) ? node3824 : node3819;
														assign node3819 = (inp[12]) ? node3821 : 4'b1110;
															assign node3821 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node3824 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node3827 = (inp[12]) ? node3829 : 4'b1110;
														assign node3829 = (inp[0]) ? node3833 : node3830;
															assign node3830 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node3833 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node3836 = (inp[12]) ? node3846 : node3837;
													assign node3837 = (inp[4]) ? node3839 : 4'b1000;
														assign node3839 = (inp[10]) ? 4'b1010 : node3840;
															assign node3840 = (inp[11]) ? 4'b1010 : node3841;
																assign node3841 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node3846 = (inp[4]) ? 4'b1000 : node3847;
														assign node3847 = (inp[11]) ? 4'b1011 : node3848;
															assign node3848 = (inp[10]) ? node3850 : 4'b1011;
																assign node3850 = (inp[0]) ? 4'b1011 : 4'b1010;
									assign node3855 = (inp[7]) ? node3961 : node3856;
										assign node3856 = (inp[4]) ? node3902 : node3857;
											assign node3857 = (inp[12]) ? node3883 : node3858;
												assign node3858 = (inp[0]) ? node3868 : node3859;
													assign node3859 = (inp[11]) ? node3861 : 4'b1100;
														assign node3861 = (inp[5]) ? node3863 : 4'b1101;
															assign node3863 = (inp[10]) ? 4'b1100 : node3864;
																assign node3864 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node3868 = (inp[10]) ? node3870 : 4'b1101;
														assign node3870 = (inp[5]) ? node3876 : node3871;
															assign node3871 = (inp[15]) ? 4'b1101 : node3872;
																assign node3872 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node3876 = (inp[15]) ? node3880 : node3877;
																assign node3877 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node3880 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node3883 = (inp[15]) ? node3893 : node3884;
													assign node3884 = (inp[0]) ? node3886 : 4'b1111;
														assign node3886 = (inp[10]) ? node3890 : node3887;
															assign node3887 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node3890 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node3893 = (inp[11]) ? 4'b1110 : node3894;
														assign node3894 = (inp[5]) ? node3896 : 4'b1110;
															assign node3896 = (inp[0]) ? 4'b1111 : node3897;
																assign node3897 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node3902 = (inp[12]) ? node3934 : node3903;
												assign node3903 = (inp[15]) ? node3917 : node3904;
													assign node3904 = (inp[0]) ? node3912 : node3905;
														assign node3905 = (inp[10]) ? node3907 : 4'b1110;
															assign node3907 = (inp[5]) ? 4'b1111 : node3908;
																assign node3908 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node3912 = (inp[10]) ? node3914 : 4'b1111;
															assign node3914 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node3917 = (inp[5]) ? node3927 : node3918;
														assign node3918 = (inp[0]) ? 4'b1110 : node3919;
															assign node3919 = (inp[10]) ? node3923 : node3920;
																assign node3920 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node3923 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node3927 = (inp[11]) ? node3929 : 4'b1011;
															assign node3929 = (inp[10]) ? node3931 : 4'b1010;
																assign node3931 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node3934 = (inp[5]) ? node3944 : node3935;
													assign node3935 = (inp[15]) ? node3939 : node3936;
														assign node3936 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node3939 = (inp[10]) ? 4'b1101 : node3940;
															assign node3940 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node3944 = (inp[15]) ? node3954 : node3945;
														assign node3945 = (inp[0]) ? 4'b1101 : node3946;
															assign node3946 = (inp[11]) ? node3950 : node3947;
																assign node3947 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node3950 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node3954 = (inp[0]) ? node3956 : 4'b1100;
															assign node3956 = (inp[11]) ? 4'b1100 : node3957;
																assign node3957 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node3961 = (inp[5]) ? node4009 : node3962;
											assign node3962 = (inp[15]) ? node3986 : node3963;
												assign node3963 = (inp[4]) ? node3975 : node3964;
													assign node3964 = (inp[12]) ? node3968 : node3965;
														assign node3965 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node3968 = (inp[0]) ? node3972 : node3969;
															assign node3969 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node3972 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node3975 = (inp[12]) ? node3981 : node3976;
														assign node3976 = (inp[10]) ? node3978 : 4'b1110;
															assign node3978 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node3981 = (inp[11]) ? node3983 : 4'b1100;
															assign node3983 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node3986 = (inp[12]) ? node4000 : node3987;
													assign node3987 = (inp[4]) ? node3993 : node3988;
														assign node3988 = (inp[0]) ? 4'b1000 : node3989;
															assign node3989 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node3993 = (inp[11]) ? 4'b1110 : node3994;
															assign node3994 = (inp[10]) ? node3996 : 4'b1111;
																assign node3996 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node4000 = (inp[4]) ? node4004 : node4001;
														assign node4001 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node4004 = (inp[0]) ? 4'b1000 : node4005;
															assign node4005 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node4009 = (inp[15]) ? node4031 : node4010;
												assign node4010 = (inp[0]) ? node4016 : node4011;
													assign node4011 = (inp[11]) ? node4013 : 4'b1011;
														assign node4013 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node4016 = (inp[10]) ? node4022 : node4017;
														assign node4017 = (inp[12]) ? 4'b1101 : node4018;
															assign node4018 = (inp[11]) ? 4'b1011 : 4'b1001;
														assign node4022 = (inp[4]) ? node4028 : node4023;
															assign node4023 = (inp[12]) ? node4025 : 4'b1000;
																assign node4025 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node4028 = (inp[11]) ? 4'b1100 : 4'b1011;
												assign node4031 = (inp[0]) ? node4051 : node4032;
													assign node4032 = (inp[4]) ? node4042 : node4033;
														assign node4033 = (inp[12]) ? node4037 : node4034;
															assign node4034 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node4037 = (inp[10]) ? node4039 : 4'b1110;
																assign node4039 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node4042 = (inp[12]) ? node4044 : 4'b1110;
															assign node4044 = (inp[11]) ? node4048 : node4045;
																assign node4045 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node4048 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node4051 = (inp[10]) ? node4057 : node4052;
														assign node4052 = (inp[12]) ? 4'b1101 : node4053;
															assign node4053 = (inp[11]) ? 4'b1110 : 4'b1100;
														assign node4057 = (inp[12]) ? node4061 : node4058;
															assign node4058 = (inp[4]) ? 4'b1111 : 4'b1101;
															assign node4061 = (inp[11]) ? 4'b1110 : node4062;
																assign node4062 = (inp[4]) ? 4'b1101 : 4'b1111;
								assign node4066 = (inp[2]) ? node4272 : node4067;
									assign node4067 = (inp[7]) ? node4163 : node4068;
										assign node4068 = (inp[4]) ? node4108 : node4069;
											assign node4069 = (inp[12]) ? node4091 : node4070;
												assign node4070 = (inp[15]) ? node4086 : node4071;
													assign node4071 = (inp[5]) ? node4079 : node4072;
														assign node4072 = (inp[11]) ? node4074 : 4'b1101;
															assign node4074 = (inp[10]) ? node4076 : 4'b1101;
																assign node4076 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node4079 = (inp[10]) ? 4'b1100 : node4080;
															assign node4080 = (inp[11]) ? 4'b1101 : node4081;
																assign node4081 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node4086 = (inp[10]) ? node4088 : 4'b1100;
														assign node4088 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node4091 = (inp[0]) ? node4097 : node4092;
													assign node4092 = (inp[10]) ? node4094 : 4'b1111;
														assign node4094 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node4097 = (inp[10]) ? node4103 : node4098;
														assign node4098 = (inp[11]) ? node4100 : 4'b1110;
															assign node4100 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node4103 = (inp[15]) ? 4'b1111 : node4104;
															assign node4104 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node4108 = (inp[12]) ? node4132 : node4109;
												assign node4109 = (inp[15]) ? node4123 : node4110;
													assign node4110 = (inp[10]) ? 4'b1110 : node4111;
														assign node4111 = (inp[0]) ? node4117 : node4112;
															assign node4112 = (inp[5]) ? 4'b1111 : node4113;
																assign node4113 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node4117 = (inp[11]) ? 4'b1110 : node4118;
																assign node4118 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node4123 = (inp[5]) ? node4127 : node4124;
														assign node4124 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node4127 = (inp[10]) ? 4'b1010 : node4128;
															assign node4128 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node4132 = (inp[10]) ? node4148 : node4133;
													assign node4133 = (inp[15]) ? node4141 : node4134;
														assign node4134 = (inp[0]) ? node4138 : node4135;
															assign node4135 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node4138 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node4141 = (inp[5]) ? 4'b1100 : node4142;
															assign node4142 = (inp[0]) ? 4'b1100 : node4143;
																assign node4143 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node4148 = (inp[0]) ? node4154 : node4149;
														assign node4149 = (inp[11]) ? node4151 : 4'b1101;
															assign node4151 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node4154 = (inp[15]) ? node4158 : node4155;
															assign node4155 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node4158 = (inp[11]) ? 4'b1100 : node4159;
																assign node4159 = (inp[5]) ? 4'b1100 : 4'b1101;
										assign node4163 = (inp[4]) ? node4219 : node4164;
											assign node4164 = (inp[12]) ? node4204 : node4165;
												assign node4165 = (inp[10]) ? node4187 : node4166;
													assign node4166 = (inp[11]) ? node4180 : node4167;
														assign node4167 = (inp[0]) ? node4175 : node4168;
															assign node4168 = (inp[15]) ? node4172 : node4169;
																assign node4169 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node4172 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node4175 = (inp[5]) ? node4177 : 4'b1001;
																assign node4177 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node4180 = (inp[15]) ? 4'b1000 : node4181;
															assign node4181 = (inp[5]) ? 4'b1000 : node4182;
																assign node4182 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node4187 = (inp[0]) ? node4199 : node4188;
														assign node4188 = (inp[5]) ? node4194 : node4189;
															assign node4189 = (inp[15]) ? node4191 : 4'b1100;
																assign node4191 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node4194 = (inp[15]) ? node4196 : 4'b1001;
																assign node4196 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node4199 = (inp[15]) ? node4201 : 4'b1100;
															assign node4201 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node4204 = (inp[15]) ? node4214 : node4205;
													assign node4205 = (inp[5]) ? node4209 : node4206;
														assign node4206 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node4209 = (inp[10]) ? node4211 : 4'b1010;
															assign node4211 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node4214 = (inp[5]) ? 4'b1111 : node4215;
														assign node4215 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node4219 = (inp[12]) ? node4245 : node4220;
												assign node4220 = (inp[5]) ? node4232 : node4221;
													assign node4221 = (inp[10]) ? node4227 : node4222;
														assign node4222 = (inp[15]) ? 4'b1111 : node4223;
															assign node4223 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node4227 = (inp[0]) ? node4229 : 4'b1110;
															assign node4229 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node4232 = (inp[15]) ? node4238 : node4233;
														assign node4233 = (inp[0]) ? 4'b1011 : node4234;
															assign node4234 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node4238 = (inp[11]) ? node4242 : node4239;
															assign node4239 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node4242 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node4245 = (inp[5]) ? node4257 : node4246;
													assign node4246 = (inp[15]) ? 4'b1001 : node4247;
														assign node4247 = (inp[11]) ? node4249 : 4'b1100;
															assign node4249 = (inp[0]) ? node4253 : node4250;
																assign node4250 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node4253 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node4257 = (inp[11]) ? node4263 : node4258;
														assign node4258 = (inp[15]) ? node4260 : 4'b1101;
															assign node4260 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node4263 = (inp[15]) ? node4265 : 4'b1100;
															assign node4265 = (inp[10]) ? node4269 : node4266;
																assign node4266 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node4269 = (inp[0]) ? 4'b1100 : 4'b1101;
									assign node4272 = (inp[7]) ? node4362 : node4273;
										assign node4273 = (inp[4]) ? node4313 : node4274;
											assign node4274 = (inp[12]) ? node4290 : node4275;
												assign node4275 = (inp[0]) ? node4283 : node4276;
													assign node4276 = (inp[10]) ? node4278 : 4'b1001;
														assign node4278 = (inp[11]) ? 4'b1000 : node4279;
															assign node4279 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node4283 = (inp[15]) ? node4285 : 4'b1000;
														assign node4285 = (inp[10]) ? 4'b1001 : node4286;
															assign node4286 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node4290 = (inp[0]) ? node4302 : node4291;
													assign node4291 = (inp[10]) ? node4297 : node4292;
														assign node4292 = (inp[11]) ? 4'b1010 : node4293;
															assign node4293 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node4297 = (inp[11]) ? 4'b1011 : node4298;
															assign node4298 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node4302 = (inp[10]) ? node4308 : node4303;
														assign node4303 = (inp[15]) ? node4305 : 4'b1011;
															assign node4305 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node4308 = (inp[15]) ? node4310 : 4'b1010;
															assign node4310 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node4313 = (inp[12]) ? node4339 : node4314;
												assign node4314 = (inp[5]) ? node4326 : node4315;
													assign node4315 = (inp[0]) ? node4321 : node4316;
														assign node4316 = (inp[10]) ? 4'b1011 : node4317;
															assign node4317 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node4321 = (inp[10]) ? 4'b1010 : node4322;
															assign node4322 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node4326 = (inp[15]) ? node4334 : node4327;
														assign node4327 = (inp[0]) ? node4331 : node4328;
															assign node4328 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node4331 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node4334 = (inp[0]) ? node4336 : 4'b1111;
															assign node4336 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node4339 = (inp[5]) ? node4349 : node4340;
													assign node4340 = (inp[15]) ? node4344 : node4341;
														assign node4341 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node4344 = (inp[10]) ? node4346 : 4'b1001;
															assign node4346 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node4349 = (inp[0]) ? node4355 : node4350;
														assign node4350 = (inp[10]) ? node4352 : 4'b1000;
															assign node4352 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node4355 = (inp[10]) ? node4357 : 4'b1001;
															assign node4357 = (inp[11]) ? 4'b1000 : node4358;
																assign node4358 = (inp[15]) ? 4'b1001 : 4'b1000;
										assign node4362 = (inp[4]) ? node4424 : node4363;
											assign node4363 = (inp[12]) ? node4397 : node4364;
												assign node4364 = (inp[11]) ? node4378 : node4365;
													assign node4365 = (inp[15]) ? node4369 : node4366;
														assign node4366 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node4369 = (inp[5]) ? node4371 : 4'b1101;
															assign node4371 = (inp[10]) ? node4375 : node4372;
																assign node4372 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node4375 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node4378 = (inp[10]) ? node4386 : node4379;
														assign node4379 = (inp[15]) ? node4383 : node4380;
															assign node4380 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node4383 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node4386 = (inp[0]) ? node4390 : node4387;
															assign node4387 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node4390 = (inp[5]) ? node4394 : node4391;
																assign node4391 = (inp[15]) ? 4'b1101 : 4'b1001;
																assign node4394 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node4397 = (inp[5]) ? node4413 : node4398;
													assign node4398 = (inp[15]) ? node4406 : node4399;
														assign node4399 = (inp[0]) ? node4403 : node4400;
															assign node4400 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node4403 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node4406 = (inp[11]) ? 4'b1110 : node4407;
															assign node4407 = (inp[10]) ? 4'b1111 : node4408;
																assign node4408 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node4413 = (inp[15]) ? node4421 : node4414;
														assign node4414 = (inp[0]) ? node4416 : 4'b1111;
															assign node4416 = (inp[11]) ? node4418 : 4'b1111;
																assign node4418 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node4421 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node4424 = (inp[12]) ? node4450 : node4425;
												assign node4425 = (inp[15]) ? node4437 : node4426;
													assign node4426 = (inp[5]) ? node4430 : node4427;
														assign node4427 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node4430 = (inp[0]) ? 4'b1111 : node4431;
															assign node4431 = (inp[11]) ? node4433 : 4'b1110;
																assign node4433 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node4437 = (inp[5]) ? node4443 : node4438;
														assign node4438 = (inp[0]) ? node4440 : 4'b1011;
															assign node4440 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node4443 = (inp[10]) ? node4445 : 4'b1010;
															assign node4445 = (inp[11]) ? node4447 : 4'b1010;
																assign node4447 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node4450 = (inp[15]) ? node4462 : node4451;
													assign node4451 = (inp[5]) ? node4457 : node4452;
														assign node4452 = (inp[0]) ? 4'b1001 : node4453;
															assign node4453 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node4457 = (inp[0]) ? 4'b1000 : node4458;
															assign node4458 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node4462 = (inp[5]) ? node4470 : node4463;
														assign node4463 = (inp[11]) ? node4467 : node4464;
															assign node4464 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node4467 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node4470 = (inp[0]) ? 4'b1001 : 4'b1000;
						assign node4473 = (inp[15]) ? node5245 : node4474;
							assign node4474 = (inp[2]) ? node4858 : node4475;
								assign node4475 = (inp[1]) ? node4665 : node4476;
									assign node4476 = (inp[5]) ? node4562 : node4477;
										assign node4477 = (inp[4]) ? node4523 : node4478;
											assign node4478 = (inp[12]) ? node4498 : node4479;
												assign node4479 = (inp[0]) ? node4487 : node4480;
													assign node4480 = (inp[10]) ? node4482 : 4'b1000;
														assign node4482 = (inp[13]) ? node4484 : 4'b1001;
															assign node4484 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node4487 = (inp[10]) ? node4493 : node4488;
														assign node4488 = (inp[11]) ? node4490 : 4'b1001;
															assign node4490 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node4493 = (inp[13]) ? node4495 : 4'b1000;
															assign node4495 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4498 = (inp[0]) ? node4514 : node4499;
													assign node4499 = (inp[13]) ? node4509 : node4500;
														assign node4500 = (inp[10]) ? node4506 : node4501;
															assign node4501 = (inp[11]) ? node4503 : 4'b1010;
																assign node4503 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node4506 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node4509 = (inp[7]) ? node4511 : 4'b1010;
															assign node4511 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node4514 = (inp[13]) ? node4516 : 4'b1011;
														assign node4516 = (inp[10]) ? 4'b1011 : node4517;
															assign node4517 = (inp[11]) ? 4'b1010 : node4518;
																assign node4518 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node4523 = (inp[12]) ? node4541 : node4524;
												assign node4524 = (inp[0]) ? node4532 : node4525;
													assign node4525 = (inp[10]) ? node4527 : 4'b1010;
														assign node4527 = (inp[13]) ? node4529 : 4'b1011;
															assign node4529 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node4532 = (inp[11]) ? node4534 : 4'b1011;
														assign node4534 = (inp[10]) ? node4538 : node4535;
															assign node4535 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node4538 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node4541 = (inp[7]) ? node4553 : node4542;
													assign node4542 = (inp[13]) ? node4544 : 4'b1100;
														assign node4544 = (inp[11]) ? 4'b1101 : node4545;
															assign node4545 = (inp[0]) ? node4549 : node4546;
																assign node4546 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node4549 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node4553 = (inp[0]) ? node4555 : 4'b1001;
														assign node4555 = (inp[13]) ? node4557 : 4'b1000;
															assign node4557 = (inp[10]) ? node4559 : 4'b1001;
																assign node4559 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node4562 = (inp[7]) ? node4614 : node4563;
											assign node4563 = (inp[10]) ? node4587 : node4564;
												assign node4564 = (inp[13]) ? node4578 : node4565;
													assign node4565 = (inp[11]) ? node4571 : node4566;
														assign node4566 = (inp[0]) ? node4568 : 4'b1000;
															assign node4568 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node4571 = (inp[4]) ? node4575 : node4572;
															assign node4572 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node4575 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node4578 = (inp[0]) ? node4580 : 4'b1011;
														assign node4580 = (inp[12]) ? node4582 : 4'b1010;
															assign node4582 = (inp[4]) ? node4584 : 4'b1010;
																assign node4584 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4587 = (inp[13]) ? node4595 : node4588;
													assign node4588 = (inp[0]) ? node4592 : node4589;
														assign node4589 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node4592 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node4595 = (inp[12]) ? node4605 : node4596;
														assign node4596 = (inp[4]) ? node4602 : node4597;
															assign node4597 = (inp[11]) ? node4599 : 4'b1001;
																assign node4599 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node4602 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node4605 = (inp[4]) ? node4607 : 4'b1010;
															assign node4607 = (inp[0]) ? node4611 : node4608;
																assign node4608 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node4611 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node4614 = (inp[12]) ? node4644 : node4615;
												assign node4615 = (inp[4]) ? node4631 : node4616;
													assign node4616 = (inp[10]) ? node4622 : node4617;
														assign node4617 = (inp[0]) ? node4619 : 4'b1101;
															assign node4619 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node4622 = (inp[13]) ? node4626 : node4623;
															assign node4623 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node4626 = (inp[11]) ? node4628 : 4'b1100;
																assign node4628 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node4631 = (inp[0]) ? node4637 : node4632;
														assign node4632 = (inp[10]) ? node4634 : 4'b1110;
															assign node4634 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node4637 = (inp[13]) ? 4'b1111 : node4638;
															assign node4638 = (inp[11]) ? 4'b1111 : node4639;
																assign node4639 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node4644 = (inp[4]) ? node4654 : node4645;
													assign node4645 = (inp[11]) ? 4'b1111 : node4646;
														assign node4646 = (inp[0]) ? 4'b1111 : node4647;
															assign node4647 = (inp[10]) ? 4'b1110 : node4648;
																assign node4648 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node4654 = (inp[13]) ? node4660 : node4655;
														assign node4655 = (inp[11]) ? 4'b1000 : node4656;
															assign node4656 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node4660 = (inp[11]) ? node4662 : 4'b1001;
															assign node4662 = (inp[10]) ? 4'b1000 : 4'b1001;
									assign node4665 = (inp[7]) ? node4757 : node4666;
										assign node4666 = (inp[12]) ? node4722 : node4667;
											assign node4667 = (inp[4]) ? node4701 : node4668;
												assign node4668 = (inp[5]) ? node4686 : node4669;
													assign node4669 = (inp[11]) ? node4675 : node4670;
														assign node4670 = (inp[0]) ? 4'b1100 : node4671;
															assign node4671 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node4675 = (inp[0]) ? node4681 : node4676;
															assign node4676 = (inp[13]) ? node4678 : 4'b1100;
																assign node4678 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node4681 = (inp[13]) ? node4683 : 4'b1101;
																assign node4683 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node4686 = (inp[13]) ? 4'b1101 : node4687;
														assign node4687 = (inp[11]) ? node4693 : node4688;
															assign node4688 = (inp[10]) ? node4690 : 4'b1101;
																assign node4690 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node4693 = (inp[0]) ? node4697 : node4694;
																assign node4694 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node4697 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node4701 = (inp[5]) ? node4711 : node4702;
													assign node4702 = (inp[10]) ? 4'b1111 : node4703;
														assign node4703 = (inp[0]) ? 4'b1111 : node4704;
															assign node4704 = (inp[11]) ? node4706 : 4'b1110;
																assign node4706 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node4711 = (inp[10]) ? node4713 : 4'b1110;
														assign node4713 = (inp[0]) ? node4719 : node4714;
															assign node4714 = (inp[13]) ? 4'b1110 : node4715;
																assign node4715 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node4719 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node4722 = (inp[4]) ? node4738 : node4723;
												assign node4723 = (inp[5]) ? node4733 : node4724;
													assign node4724 = (inp[0]) ? node4726 : 4'b1110;
														assign node4726 = (inp[10]) ? node4728 : 4'b1111;
															assign node4728 = (inp[13]) ? node4730 : 4'b1111;
																assign node4730 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node4733 = (inp[13]) ? 4'b1111 : node4734;
														assign node4734 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node4738 = (inp[5]) ? node4750 : node4739;
													assign node4739 = (inp[11]) ? node4741 : 4'b1000;
														assign node4741 = (inp[13]) ? 4'b1001 : node4742;
															assign node4742 = (inp[0]) ? node4746 : node4743;
																assign node4743 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node4746 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node4750 = (inp[13]) ? 4'b1101 : node4751;
														assign node4751 = (inp[10]) ? node4753 : 4'b1100;
															assign node4753 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node4757 = (inp[5]) ? node4795 : node4758;
											assign node4758 = (inp[13]) ? node4778 : node4759;
												assign node4759 = (inp[11]) ? node4767 : node4760;
													assign node4760 = (inp[0]) ? node4762 : 4'b1111;
														assign node4762 = (inp[4]) ? 4'b1101 : node4763;
															assign node4763 = (inp[12]) ? 4'b1110 : 4'b1101;
													assign node4767 = (inp[12]) ? node4775 : node4768;
														assign node4768 = (inp[4]) ? 4'b1110 : node4769;
															assign node4769 = (inp[0]) ? 4'b1101 : node4770;
																assign node4770 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node4775 = (inp[4]) ? 4'b1101 : 4'b1111;
												assign node4778 = (inp[11]) ? node4786 : node4779;
													assign node4779 = (inp[0]) ? node4781 : 4'b1100;
														assign node4781 = (inp[12]) ? 4'b1100 : node4782;
															assign node4782 = (inp[4]) ? 4'b1110 : 4'b1100;
													assign node4786 = (inp[0]) ? node4790 : node4787;
														assign node4787 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node4790 = (inp[4]) ? node4792 : 4'b1111;
															assign node4792 = (inp[12]) ? 4'b1101 : 4'b1111;
											assign node4795 = (inp[12]) ? node4833 : node4796;
												assign node4796 = (inp[4]) ? node4810 : node4797;
													assign node4797 = (inp[10]) ? node4807 : node4798;
														assign node4798 = (inp[0]) ? node4804 : node4799;
															assign node4799 = (inp[13]) ? 4'b1000 : node4800;
																assign node4800 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node4804 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node4807 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node4810 = (inp[11]) ? node4826 : node4811;
														assign node4811 = (inp[13]) ? node4819 : node4812;
															assign node4812 = (inp[0]) ? node4816 : node4813;
																assign node4813 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node4816 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node4819 = (inp[0]) ? node4823 : node4820;
																assign node4820 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node4823 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node4826 = (inp[13]) ? node4828 : 4'b1011;
															assign node4828 = (inp[0]) ? node4830 : 4'b1011;
																assign node4830 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node4833 = (inp[4]) ? node4847 : node4834;
													assign node4834 = (inp[10]) ? node4840 : node4835;
														assign node4835 = (inp[0]) ? 4'b1010 : node4836;
															assign node4836 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node4840 = (inp[11]) ? node4842 : 4'b1011;
															assign node4842 = (inp[13]) ? node4844 : 4'b1010;
																assign node4844 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node4847 = (inp[11]) ? 4'b1100 : node4848;
														assign node4848 = (inp[0]) ? node4850 : 4'b1101;
															assign node4850 = (inp[10]) ? node4854 : node4851;
																assign node4851 = (inp[13]) ? 4'b1101 : 4'b1100;
																assign node4854 = (inp[13]) ? 4'b1100 : 4'b1101;
								assign node4858 = (inp[1]) ? node5046 : node4859;
									assign node4859 = (inp[5]) ? node4947 : node4860;
										assign node4860 = (inp[12]) ? node4904 : node4861;
											assign node4861 = (inp[4]) ? node4883 : node4862;
												assign node4862 = (inp[7]) ? node4872 : node4863;
													assign node4863 = (inp[13]) ? 4'b1101 : node4864;
														assign node4864 = (inp[0]) ? node4868 : node4865;
															assign node4865 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node4868 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node4872 = (inp[0]) ? 4'b1100 : node4873;
														assign node4873 = (inp[11]) ? node4877 : node4874;
															assign node4874 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node4877 = (inp[13]) ? node4879 : 4'b1101;
																assign node4879 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node4883 = (inp[13]) ? node4891 : node4884;
													assign node4884 = (inp[10]) ? node4888 : node4885;
														assign node4885 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node4888 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node4891 = (inp[0]) ? node4897 : node4892;
														assign node4892 = (inp[10]) ? node4894 : 4'b1111;
															assign node4894 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node4897 = (inp[10]) ? node4901 : node4898;
															assign node4898 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node4901 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node4904 = (inp[4]) ? node4922 : node4905;
												assign node4905 = (inp[10]) ? node4919 : node4906;
													assign node4906 = (inp[0]) ? node4912 : node4907;
														assign node4907 = (inp[7]) ? node4909 : 4'b1110;
															assign node4909 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node4912 = (inp[7]) ? node4914 : 4'b1111;
															assign node4914 = (inp[13]) ? 4'b1110 : node4915;
																assign node4915 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node4919 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node4922 = (inp[7]) ? node4936 : node4923;
													assign node4923 = (inp[0]) ? 4'b1000 : node4924;
														assign node4924 = (inp[10]) ? node4930 : node4925;
															assign node4925 = (inp[11]) ? 4'b1000 : node4926;
																assign node4926 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node4930 = (inp[11]) ? 4'b1001 : node4931;
																assign node4931 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node4936 = (inp[0]) ? node4940 : node4937;
														assign node4937 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node4940 = (inp[10]) ? node4942 : 4'b1101;
															assign node4942 = (inp[13]) ? node4944 : 4'b1100;
																assign node4944 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node4947 = (inp[7]) ? node4997 : node4948;
											assign node4948 = (inp[12]) ? node4980 : node4949;
												assign node4949 = (inp[4]) ? node4963 : node4950;
													assign node4950 = (inp[11]) ? 4'b1100 : node4951;
														assign node4951 = (inp[13]) ? node4957 : node4952;
															assign node4952 = (inp[0]) ? node4954 : 4'b1101;
																assign node4954 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node4957 = (inp[10]) ? node4959 : 4'b1100;
																assign node4959 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node4963 = (inp[11]) ? node4969 : node4964;
														assign node4964 = (inp[13]) ? 4'b1111 : node4965;
															assign node4965 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node4969 = (inp[13]) ? node4975 : node4970;
															assign node4970 = (inp[10]) ? node4972 : 4'b1111;
																assign node4972 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node4975 = (inp[0]) ? node4977 : 4'b1110;
																assign node4977 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node4980 = (inp[4]) ? node4984 : node4981;
													assign node4981 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node4984 = (inp[11]) ? node4992 : node4985;
														assign node4985 = (inp[10]) ? node4989 : node4986;
															assign node4986 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node4989 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node4992 = (inp[13]) ? 4'b1101 : node4993;
															assign node4993 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node4997 = (inp[4]) ? node5025 : node4998;
												assign node4998 = (inp[12]) ? node5014 : node4999;
													assign node4999 = (inp[0]) ? node5005 : node5000;
														assign node5000 = (inp[10]) ? node5002 : 4'b1000;
															assign node5002 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node5005 = (inp[10]) ? node5011 : node5006;
															assign node5006 = (inp[11]) ? 4'b1001 : node5007;
																assign node5007 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node5011 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5014 = (inp[0]) ? node5020 : node5015;
														assign node5015 = (inp[11]) ? 4'b1011 : node5016;
															assign node5016 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node5020 = (inp[10]) ? 4'b1010 : node5021;
															assign node5021 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node5025 = (inp[12]) ? node5031 : node5026;
													assign node5026 = (inp[0]) ? node5028 : 4'b1011;
														assign node5028 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node5031 = (inp[11]) ? node5041 : node5032;
														assign node5032 = (inp[10]) ? node5034 : 4'b1101;
															assign node5034 = (inp[13]) ? node5038 : node5035;
																assign node5035 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node5038 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5041 = (inp[13]) ? node5043 : 4'b1100;
															assign node5043 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node5046 = (inp[5]) ? node5146 : node5047;
										assign node5047 = (inp[4]) ? node5097 : node5048;
											assign node5048 = (inp[12]) ? node5068 : node5049;
												assign node5049 = (inp[10]) ? node5059 : node5050;
													assign node5050 = (inp[0]) ? node5056 : node5051;
														assign node5051 = (inp[13]) ? 4'b1001 : node5052;
															assign node5052 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node5056 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5059 = (inp[0]) ? node5065 : node5060;
														assign node5060 = (inp[11]) ? 4'b1000 : node5061;
															assign node5061 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node5065 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node5068 = (inp[7]) ? node5084 : node5069;
													assign node5069 = (inp[11]) ? 4'b1011 : node5070;
														assign node5070 = (inp[0]) ? node5076 : node5071;
															assign node5071 = (inp[13]) ? node5073 : 4'b1011;
																assign node5073 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node5076 = (inp[13]) ? node5080 : node5077;
																assign node5077 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node5080 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node5084 = (inp[13]) ? node5090 : node5085;
														assign node5085 = (inp[10]) ? 4'b1010 : node5086;
															assign node5086 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5090 = (inp[11]) ? 4'b1011 : node5091;
															assign node5091 = (inp[10]) ? node5093 : 4'b1010;
																assign node5093 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node5097 = (inp[12]) ? node5113 : node5098;
												assign node5098 = (inp[10]) ? node5106 : node5099;
													assign node5099 = (inp[0]) ? node5101 : 4'b1010;
														assign node5101 = (inp[7]) ? 4'b1011 : node5102;
															assign node5102 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node5106 = (inp[7]) ? 4'b1011 : node5107;
														assign node5107 = (inp[13]) ? node5109 : 4'b1010;
															assign node5109 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5113 = (inp[7]) ? node5125 : node5114;
													assign node5114 = (inp[13]) ? node5122 : node5115;
														assign node5115 = (inp[0]) ? 4'b1101 : node5116;
															assign node5116 = (inp[10]) ? node5118 : 4'b1100;
																assign node5118 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node5122 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5125 = (inp[13]) ? node5133 : node5126;
														assign node5126 = (inp[0]) ? node5128 : 4'b1000;
															assign node5128 = (inp[11]) ? 4'b1000 : node5129;
																assign node5129 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node5133 = (inp[11]) ? node5139 : node5134;
															assign node5134 = (inp[10]) ? node5136 : 4'b1000;
																assign node5136 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node5139 = (inp[10]) ? node5143 : node5140;
																assign node5140 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node5143 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node5146 = (inp[7]) ? node5182 : node5147;
											assign node5147 = (inp[0]) ? node5163 : node5148;
												assign node5148 = (inp[13]) ? node5150 : 4'b1001;
													assign node5150 = (inp[10]) ? node5156 : node5151;
														assign node5151 = (inp[11]) ? node5153 : 4'b1010;
															assign node5153 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node5156 = (inp[4]) ? node5160 : node5157;
															assign node5157 = (inp[12]) ? 4'b1011 : 4'b1000;
															assign node5160 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node5163 = (inp[12]) ? node5173 : node5164;
													assign node5164 = (inp[4]) ? node5168 : node5165;
														assign node5165 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node5168 = (inp[10]) ? node5170 : 4'b1010;
															assign node5170 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node5173 = (inp[4]) ? node5179 : node5174;
														assign node5174 = (inp[11]) ? node5176 : 4'b1010;
															assign node5176 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5179 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node5182 = (inp[4]) ? node5212 : node5183;
												assign node5183 = (inp[12]) ? node5189 : node5184;
													assign node5184 = (inp[13]) ? node5186 : 4'b1101;
														assign node5186 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5189 = (inp[13]) ? node5197 : node5190;
														assign node5190 = (inp[11]) ? 4'b1110 : node5191;
															assign node5191 = (inp[10]) ? node5193 : 4'b1110;
																assign node5193 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node5197 = (inp[10]) ? node5205 : node5198;
															assign node5198 = (inp[0]) ? node5202 : node5199;
																assign node5199 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node5202 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node5205 = (inp[11]) ? node5209 : node5206;
																assign node5206 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node5209 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node5212 = (inp[12]) ? node5226 : node5213;
													assign node5213 = (inp[13]) ? node5219 : node5214;
														assign node5214 = (inp[0]) ? 4'b1110 : node5215;
															assign node5215 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node5219 = (inp[11]) ? node5221 : 4'b1110;
															assign node5221 = (inp[10]) ? 4'b1111 : node5222;
																assign node5222 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5226 = (inp[0]) ? node5236 : node5227;
														assign node5227 = (inp[13]) ? node5229 : 4'b1000;
															assign node5229 = (inp[10]) ? node5233 : node5230;
																assign node5230 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node5233 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node5236 = (inp[10]) ? node5240 : node5237;
															assign node5237 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node5240 = (inp[13]) ? node5242 : 4'b1001;
																assign node5242 = (inp[11]) ? 4'b1000 : 4'b1001;
							assign node5245 = (inp[1]) ? node5637 : node5246;
								assign node5246 = (inp[2]) ? node5428 : node5247;
									assign node5247 = (inp[7]) ? node5331 : node5248;
										assign node5248 = (inp[5]) ? node5298 : node5249;
											assign node5249 = (inp[4]) ? node5273 : node5250;
												assign node5250 = (inp[12]) ? node5266 : node5251;
													assign node5251 = (inp[10]) ? node5261 : node5252;
														assign node5252 = (inp[11]) ? 4'b1001 : node5253;
															assign node5253 = (inp[13]) ? node5257 : node5254;
																assign node5254 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node5257 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5261 = (inp[11]) ? node5263 : 4'b1001;
															assign node5263 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node5266 = (inp[10]) ? node5268 : 4'b1011;
														assign node5268 = (inp[13]) ? 4'b1011 : node5269;
															assign node5269 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5273 = (inp[12]) ? node5289 : node5274;
													assign node5274 = (inp[13]) ? node5280 : node5275;
														assign node5275 = (inp[0]) ? node5277 : 4'b1010;
															assign node5277 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5280 = (inp[10]) ? 4'b1011 : node5281;
															assign node5281 = (inp[0]) ? node5285 : node5282;
																assign node5282 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node5285 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node5289 = (inp[13]) ? node5291 : 4'b1001;
														assign node5291 = (inp[10]) ? node5295 : node5292;
															assign node5292 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node5295 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node5298 = (inp[12]) ? node5316 : node5299;
												assign node5299 = (inp[4]) ? node5307 : node5300;
													assign node5300 = (inp[0]) ? node5302 : 4'b1001;
														assign node5302 = (inp[13]) ? node5304 : 4'b1000;
															assign node5304 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5307 = (inp[13]) ? node5309 : 4'b1110;
														assign node5309 = (inp[10]) ? node5313 : node5310;
															assign node5310 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5313 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node5316 = (inp[4]) ? node5324 : node5317;
													assign node5317 = (inp[11]) ? node5319 : 4'b1011;
														assign node5319 = (inp[0]) ? node5321 : 4'b1010;
															assign node5321 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node5324 = (inp[10]) ? 4'b1001 : node5325;
														assign node5325 = (inp[11]) ? node5327 : 4'b1000;
															assign node5327 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node5331 = (inp[5]) ? node5377 : node5332;
											assign node5332 = (inp[4]) ? node5356 : node5333;
												assign node5333 = (inp[12]) ? node5343 : node5334;
													assign node5334 = (inp[10]) ? node5338 : node5335;
														assign node5335 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node5338 = (inp[13]) ? node5340 : 4'b1100;
															assign node5340 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node5343 = (inp[11]) ? node5349 : node5344;
														assign node5344 = (inp[0]) ? 4'b1110 : node5345;
															assign node5345 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5349 = (inp[13]) ? 4'b1111 : node5350;
															assign node5350 = (inp[0]) ? 4'b1111 : node5351;
																assign node5351 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node5356 = (inp[12]) ? node5370 : node5357;
													assign node5357 = (inp[10]) ? node5365 : node5358;
														assign node5358 = (inp[0]) ? 4'b1011 : node5359;
															assign node5359 = (inp[11]) ? node5361 : 4'b1010;
																assign node5361 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node5365 = (inp[0]) ? 4'b1010 : node5366;
															assign node5366 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node5370 = (inp[0]) ? 4'b1100 : node5371;
														assign node5371 = (inp[11]) ? 4'b1101 : node5372;
															assign node5372 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node5377 = (inp[0]) ? node5401 : node5378;
												assign node5378 = (inp[13]) ? node5392 : node5379;
													assign node5379 = (inp[12]) ? node5387 : node5380;
														assign node5380 = (inp[4]) ? node5384 : node5381;
															assign node5381 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node5384 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node5387 = (inp[4]) ? 4'b1001 : node5388;
															assign node5388 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node5392 = (inp[12]) ? node5398 : node5393;
														assign node5393 = (inp[11]) ? 4'b1010 : node5394;
															assign node5394 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5398 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node5401 = (inp[13]) ? node5417 : node5402;
													assign node5402 = (inp[11]) ? node5408 : node5403;
														assign node5403 = (inp[12]) ? 4'b1010 : node5404;
															assign node5404 = (inp[4]) ? 4'b1010 : 4'b1001;
														assign node5408 = (inp[4]) ? node5412 : node5409;
															assign node5409 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node5412 = (inp[12]) ? node5414 : 4'b1011;
																assign node5414 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node5417 = (inp[12]) ? node5425 : node5418;
														assign node5418 = (inp[4]) ? node5420 : 4'b1001;
															assign node5420 = (inp[11]) ? node5422 : 4'b1011;
																assign node5422 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5425 = (inp[4]) ? 4'b1001 : 4'b1011;
									assign node5428 = (inp[7]) ? node5518 : node5429;
										assign node5429 = (inp[5]) ? node5479 : node5430;
											assign node5430 = (inp[4]) ? node5452 : node5431;
												assign node5431 = (inp[12]) ? node5441 : node5432;
													assign node5432 = (inp[11]) ? node5434 : 4'b1100;
														assign node5434 = (inp[13]) ? node5438 : node5435;
															assign node5435 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node5438 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node5441 = (inp[10]) ? node5447 : node5442;
														assign node5442 = (inp[0]) ? node5444 : 4'b1110;
															assign node5444 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node5447 = (inp[0]) ? node5449 : 4'b1111;
															assign node5449 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node5452 = (inp[12]) ? node5470 : node5453;
													assign node5453 = (inp[11]) ? node5463 : node5454;
														assign node5454 = (inp[0]) ? node5456 : 4'b1110;
															assign node5456 = (inp[10]) ? node5460 : node5457;
																assign node5457 = (inp[13]) ? 4'b1111 : 4'b1110;
																assign node5460 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node5463 = (inp[13]) ? node5465 : 4'b1111;
															assign node5465 = (inp[0]) ? 4'b1111 : node5466;
																assign node5466 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node5470 = (inp[11]) ? 4'b1100 : node5471;
														assign node5471 = (inp[13]) ? node5475 : node5472;
															assign node5472 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5475 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node5479 = (inp[4]) ? node5501 : node5480;
												assign node5480 = (inp[12]) ? node5488 : node5481;
													assign node5481 = (inp[0]) ? 4'b1100 : node5482;
														assign node5482 = (inp[10]) ? 4'b1101 : node5483;
															assign node5483 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node5488 = (inp[13]) ? node5494 : node5489;
														assign node5489 = (inp[10]) ? node5491 : 4'b1110;
															assign node5491 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5494 = (inp[10]) ? node5496 : 4'b1111;
															assign node5496 = (inp[0]) ? 4'b1110 : node5497;
																assign node5497 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node5501 = (inp[12]) ? 4'b1100 : node5502;
													assign node5502 = (inp[0]) ? node5514 : node5503;
														assign node5503 = (inp[10]) ? node5509 : node5504;
															assign node5504 = (inp[13]) ? node5506 : 4'b1010;
																assign node5506 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node5509 = (inp[11]) ? 4'b1011 : node5510;
																assign node5510 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node5514 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node5518 = (inp[5]) ? node5570 : node5519;
											assign node5519 = (inp[12]) ? node5543 : node5520;
												assign node5520 = (inp[4]) ? node5536 : node5521;
													assign node5521 = (inp[13]) ? 4'b1000 : node5522;
														assign node5522 = (inp[0]) ? node5528 : node5523;
															assign node5523 = (inp[11]) ? node5525 : 4'b1000;
																assign node5525 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node5528 = (inp[10]) ? node5532 : node5529;
																assign node5529 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node5532 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5536 = (inp[11]) ? 4'b1111 : node5537;
														assign node5537 = (inp[10]) ? node5539 : 4'b1110;
															assign node5539 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node5543 = (inp[4]) ? node5555 : node5544;
													assign node5544 = (inp[0]) ? node5546 : 4'b1011;
														assign node5546 = (inp[10]) ? node5550 : node5547;
															assign node5547 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node5550 = (inp[13]) ? node5552 : 4'b1011;
																assign node5552 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node5555 = (inp[11]) ? node5565 : node5556;
														assign node5556 = (inp[13]) ? node5560 : node5557;
															assign node5557 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node5560 = (inp[10]) ? node5562 : 4'b1001;
																assign node5562 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5565 = (inp[13]) ? node5567 : 4'b1000;
															assign node5567 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node5570 = (inp[11]) ? node5606 : node5571;
												assign node5571 = (inp[13]) ? node5591 : node5572;
													assign node5572 = (inp[12]) ? node5584 : node5573;
														assign node5573 = (inp[4]) ? node5581 : node5574;
															assign node5574 = (inp[10]) ? node5578 : node5575;
																assign node5575 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node5578 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5581 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5584 = (inp[4]) ? node5586 : 4'b1110;
															assign node5586 = (inp[10]) ? 4'b1100 : node5587;
																assign node5587 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node5591 = (inp[0]) ? node5603 : node5592;
														assign node5592 = (inp[10]) ? node5600 : node5593;
															assign node5593 = (inp[12]) ? node5597 : node5594;
																assign node5594 = (inp[4]) ? 4'b1110 : 4'b1101;
																assign node5597 = (inp[4]) ? 4'b1101 : 4'b1111;
															assign node5600 = (inp[4]) ? 4'b1100 : 4'b1110;
														assign node5603 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node5606 = (inp[13]) ? node5614 : node5607;
													assign node5607 = (inp[10]) ? node5611 : node5608;
														assign node5608 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node5611 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node5614 = (inp[4]) ? node5624 : node5615;
														assign node5615 = (inp[12]) ? node5619 : node5616;
															assign node5616 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node5619 = (inp[10]) ? node5621 : 4'b1111;
																assign node5621 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5624 = (inp[12]) ? node5630 : node5625;
															assign node5625 = (inp[10]) ? node5627 : 4'b1110;
																assign node5627 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5630 = (inp[10]) ? node5634 : node5631;
																assign node5631 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node5634 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node5637 = (inp[2]) ? node5809 : node5638;
									assign node5638 = (inp[5]) ? node5742 : node5639;
										assign node5639 = (inp[7]) ? node5691 : node5640;
											assign node5640 = (inp[13]) ? node5674 : node5641;
												assign node5641 = (inp[4]) ? node5661 : node5642;
													assign node5642 = (inp[12]) ? node5650 : node5643;
														assign node5643 = (inp[10]) ? node5645 : 4'b1100;
															assign node5645 = (inp[11]) ? 4'b1100 : node5646;
																assign node5646 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5650 = (inp[0]) ? node5656 : node5651;
															assign node5651 = (inp[11]) ? node5653 : 4'b1110;
																assign node5653 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node5656 = (inp[11]) ? node5658 : 4'b1111;
																assign node5658 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node5661 = (inp[12]) ? node5671 : node5662;
														assign node5662 = (inp[0]) ? node5664 : 4'b1111;
															assign node5664 = (inp[11]) ? node5668 : node5665;
																assign node5665 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node5668 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5671 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node5674 = (inp[10]) ? node5680 : node5675;
													assign node5675 = (inp[0]) ? 4'b1101 : node5676;
														assign node5676 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node5680 = (inp[12]) ? node5686 : node5681;
														assign node5681 = (inp[0]) ? node5683 : 4'b1111;
															assign node5683 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node5686 = (inp[4]) ? 4'b1101 : node5687;
															assign node5687 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5691 = (inp[4]) ? node5723 : node5692;
												assign node5692 = (inp[12]) ? node5706 : node5693;
													assign node5693 = (inp[13]) ? node5701 : node5694;
														assign node5694 = (inp[0]) ? node5698 : node5695;
															assign node5695 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node5698 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node5701 = (inp[10]) ? node5703 : 4'b1001;
															assign node5703 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node5706 = (inp[11]) ? node5714 : node5707;
														assign node5707 = (inp[13]) ? node5709 : 4'b1010;
															assign node5709 = (inp[10]) ? 4'b1010 : node5710;
																assign node5710 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5714 = (inp[0]) ? 4'b1011 : node5715;
															assign node5715 = (inp[10]) ? node5719 : node5716;
																assign node5716 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node5719 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node5723 = (inp[12]) ? node5731 : node5724;
													assign node5724 = (inp[13]) ? node5726 : 4'b1111;
														assign node5726 = (inp[0]) ? node5728 : 4'b1110;
															assign node5728 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5731 = (inp[0]) ? node5737 : node5732;
														assign node5732 = (inp[13]) ? node5734 : 4'b1000;
															assign node5734 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node5737 = (inp[10]) ? 4'b1001 : node5738;
															assign node5738 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node5742 = (inp[4]) ? node5788 : node5743;
											assign node5743 = (inp[12]) ? node5765 : node5744;
												assign node5744 = (inp[13]) ? node5756 : node5745;
													assign node5745 = (inp[10]) ? node5751 : node5746;
														assign node5746 = (inp[0]) ? 4'b1101 : node5747;
															assign node5747 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node5751 = (inp[7]) ? node5753 : 4'b1100;
															assign node5753 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5756 = (inp[0]) ? node5762 : node5757;
														assign node5757 = (inp[11]) ? 4'b1100 : node5758;
															assign node5758 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node5762 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node5765 = (inp[7]) ? node5775 : node5766;
													assign node5766 = (inp[13]) ? 4'b1111 : node5767;
														assign node5767 = (inp[11]) ? node5769 : 4'b1110;
															assign node5769 = (inp[10]) ? node5771 : 4'b1111;
																assign node5771 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node5775 = (inp[0]) ? node5783 : node5776;
														assign node5776 = (inp[10]) ? node5780 : node5777;
															assign node5777 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node5780 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node5783 = (inp[10]) ? node5785 : 4'b1110;
															assign node5785 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node5788 = (inp[12]) ? node5796 : node5789;
												assign node5789 = (inp[13]) ? node5791 : 4'b1111;
													assign node5791 = (inp[7]) ? 4'b1110 : node5792;
														assign node5792 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node5796 = (inp[10]) ? node5802 : node5797;
													assign node5797 = (inp[0]) ? 4'b1101 : node5798;
														assign node5798 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node5802 = (inp[0]) ? node5804 : 4'b1101;
														assign node5804 = (inp[11]) ? node5806 : 4'b1100;
															assign node5806 = (inp[13]) ? 4'b1100 : 4'b1101;
									assign node5809 = (inp[7]) ? node5889 : node5810;
										assign node5810 = (inp[4]) ? node5850 : node5811;
											assign node5811 = (inp[12]) ? node5835 : node5812;
												assign node5812 = (inp[10]) ? node5824 : node5813;
													assign node5813 = (inp[0]) ? node5819 : node5814;
														assign node5814 = (inp[11]) ? 4'b1001 : node5815;
															assign node5815 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node5819 = (inp[13]) ? node5821 : 4'b1000;
															assign node5821 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5824 = (inp[13]) ? node5828 : node5825;
														assign node5825 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node5828 = (inp[5]) ? 4'b1000 : node5829;
															assign node5829 = (inp[11]) ? 4'b1000 : node5830;
																assign node5830 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node5835 = (inp[10]) ? node5845 : node5836;
													assign node5836 = (inp[11]) ? 4'b1010 : node5837;
														assign node5837 = (inp[5]) ? node5839 : 4'b1011;
															assign node5839 = (inp[0]) ? node5841 : 4'b1010;
																assign node5841 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node5845 = (inp[0]) ? node5847 : 4'b1011;
														assign node5847 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node5850 = (inp[12]) ? node5876 : node5851;
												assign node5851 = (inp[5]) ? node5863 : node5852;
													assign node5852 = (inp[10]) ? node5860 : node5853;
														assign node5853 = (inp[0]) ? node5857 : node5854;
															assign node5854 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node5857 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node5860 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5863 = (inp[13]) ? node5871 : node5864;
														assign node5864 = (inp[10]) ? 4'b1110 : node5865;
															assign node5865 = (inp[0]) ? node5867 : 4'b1111;
																assign node5867 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node5871 = (inp[0]) ? 4'b1111 : node5872;
															assign node5872 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node5876 = (inp[11]) ? node5882 : node5877;
													assign node5877 = (inp[0]) ? 4'b1001 : node5878;
														assign node5878 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node5882 = (inp[13]) ? 4'b1000 : node5883;
														assign node5883 = (inp[10]) ? node5885 : 4'b1000;
															assign node5885 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node5889 = (inp[5]) ? node5935 : node5890;
											assign node5890 = (inp[12]) ? node5916 : node5891;
												assign node5891 = (inp[4]) ? node5903 : node5892;
													assign node5892 = (inp[10]) ? 4'b1101 : node5893;
														assign node5893 = (inp[13]) ? node5895 : 4'b1101;
															assign node5895 = (inp[11]) ? node5899 : node5896;
																assign node5896 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node5899 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5903 = (inp[13]) ? node5911 : node5904;
														assign node5904 = (inp[10]) ? node5906 : 4'b1011;
															assign node5906 = (inp[0]) ? node5908 : 4'b1010;
																assign node5908 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node5911 = (inp[10]) ? 4'b1011 : node5912;
															assign node5912 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node5916 = (inp[4]) ? node5928 : node5917;
													assign node5917 = (inp[10]) ? node5923 : node5918;
														assign node5918 = (inp[0]) ? node5920 : 4'b1110;
															assign node5920 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node5923 = (inp[0]) ? node5925 : 4'b1111;
															assign node5925 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node5928 = (inp[10]) ? node5930 : 4'b1100;
														assign node5930 = (inp[0]) ? node5932 : 4'b1101;
															assign node5932 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node5935 = (inp[10]) ? node5947 : node5936;
												assign node5936 = (inp[0]) ? node5944 : node5937;
													assign node5937 = (inp[12]) ? node5941 : node5938;
														assign node5938 = (inp[13]) ? 4'b1000 : 4'b1010;
														assign node5941 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node5944 = (inp[13]) ? 4'b1011 : 4'b1001;
												assign node5947 = (inp[0]) ? node5965 : node5948;
													assign node5948 = (inp[11]) ? node5956 : node5949;
														assign node5949 = (inp[13]) ? node5951 : 4'b1011;
															assign node5951 = (inp[12]) ? node5953 : 4'b1001;
																assign node5953 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node5956 = (inp[13]) ? node5960 : node5957;
															assign node5957 = (inp[12]) ? 4'b1001 : 4'b1000;
															assign node5960 = (inp[12]) ? node5962 : 4'b1001;
																assign node5962 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node5965 = (inp[4]) ? node5973 : node5966;
														assign node5966 = (inp[12]) ? 4'b1010 : node5967;
															assign node5967 = (inp[13]) ? 4'b1000 : node5968;
																assign node5968 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node5973 = (inp[12]) ? node5977 : node5974;
															assign node5974 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node5977 = (inp[11]) ? 4'b1000 : 4'b1001;
				assign node5980 = (inp[5]) ? node8896 : node5981;
					assign node5981 = (inp[0]) ? node7379 : node5982;
						assign node5982 = (inp[10]) ? node6708 : node5983;
							assign node5983 = (inp[8]) ? node6371 : node5984;
								assign node5984 = (inp[12]) ? node6174 : node5985;
									assign node5985 = (inp[7]) ? node6073 : node5986;
										assign node5986 = (inp[4]) ? node6026 : node5987;
											assign node5987 = (inp[15]) ? node6005 : node5988;
												assign node5988 = (inp[9]) ? node5998 : node5989;
													assign node5989 = (inp[13]) ? node5991 : 4'b1100;
														assign node5991 = (inp[2]) ? node5995 : node5992;
															assign node5992 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node5995 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5998 = (inp[2]) ? node6002 : node5999;
														assign node5999 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node6002 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node6005 = (inp[9]) ? node6017 : node6006;
													assign node6006 = (inp[2]) ? node6010 : node6007;
														assign node6007 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node6010 = (inp[13]) ? 4'b1010 : node6011;
															assign node6011 = (inp[11]) ? 4'b1110 : node6012;
																assign node6012 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node6017 = (inp[11]) ? node6019 : 4'b1011;
														assign node6019 = (inp[1]) ? node6021 : 4'b1010;
															assign node6021 = (inp[2]) ? 4'b1011 : node6022;
																assign node6022 = (inp[13]) ? 4'b1110 : 4'b1011;
											assign node6026 = (inp[13]) ? node6054 : node6027;
												assign node6027 = (inp[11]) ? node6039 : node6028;
													assign node6028 = (inp[9]) ? node6034 : node6029;
														assign node6029 = (inp[2]) ? 4'b1101 : node6030;
															assign node6030 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node6034 = (inp[15]) ? node6036 : 4'b1100;
															assign node6036 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node6039 = (inp[2]) ? node6047 : node6040;
														assign node6040 = (inp[15]) ? node6044 : node6041;
															assign node6041 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node6044 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node6047 = (inp[15]) ? node6049 : 4'b1100;
															assign node6049 = (inp[9]) ? node6051 : 4'b1000;
																assign node6051 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node6054 = (inp[2]) ? node6062 : node6055;
													assign node6055 = (inp[15]) ? node6057 : 4'b1101;
														assign node6057 = (inp[11]) ? node6059 : 4'b1001;
															assign node6059 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node6062 = (inp[15]) ? node6068 : node6063;
														assign node6063 = (inp[11]) ? 4'b1001 : node6064;
															assign node6064 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6068 = (inp[1]) ? 4'b1100 : node6069;
															assign node6069 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node6073 = (inp[15]) ? node6125 : node6074;
											assign node6074 = (inp[4]) ? node6098 : node6075;
												assign node6075 = (inp[9]) ? node6087 : node6076;
													assign node6076 = (inp[13]) ? node6080 : node6077;
														assign node6077 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node6080 = (inp[2]) ? node6084 : node6081;
															assign node6081 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node6084 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node6087 = (inp[2]) ? node6093 : node6088;
														assign node6088 = (inp[13]) ? 4'b1111 : node6089;
															assign node6089 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node6093 = (inp[13]) ? node6095 : 4'b1111;
															assign node6095 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node6098 = (inp[11]) ? node6112 : node6099;
													assign node6099 = (inp[9]) ? node6107 : node6100;
														assign node6100 = (inp[1]) ? node6104 : node6101;
															assign node6101 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node6104 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node6107 = (inp[2]) ? 4'b1011 : node6108;
															assign node6108 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node6112 = (inp[9]) ? node6116 : node6113;
														assign node6113 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node6116 = (inp[1]) ? 4'b1110 : node6117;
															assign node6117 = (inp[2]) ? node6121 : node6118;
																assign node6118 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node6121 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node6125 = (inp[4]) ? node6153 : node6126;
												assign node6126 = (inp[11]) ? node6142 : node6127;
													assign node6127 = (inp[13]) ? 4'b1100 : node6128;
														assign node6128 = (inp[9]) ? node6136 : node6129;
															assign node6129 = (inp[2]) ? node6133 : node6130;
																assign node6130 = (inp[1]) ? 4'b1001 : 4'b1100;
																assign node6133 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node6136 = (inp[1]) ? node6138 : 4'b1101;
																assign node6138 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node6142 = (inp[1]) ? node6150 : node6143;
														assign node6143 = (inp[9]) ? node6147 : node6144;
															assign node6144 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node6147 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node6150 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node6153 = (inp[9]) ? node6159 : node6154;
													assign node6154 = (inp[2]) ? node6156 : 4'b1111;
														assign node6156 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node6159 = (inp[11]) ? 4'b1011 : node6160;
														assign node6160 = (inp[1]) ? node6166 : node6161;
															assign node6161 = (inp[13]) ? 4'b1010 : node6162;
																assign node6162 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node6166 = (inp[13]) ? node6170 : node6167;
																assign node6167 = (inp[2]) ? 4'b1111 : 4'b1010;
																assign node6170 = (inp[2]) ? 4'b1011 : 4'b1111;
									assign node6174 = (inp[7]) ? node6274 : node6175;
										assign node6175 = (inp[4]) ? node6227 : node6176;
											assign node6176 = (inp[15]) ? node6208 : node6177;
												assign node6177 = (inp[2]) ? node6197 : node6178;
													assign node6178 = (inp[13]) ? node6190 : node6179;
														assign node6179 = (inp[1]) ? node6187 : node6180;
															assign node6180 = (inp[9]) ? node6184 : node6181;
																assign node6181 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node6184 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node6187 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6190 = (inp[1]) ? 4'b1011 : node6191;
															assign node6191 = (inp[9]) ? 4'b1111 : node6192;
																assign node6192 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node6197 = (inp[9]) ? node6205 : node6198;
														assign node6198 = (inp[11]) ? node6202 : node6199;
															assign node6199 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node6202 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node6205 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node6208 = (inp[13]) ? node6216 : node6209;
													assign node6209 = (inp[2]) ? node6211 : 4'b1101;
														assign node6211 = (inp[9]) ? node6213 : 4'b1000;
															assign node6213 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node6216 = (inp[2]) ? node6222 : node6217;
														assign node6217 = (inp[11]) ? node6219 : 4'b1000;
															assign node6219 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6222 = (inp[9]) ? 4'b1100 : node6223;
															assign node6223 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node6227 = (inp[9]) ? node6249 : node6228;
												assign node6228 = (inp[13]) ? node6240 : node6229;
													assign node6229 = (inp[15]) ? node6235 : node6230;
														assign node6230 = (inp[11]) ? 4'b1110 : node6231;
															assign node6231 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node6235 = (inp[1]) ? node6237 : 4'b1010;
															assign node6237 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node6240 = (inp[2]) ? node6242 : 4'b1111;
														assign node6242 = (inp[15]) ? node6246 : node6243;
															assign node6243 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node6246 = (inp[1]) ? 4'b1110 : 4'b1011;
												assign node6249 = (inp[1]) ? node6259 : node6250;
													assign node6250 = (inp[13]) ? 4'b1110 : node6251;
														assign node6251 = (inp[11]) ? node6253 : 4'b1111;
															assign node6253 = (inp[2]) ? 4'b1110 : node6254;
																assign node6254 = (inp[15]) ? 4'b1011 : 4'b1110;
													assign node6259 = (inp[2]) ? node6267 : node6260;
														assign node6260 = (inp[13]) ? node6264 : node6261;
															assign node6261 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node6264 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node6267 = (inp[11]) ? 4'b1111 : node6268;
															assign node6268 = (inp[15]) ? 4'b1110 : node6269;
																assign node6269 = (inp[13]) ? 4'b1010 : 4'b1110;
										assign node6274 = (inp[4]) ? node6318 : node6275;
											assign node6275 = (inp[15]) ? node6297 : node6276;
												assign node6276 = (inp[1]) ? node6290 : node6277;
													assign node6277 = (inp[13]) ? node6285 : node6278;
														assign node6278 = (inp[2]) ? node6282 : node6279;
															assign node6279 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node6282 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6285 = (inp[2]) ? node6287 : 4'b1001;
															assign node6287 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node6290 = (inp[11]) ? 4'b1101 : node6291;
														assign node6291 = (inp[9]) ? 4'b1100 : node6292;
															assign node6292 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node6297 = (inp[11]) ? node6315 : node6298;
													assign node6298 = (inp[9]) ? node6310 : node6299;
														assign node6299 = (inp[1]) ? node6303 : node6300;
															assign node6300 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node6303 = (inp[13]) ? node6307 : node6304;
																assign node6304 = (inp[2]) ? 4'b1111 : 4'b1010;
																assign node6307 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node6310 = (inp[2]) ? node6312 : 4'b1110;
															assign node6312 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node6315 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node6318 = (inp[1]) ? node6338 : node6319;
												assign node6319 = (inp[11]) ? node6333 : node6320;
													assign node6320 = (inp[9]) ? node6328 : node6321;
														assign node6321 = (inp[2]) ? node6325 : node6322;
															assign node6322 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node6325 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node6328 = (inp[13]) ? 4'b1000 : node6329;
															assign node6329 = (inp[2]) ? 4'b1101 : 4'b1000;
													assign node6333 = (inp[9]) ? node6335 : 4'b1001;
														assign node6335 = (inp[15]) ? 4'b1101 : 4'b1001;
												assign node6338 = (inp[9]) ? node6350 : node6339;
													assign node6339 = (inp[11]) ? node6347 : node6340;
														assign node6340 = (inp[13]) ? node6344 : node6341;
															assign node6341 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node6344 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node6347 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node6350 = (inp[11]) ? node6360 : node6351;
														assign node6351 = (inp[15]) ? 4'b1101 : node6352;
															assign node6352 = (inp[13]) ? node6356 : node6353;
																assign node6353 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node6356 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node6360 = (inp[13]) ? node6368 : node6361;
															assign node6361 = (inp[2]) ? node6365 : node6362;
																assign node6362 = (inp[15]) ? 4'b1001 : 4'b1000;
																assign node6365 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node6368 = (inp[2]) ? 4'b1000 : 4'b1100;
								assign node6371 = (inp[11]) ? node6511 : node6372;
									assign node6372 = (inp[2]) ? node6432 : node6373;
										assign node6373 = (inp[1]) ? node6399 : node6374;
											assign node6374 = (inp[12]) ? node6386 : node6375;
												assign node6375 = (inp[4]) ? node6381 : node6376;
													assign node6376 = (inp[9]) ? node6378 : 4'b1000;
														assign node6378 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node6381 = (inp[15]) ? node6383 : 4'b1010;
														assign node6383 = (inp[7]) ? 4'b1010 : 4'b1111;
												assign node6386 = (inp[4]) ? node6392 : node6387;
													assign node6387 = (inp[15]) ? node6389 : 4'b1010;
														assign node6389 = (inp[7]) ? 4'b1010 : 4'b1111;
													assign node6392 = (inp[7]) ? 4'b1001 : node6393;
														assign node6393 = (inp[15]) ? 4'b1100 : node6394;
															assign node6394 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node6399 = (inp[12]) ? node6413 : node6400;
												assign node6400 = (inp[4]) ? node6406 : node6401;
													assign node6401 = (inp[13]) ? 4'b1100 : node6402;
														assign node6402 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node6406 = (inp[7]) ? node6408 : 4'b1010;
														assign node6408 = (inp[13]) ? 4'b1110 : node6409;
															assign node6409 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node6413 = (inp[4]) ? node6423 : node6414;
													assign node6414 = (inp[7]) ? node6420 : node6415;
														assign node6415 = (inp[15]) ? node6417 : 4'b1111;
															assign node6417 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node6420 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node6423 = (inp[7]) ? node6427 : node6424;
														assign node6424 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node6427 = (inp[13]) ? 4'b1100 : node6428;
															assign node6428 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node6432 = (inp[1]) ? node6480 : node6433;
											assign node6433 = (inp[7]) ? node6457 : node6434;
												assign node6434 = (inp[15]) ? node6448 : node6435;
													assign node6435 = (inp[13]) ? node6441 : node6436;
														assign node6436 = (inp[4]) ? node6438 : 4'b1100;
															assign node6438 = (inp[12]) ? 4'b1100 : 4'b1111;
														assign node6441 = (inp[4]) ? node6445 : node6442;
															assign node6442 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node6445 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node6448 = (inp[12]) ? node6452 : node6449;
														assign node6449 = (inp[4]) ? 4'b1011 : 4'b1100;
														assign node6452 = (inp[4]) ? 4'b1000 : node6453;
															assign node6453 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node6457 = (inp[4]) ? node6467 : node6458;
													assign node6458 = (inp[12]) ? node6464 : node6459;
														assign node6459 = (inp[13]) ? node6461 : 4'b1101;
															assign node6461 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node6464 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node6467 = (inp[12]) ? node6473 : node6468;
														assign node6468 = (inp[13]) ? 4'b1110 : node6469;
															assign node6469 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node6473 = (inp[9]) ? node6475 : 4'b1101;
															assign node6475 = (inp[13]) ? node6477 : 4'b1100;
																assign node6477 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node6480 = (inp[4]) ? node6494 : node6481;
												assign node6481 = (inp[12]) ? node6487 : node6482;
													assign node6482 = (inp[7]) ? node6484 : 4'b1001;
														assign node6484 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node6487 = (inp[7]) ? node6491 : node6488;
														assign node6488 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node6491 = (inp[15]) ? 4'b1011 : 4'b1111;
												assign node6494 = (inp[12]) ? node6500 : node6495;
													assign node6495 = (inp[15]) ? node6497 : 4'b1010;
														assign node6497 = (inp[7]) ? 4'b1011 : 4'b1110;
													assign node6500 = (inp[15]) ? node6506 : node6501;
														assign node6501 = (inp[13]) ? 4'b1000 : node6502;
															assign node6502 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node6506 = (inp[7]) ? 4'b1000 : node6507;
															assign node6507 = (inp[13]) ? 4'b1101 : 4'b1100;
									assign node6511 = (inp[7]) ? node6631 : node6512;
										assign node6512 = (inp[15]) ? node6564 : node6513;
											assign node6513 = (inp[13]) ? node6541 : node6514;
												assign node6514 = (inp[4]) ? node6528 : node6515;
													assign node6515 = (inp[12]) ? node6521 : node6516;
														assign node6516 = (inp[2]) ? 4'b1100 : node6517;
															assign node6517 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node6521 = (inp[1]) ? node6525 : node6522;
															assign node6522 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node6525 = (inp[2]) ? 4'b1011 : 4'b1110;
													assign node6528 = (inp[12]) ? node6536 : node6529;
														assign node6529 = (inp[2]) ? node6533 : node6530;
															assign node6530 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node6533 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6536 = (inp[1]) ? node6538 : 4'b1000;
															assign node6538 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node6541 = (inp[12]) ? node6555 : node6542;
													assign node6542 = (inp[4]) ? node6548 : node6543;
														assign node6543 = (inp[1]) ? 4'b1100 : node6544;
															assign node6544 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node6548 = (inp[2]) ? node6552 : node6549;
															assign node6549 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node6552 = (inp[1]) ? 4'b1010 : 4'b1111;
													assign node6555 = (inp[4]) ? 4'b1001 : node6556;
														assign node6556 = (inp[1]) ? node6560 : node6557;
															assign node6557 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node6560 = (inp[2]) ? 4'b1010 : 4'b1111;
											assign node6564 = (inp[13]) ? node6594 : node6565;
												assign node6565 = (inp[2]) ? node6579 : node6566;
													assign node6566 = (inp[4]) ? node6572 : node6567;
														assign node6567 = (inp[12]) ? node6569 : 4'b1001;
															assign node6569 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6572 = (inp[12]) ? node6576 : node6573;
															assign node6573 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node6576 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node6579 = (inp[1]) ? node6587 : node6580;
														assign node6580 = (inp[12]) ? node6584 : node6581;
															assign node6581 = (inp[4]) ? 4'b1011 : 4'b1100;
															assign node6584 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node6587 = (inp[9]) ? 4'b1101 : node6588;
															assign node6588 = (inp[4]) ? 4'b1110 : node6589;
																assign node6589 = (inp[12]) ? 4'b1110 : 4'b1001;
												assign node6594 = (inp[9]) ? node6610 : node6595;
													assign node6595 = (inp[4]) ? node6599 : node6596;
														assign node6596 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node6599 = (inp[12]) ? node6605 : node6600;
															assign node6600 = (inp[2]) ? node6602 : 4'b1111;
																assign node6602 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node6605 = (inp[2]) ? 4'b1101 : node6606;
																assign node6606 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node6610 = (inp[4]) ? node6618 : node6611;
														assign node6611 = (inp[12]) ? node6615 : node6612;
															assign node6612 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6615 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node6618 = (inp[12]) ? node6624 : node6619;
															assign node6619 = (inp[1]) ? 4'b1111 : node6620;
																assign node6620 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node6624 = (inp[2]) ? node6628 : node6625;
																assign node6625 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node6628 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node6631 = (inp[15]) ? node6673 : node6632;
											assign node6632 = (inp[13]) ? node6652 : node6633;
												assign node6633 = (inp[1]) ? node6639 : node6634;
													assign node6634 = (inp[2]) ? 4'b1100 : node6635;
														assign node6635 = (inp[12]) ? 4'b1000 : 4'b1011;
													assign node6639 = (inp[2]) ? node6645 : node6640;
														assign node6640 = (inp[12]) ? 4'b1011 : node6641;
															assign node6641 = (inp[4]) ? 4'b1111 : 4'b1101;
														assign node6645 = (inp[4]) ? node6649 : node6646;
															assign node6646 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node6649 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node6652 = (inp[9]) ? node6658 : node6653;
													assign node6653 = (inp[4]) ? 4'b1100 : node6654;
														assign node6654 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node6658 = (inp[4]) ? node6662 : node6659;
														assign node6659 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node6662 = (inp[12]) ? node6668 : node6663;
															assign node6663 = (inp[1]) ? node6665 : 4'b1010;
																assign node6665 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node6668 = (inp[2]) ? node6670 : 4'b1001;
																assign node6670 = (inp[1]) ? 4'b1000 : 4'b1100;
											assign node6673 = (inp[2]) ? node6687 : node6674;
												assign node6674 = (inp[1]) ? node6680 : node6675;
													assign node6675 = (inp[12]) ? 4'b1000 : node6676;
														assign node6676 = (inp[9]) ? 4'b1001 : 4'b1011;
													assign node6680 = (inp[12]) ? node6684 : node6681;
														assign node6681 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node6684 = (inp[4]) ? 4'b1100 : 4'b1111;
												assign node6687 = (inp[1]) ? node6699 : node6688;
													assign node6688 = (inp[13]) ? node6694 : node6689;
														assign node6689 = (inp[4]) ? node6691 : 4'b1100;
															assign node6691 = (inp[12]) ? 4'b1100 : 4'b1111;
														assign node6694 = (inp[4]) ? 4'b1111 : node6695;
															assign node6695 = (inp[12]) ? 4'b1110 : 4'b1100;
													assign node6699 = (inp[4]) ? node6705 : node6700;
														assign node6700 = (inp[12]) ? node6702 : 4'b1001;
															assign node6702 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node6705 = (inp[12]) ? 4'b1000 : 4'b1010;
							assign node6708 = (inp[7]) ? node7078 : node6709;
								assign node6709 = (inp[12]) ? node6879 : node6710;
									assign node6710 = (inp[15]) ? node6792 : node6711;
										assign node6711 = (inp[4]) ? node6749 : node6712;
											assign node6712 = (inp[1]) ? node6734 : node6713;
												assign node6713 = (inp[2]) ? node6723 : node6714;
													assign node6714 = (inp[8]) ? 4'b1001 : node6715;
														assign node6715 = (inp[13]) ? node6717 : 4'b1001;
															assign node6717 = (inp[11]) ? 4'b1101 : node6718;
																assign node6718 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node6723 = (inp[11]) ? node6729 : node6724;
														assign node6724 = (inp[9]) ? 4'b1100 : node6725;
															assign node6725 = (inp[8]) ? 4'b1100 : 4'b1000;
														assign node6729 = (inp[8]) ? 4'b1101 : node6730;
															assign node6730 = (inp[13]) ? 4'b1001 : 4'b1100;
												assign node6734 = (inp[2]) ? 4'b1000 : node6735;
													assign node6735 = (inp[8]) ? node6743 : node6736;
														assign node6736 = (inp[13]) ? 4'b1100 : node6737;
															assign node6737 = (inp[11]) ? 4'b1000 : node6738;
																assign node6738 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6743 = (inp[11]) ? node6745 : 4'b1101;
															assign node6745 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node6749 = (inp[8]) ? node6773 : node6750;
												assign node6750 = (inp[9]) ? node6764 : node6751;
													assign node6751 = (inp[11]) ? node6757 : node6752;
														assign node6752 = (inp[13]) ? 4'b1001 : node6753;
															assign node6753 = (inp[2]) ? 4'b1100 : 4'b1001;
														assign node6757 = (inp[2]) ? node6761 : node6758;
															assign node6758 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node6761 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node6764 = (inp[11]) ? node6766 : 4'b1101;
														assign node6766 = (inp[13]) ? node6770 : node6767;
															assign node6767 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node6770 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node6773 = (inp[13]) ? node6787 : node6774;
													assign node6774 = (inp[11]) ? node6782 : node6775;
														assign node6775 = (inp[2]) ? node6779 : node6776;
															assign node6776 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node6779 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node6782 = (inp[2]) ? 4'b1110 : node6783;
															assign node6783 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node6787 = (inp[2]) ? 4'b1011 : node6788;
														assign node6788 = (inp[1]) ? 4'b1111 : 4'b1011;
										assign node6792 = (inp[1]) ? node6830 : node6793;
											assign node6793 = (inp[2]) ? node6809 : node6794;
												assign node6794 = (inp[4]) ? node6804 : node6795;
													assign node6795 = (inp[8]) ? node6801 : node6796;
														assign node6796 = (inp[13]) ? node6798 : 4'b1010;
															assign node6798 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node6801 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node6804 = (inp[8]) ? 4'b1110 : node6805;
														assign node6805 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node6809 = (inp[4]) ? node6821 : node6810;
													assign node6810 = (inp[13]) ? node6816 : node6811;
														assign node6811 = (inp[8]) ? 4'b1101 : node6812;
															assign node6812 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6816 = (inp[9]) ? 4'b1010 : node6817;
															assign node6817 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node6821 = (inp[8]) ? node6825 : node6822;
														assign node6822 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node6825 = (inp[13]) ? 4'b1010 : node6826;
															assign node6826 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node6830 = (inp[8]) ? node6858 : node6831;
												assign node6831 = (inp[4]) ? node6845 : node6832;
													assign node6832 = (inp[9]) ? node6838 : node6833;
														assign node6833 = (inp[2]) ? 4'b1011 : node6834;
															assign node6834 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node6838 = (inp[2]) ? node6840 : 4'b1010;
															assign node6840 = (inp[13]) ? 4'b1010 : node6841;
																assign node6841 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node6845 = (inp[2]) ? node6851 : node6846;
														assign node6846 = (inp[9]) ? 4'b1000 : node6847;
															assign node6847 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node6851 = (inp[13]) ? node6855 : node6852;
															assign node6852 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node6855 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node6858 = (inp[4]) ? node6868 : node6859;
													assign node6859 = (inp[2]) ? node6865 : node6860;
														assign node6860 = (inp[13]) ? node6862 : 4'b1101;
															assign node6862 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node6865 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node6868 = (inp[2]) ? node6874 : node6869;
														assign node6869 = (inp[11]) ? 4'b1011 : node6870;
															assign node6870 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node6874 = (inp[9]) ? 4'b1111 : node6875;
															assign node6875 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node6879 = (inp[15]) ? node6985 : node6880;
										assign node6880 = (inp[8]) ? node6952 : node6881;
											assign node6881 = (inp[11]) ? node6923 : node6882;
												assign node6882 = (inp[2]) ? node6908 : node6883;
													assign node6883 = (inp[4]) ? node6895 : node6884;
														assign node6884 = (inp[1]) ? node6890 : node6885;
															assign node6885 = (inp[13]) ? 4'b1110 : node6886;
																assign node6886 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node6890 = (inp[9]) ? 4'b1011 : node6891;
																assign node6891 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node6895 = (inp[1]) ? node6901 : node6896;
															assign node6896 = (inp[13]) ? 4'b1011 : node6897;
																assign node6897 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node6901 = (inp[13]) ? node6905 : node6902;
																assign node6902 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node6905 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6908 = (inp[4]) ? node6914 : node6909;
														assign node6909 = (inp[9]) ? 4'b1011 : node6910;
															assign node6910 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6914 = (inp[1]) ? node6918 : node6915;
															assign node6915 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node6918 = (inp[13]) ? node6920 : 4'b1111;
																assign node6920 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node6923 = (inp[9]) ? node6945 : node6924;
													assign node6924 = (inp[1]) ? node6936 : node6925;
														assign node6925 = (inp[2]) ? node6931 : node6926;
															assign node6926 = (inp[13]) ? 4'b1011 : node6927;
																assign node6927 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node6931 = (inp[4]) ? node6933 : 4'b1111;
																assign node6933 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node6936 = (inp[13]) ? node6940 : node6937;
															assign node6937 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node6940 = (inp[4]) ? node6942 : 4'b1110;
																assign node6942 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node6945 = (inp[4]) ? node6947 : 4'b1111;
														assign node6947 = (inp[2]) ? node6949 : 4'b1010;
															assign node6949 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node6952 = (inp[4]) ? node6974 : node6953;
												assign node6953 = (inp[1]) ? node6965 : node6954;
													assign node6954 = (inp[2]) ? node6960 : node6955;
														assign node6955 = (inp[11]) ? node6957 : 4'b1011;
															assign node6957 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node6960 = (inp[13]) ? node6962 : 4'b1111;
															assign node6962 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node6965 = (inp[2]) ? node6971 : node6966;
														assign node6966 = (inp[11]) ? node6968 : 4'b1110;
															assign node6968 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node6971 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node6974 = (inp[1]) ? node6978 : node6975;
													assign node6975 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node6978 = (inp[2]) ? node6982 : node6979;
														assign node6979 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6982 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node6985 = (inp[2]) ? node7029 : node6986;
											assign node6986 = (inp[13]) ? node7006 : node6987;
												assign node6987 = (inp[1]) ? node6997 : node6988;
													assign node6988 = (inp[4]) ? node6994 : node6989;
														assign node6989 = (inp[11]) ? 4'b1110 : node6990;
															assign node6990 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node6994 = (inp[8]) ? 4'b1101 : 4'b1011;
													assign node6997 = (inp[8]) ? node7003 : node6998;
														assign node6998 = (inp[4]) ? 4'b1110 : node6999;
															assign node6999 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node7003 = (inp[4]) ? 4'b1001 : 4'b1010;
												assign node7006 = (inp[1]) ? node7018 : node7007;
													assign node7007 = (inp[4]) ? node7013 : node7008;
														assign node7008 = (inp[8]) ? 4'b1110 : node7009;
															assign node7009 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node7013 = (inp[9]) ? node7015 : 4'b1110;
															assign node7015 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node7018 = (inp[4]) ? node7022 : node7019;
														assign node7019 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node7022 = (inp[8]) ? node7026 : node7023;
															assign node7023 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node7026 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node7029 = (inp[1]) ? node7053 : node7030;
												assign node7030 = (inp[8]) ? node7046 : node7031;
													assign node7031 = (inp[4]) ? node7039 : node7032;
														assign node7032 = (inp[9]) ? node7036 : node7033;
															assign node7033 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node7036 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node7039 = (inp[13]) ? node7043 : node7040;
															assign node7040 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node7043 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node7046 = (inp[4]) ? 4'b1001 : node7047;
														assign node7047 = (inp[11]) ? 4'b1011 : node7048;
															assign node7048 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node7053 = (inp[13]) ? node7067 : node7054;
													assign node7054 = (inp[8]) ? node7062 : node7055;
														assign node7055 = (inp[4]) ? node7059 : node7056;
															assign node7056 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node7059 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node7062 = (inp[4]) ? node7064 : 4'b1111;
															assign node7064 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node7067 = (inp[11]) ? node7073 : node7068;
														assign node7068 = (inp[8]) ? 4'b1111 : node7069;
															assign node7069 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node7073 = (inp[8]) ? 4'b1110 : node7074;
															assign node7074 = (inp[9]) ? 4'b1110 : 4'b1111;
								assign node7078 = (inp[12]) ? node7228 : node7079;
									assign node7079 = (inp[4]) ? node7165 : node7080;
										assign node7080 = (inp[15]) ? node7114 : node7081;
											assign node7081 = (inp[8]) ? node7103 : node7082;
												assign node7082 = (inp[2]) ? node7092 : node7083;
													assign node7083 = (inp[13]) ? node7089 : node7084;
														assign node7084 = (inp[11]) ? 4'b1010 : node7085;
															assign node7085 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node7089 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node7092 = (inp[13]) ? node7094 : 4'b1111;
														assign node7094 = (inp[1]) ? 4'b1011 : node7095;
															assign node7095 = (inp[9]) ? node7099 : node7096;
																assign node7096 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node7099 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node7103 = (inp[2]) ? node7107 : node7104;
													assign node7104 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node7107 = (inp[1]) ? 4'b1000 : node7108;
														assign node7108 = (inp[13]) ? node7110 : 4'b1101;
															assign node7110 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node7114 = (inp[9]) ? node7140 : node7115;
												assign node7115 = (inp[8]) ? node7129 : node7116;
													assign node7116 = (inp[2]) ? node7122 : node7117;
														assign node7117 = (inp[11]) ? node7119 : 4'b1000;
															assign node7119 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node7122 = (inp[1]) ? node7126 : node7123;
															assign node7123 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node7126 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node7129 = (inp[1]) ? node7135 : node7130;
														assign node7130 = (inp[2]) ? node7132 : 4'b1000;
															assign node7132 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node7135 = (inp[2]) ? node7137 : 4'b1101;
															assign node7137 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node7140 = (inp[11]) ? node7152 : node7141;
													assign node7141 = (inp[1]) ? node7143 : 4'b1001;
														assign node7143 = (inp[8]) ? node7149 : node7144;
															assign node7144 = (inp[13]) ? 4'b1001 : node7145;
																assign node7145 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node7149 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node7152 = (inp[2]) ? node7158 : node7153;
														assign node7153 = (inp[13]) ? node7155 : 4'b1101;
															assign node7155 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node7158 = (inp[1]) ? node7162 : node7159;
															assign node7159 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node7162 = (inp[13]) ? 4'b1000 : 4'b1101;
										assign node7165 = (inp[13]) ? node7203 : node7166;
											assign node7166 = (inp[2]) ? node7188 : node7167;
												assign node7167 = (inp[1]) ? node7173 : node7168;
													assign node7168 = (inp[11]) ? node7170 : 4'b1011;
														assign node7170 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node7173 = (inp[8]) ? node7185 : node7174;
														assign node7174 = (inp[15]) ? node7180 : node7175;
															assign node7175 = (inp[11]) ? node7177 : 4'b1010;
																assign node7177 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node7180 = (inp[9]) ? node7182 : 4'b1011;
																assign node7182 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node7185 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node7188 = (inp[15]) ? node7190 : 4'b1110;
													assign node7190 = (inp[8]) ? node7196 : node7191;
														assign node7191 = (inp[9]) ? node7193 : 4'b1111;
															assign node7193 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node7196 = (inp[1]) ? node7200 : node7197;
															assign node7197 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node7200 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node7203 = (inp[2]) ? node7219 : node7204;
												assign node7204 = (inp[8]) ? node7212 : node7205;
													assign node7205 = (inp[1]) ? 4'b1111 : node7206;
														assign node7206 = (inp[11]) ? node7208 : 4'b1110;
															assign node7208 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node7212 = (inp[1]) ? 4'b1111 : node7213;
														assign node7213 = (inp[15]) ? node7215 : 4'b1011;
															assign node7215 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node7219 = (inp[1]) ? node7223 : node7220;
													assign node7220 = (inp[8]) ? 4'b1110 : 4'b1011;
													assign node7223 = (inp[15]) ? 4'b1011 : node7224;
														assign node7224 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node7228 = (inp[4]) ? node7312 : node7229;
										assign node7229 = (inp[8]) ? node7281 : node7230;
											assign node7230 = (inp[15]) ? node7258 : node7231;
												assign node7231 = (inp[11]) ? node7243 : node7232;
													assign node7232 = (inp[2]) ? 4'b1101 : node7233;
														assign node7233 = (inp[13]) ? 4'b1000 : node7234;
															assign node7234 = (inp[9]) ? node7238 : node7235;
																assign node7235 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node7238 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node7243 = (inp[2]) ? node7253 : node7244;
														assign node7244 = (inp[13]) ? node7250 : node7245;
															assign node7245 = (inp[9]) ? node7247 : 4'b1100;
																assign node7247 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7250 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7253 = (inp[1]) ? node7255 : 4'b1100;
															assign node7255 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node7258 = (inp[11]) ? node7270 : node7259;
													assign node7259 = (inp[13]) ? node7263 : node7260;
														assign node7260 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node7263 = (inp[2]) ? node7267 : node7264;
															assign node7264 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node7267 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node7270 = (inp[13]) ? node7276 : node7271;
														assign node7271 = (inp[9]) ? 4'b1110 : node7272;
															assign node7272 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node7276 = (inp[2]) ? 4'b1011 : node7277;
															assign node7277 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node7281 = (inp[11]) ? node7299 : node7282;
												assign node7282 = (inp[1]) ? node7292 : node7283;
													assign node7283 = (inp[13]) ? 4'b1110 : node7284;
														assign node7284 = (inp[9]) ? 4'b1110 : node7285;
															assign node7285 = (inp[2]) ? 4'b1010 : node7286;
																assign node7286 = (inp[15]) ? 4'b1010 : 4'b1111;
													assign node7292 = (inp[15]) ? node7296 : node7293;
														assign node7293 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node7296 = (inp[2]) ? 4'b1010 : 4'b1111;
												assign node7299 = (inp[15]) ? node7307 : node7300;
													assign node7300 = (inp[2]) ? 4'b1111 : node7301;
														assign node7301 = (inp[1]) ? node7303 : 4'b1111;
															assign node7303 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node7307 = (inp[1]) ? node7309 : 4'b1011;
														assign node7309 = (inp[2]) ? 4'b1011 : 4'b1110;
										assign node7312 = (inp[13]) ? node7354 : node7313;
											assign node7313 = (inp[2]) ? node7333 : node7314;
												assign node7314 = (inp[1]) ? node7324 : node7315;
													assign node7315 = (inp[8]) ? 4'b1000 : node7316;
														assign node7316 = (inp[11]) ? node7318 : 4'b1001;
															assign node7318 = (inp[15]) ? 4'b1000 : node7319;
																assign node7319 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7324 = (inp[8]) ? node7328 : node7325;
														assign node7325 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node7328 = (inp[15]) ? node7330 : 4'b1101;
															assign node7330 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node7333 = (inp[1]) ? node7341 : node7334;
													assign node7334 = (inp[11]) ? 4'b1101 : node7335;
														assign node7335 = (inp[8]) ? node7337 : 4'b1100;
															assign node7337 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node7341 = (inp[8]) ? node7349 : node7342;
														assign node7342 = (inp[9]) ? node7346 : node7343;
															assign node7343 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node7346 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node7349 = (inp[15]) ? node7351 : 4'b1000;
															assign node7351 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node7354 = (inp[2]) ? node7368 : node7355;
												assign node7355 = (inp[11]) ? node7363 : node7356;
													assign node7356 = (inp[9]) ? node7358 : 4'b1101;
														assign node7358 = (inp[8]) ? 4'b1101 : node7359;
															assign node7359 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node7363 = (inp[1]) ? 4'b1101 : node7364;
														assign node7364 = (inp[8]) ? 4'b1001 : 4'b1101;
												assign node7368 = (inp[8]) ? node7376 : node7369;
													assign node7369 = (inp[15]) ? node7371 : 4'b1000;
														assign node7371 = (inp[9]) ? node7373 : 4'b1000;
															assign node7373 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node7376 = (inp[1]) ? 4'b1001 : 4'b1101;
						assign node7379 = (inp[10]) ? node8115 : node7380;
							assign node7380 = (inp[11]) ? node7732 : node7381;
								assign node7381 = (inp[8]) ? node7593 : node7382;
									assign node7382 = (inp[9]) ? node7500 : node7383;
										assign node7383 = (inp[13]) ? node7441 : node7384;
											assign node7384 = (inp[15]) ? node7404 : node7385;
												assign node7385 = (inp[4]) ? node7395 : node7386;
													assign node7386 = (inp[1]) ? node7388 : 4'b1000;
														assign node7388 = (inp[2]) ? node7392 : node7389;
															assign node7389 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node7392 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node7395 = (inp[12]) ? node7397 : 4'b1110;
														assign node7397 = (inp[7]) ? node7401 : node7398;
															assign node7398 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node7401 = (inp[1]) ? 4'b1100 : 4'b1001;
												assign node7404 = (inp[2]) ? node7424 : node7405;
													assign node7405 = (inp[7]) ? node7413 : node7406;
														assign node7406 = (inp[12]) ? node7408 : 4'b1101;
															assign node7408 = (inp[4]) ? node7410 : 4'b1100;
																assign node7410 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node7413 = (inp[1]) ? node7419 : node7414;
															assign node7414 = (inp[12]) ? node7416 : 4'b1011;
																assign node7416 = (inp[4]) ? 4'b1000 : 4'b1011;
															assign node7419 = (inp[4]) ? 4'b1011 : node7420;
																assign node7420 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node7424 = (inp[7]) ? node7430 : node7425;
														assign node7425 = (inp[12]) ? 4'b1001 : node7426;
															assign node7426 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node7430 = (inp[1]) ? node7438 : node7431;
															assign node7431 = (inp[12]) ? node7435 : node7432;
																assign node7432 = (inp[4]) ? 4'b1110 : 4'b1001;
																assign node7435 = (inp[4]) ? 4'b1101 : 4'b1110;
															assign node7438 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node7441 = (inp[2]) ? node7471 : node7442;
												assign node7442 = (inp[1]) ? node7460 : node7443;
													assign node7443 = (inp[12]) ? node7453 : node7444;
														assign node7444 = (inp[15]) ? node7448 : node7445;
															assign node7445 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node7448 = (inp[4]) ? 4'b1000 : node7449;
																assign node7449 = (inp[7]) ? 4'b1000 : 4'b1111;
														assign node7453 = (inp[4]) ? 4'b1101 : node7454;
															assign node7454 = (inp[15]) ? node7456 : 4'b1001;
																assign node7456 = (inp[7]) ? 4'b1110 : 4'b1000;
													assign node7460 = (inp[15]) ? node7462 : 4'b1110;
														assign node7462 = (inp[7]) ? node7464 : 4'b1000;
															assign node7464 = (inp[4]) ? node7468 : node7465;
																assign node7465 = (inp[12]) ? 4'b1110 : 4'b1100;
																assign node7468 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node7471 = (inp[4]) ? node7487 : node7472;
													assign node7472 = (inp[12]) ? node7478 : node7473;
														assign node7473 = (inp[1]) ? 4'b1011 : node7474;
															assign node7474 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node7478 = (inp[1]) ? node7484 : node7479;
															assign node7479 = (inp[15]) ? 4'b1100 : node7480;
																assign node7480 = (inp[7]) ? 4'b1100 : 4'b1011;
															assign node7484 = (inp[15]) ? 4'b1011 : 4'b1110;
													assign node7487 = (inp[1]) ? node7493 : node7488;
														assign node7488 = (inp[12]) ? node7490 : 4'b1101;
															assign node7490 = (inp[15]) ? 4'b1010 : 4'b1001;
														assign node7493 = (inp[12]) ? node7497 : node7494;
															assign node7494 = (inp[7]) ? 4'b1010 : 4'b1100;
															assign node7497 = (inp[7]) ? 4'b1000 : 4'b1010;
										assign node7500 = (inp[4]) ? node7546 : node7501;
											assign node7501 = (inp[2]) ? node7525 : node7502;
												assign node7502 = (inp[13]) ? node7510 : node7503;
													assign node7503 = (inp[12]) ? 4'b1010 : node7504;
														assign node7504 = (inp[1]) ? node7506 : 4'b1101;
															assign node7506 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node7510 = (inp[7]) ? node7518 : node7511;
														assign node7511 = (inp[15]) ? node7515 : node7512;
															assign node7512 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node7515 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node7518 = (inp[12]) ? 4'b1001 : node7519;
															assign node7519 = (inp[15]) ? node7521 : 4'b1111;
																assign node7521 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node7525 = (inp[7]) ? node7535 : node7526;
													assign node7526 = (inp[12]) ? node7532 : node7527;
														assign node7527 = (inp[13]) ? 4'b1000 : node7528;
															assign node7528 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node7532 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node7535 = (inp[12]) ? node7539 : node7536;
														assign node7536 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node7539 = (inp[15]) ? node7543 : node7540;
															assign node7540 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node7543 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node7546 = (inp[7]) ? node7566 : node7547;
												assign node7547 = (inp[12]) ? node7561 : node7548;
													assign node7548 = (inp[15]) ? node7556 : node7549;
														assign node7549 = (inp[2]) ? node7553 : node7550;
															assign node7550 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node7553 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node7556 = (inp[2]) ? node7558 : 4'b1001;
															assign node7558 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node7561 = (inp[13]) ? node7563 : 4'b1111;
														assign node7563 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node7566 = (inp[12]) ? node7582 : node7567;
													assign node7567 = (inp[15]) ? node7575 : node7568;
														assign node7568 = (inp[13]) ? node7572 : node7569;
															assign node7569 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node7572 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node7575 = (inp[13]) ? node7579 : node7576;
															assign node7576 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node7579 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node7582 = (inp[1]) ? node7590 : node7583;
														assign node7583 = (inp[2]) ? 4'b1100 : node7584;
															assign node7584 = (inp[13]) ? 4'b1100 : node7585;
																assign node7585 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node7590 = (inp[2]) ? 4'b1001 : 4'b1101;
									assign node7593 = (inp[2]) ? node7663 : node7594;
										assign node7594 = (inp[1]) ? node7632 : node7595;
											assign node7595 = (inp[12]) ? node7611 : node7596;
												assign node7596 = (inp[4]) ? node7604 : node7597;
													assign node7597 = (inp[7]) ? 4'b1001 : node7598;
														assign node7598 = (inp[15]) ? node7600 : 4'b1001;
															assign node7600 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node7604 = (inp[7]) ? 4'b1011 : node7605;
														assign node7605 = (inp[15]) ? node7607 : 4'b1011;
															assign node7607 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node7611 = (inp[4]) ? node7627 : node7612;
													assign node7612 = (inp[9]) ? node7620 : node7613;
														assign node7613 = (inp[13]) ? 4'b1011 : node7614;
															assign node7614 = (inp[15]) ? 4'b1111 : node7615;
																assign node7615 = (inp[7]) ? 4'b1111 : 4'b1011;
														assign node7620 = (inp[15]) ? 4'b1110 : node7621;
															assign node7621 = (inp[7]) ? node7623 : 4'b1011;
																assign node7623 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node7627 = (inp[15]) ? node7629 : 4'b1000;
														assign node7629 = (inp[7]) ? 4'b1000 : 4'b1101;
											assign node7632 = (inp[12]) ? node7646 : node7633;
												assign node7633 = (inp[4]) ? node7641 : node7634;
													assign node7634 = (inp[15]) ? node7636 : 4'b1101;
														assign node7636 = (inp[7]) ? node7638 : 4'b1101;
															assign node7638 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node7641 = (inp[15]) ? node7643 : 4'b1111;
														assign node7643 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node7646 = (inp[4]) ? node7654 : node7647;
													assign node7647 = (inp[15]) ? node7651 : node7648;
														assign node7648 = (inp[7]) ? 4'b1011 : 4'b1110;
														assign node7651 = (inp[7]) ? 4'b1111 : 4'b1011;
													assign node7654 = (inp[7]) ? node7658 : node7655;
														assign node7655 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node7658 = (inp[13]) ? 4'b1101 : node7659;
															assign node7659 = (inp[15]) ? 4'b1100 : 4'b1101;
										assign node7663 = (inp[1]) ? node7703 : node7664;
											assign node7664 = (inp[15]) ? node7688 : node7665;
												assign node7665 = (inp[13]) ? node7677 : node7666;
													assign node7666 = (inp[7]) ? node7670 : node7667;
														assign node7667 = (inp[4]) ? 4'b1101 : 4'b1111;
														assign node7670 = (inp[12]) ? node7674 : node7671;
															assign node7671 = (inp[4]) ? 4'b1110 : 4'b1101;
															assign node7674 = (inp[4]) ? 4'b1101 : 4'b1010;
													assign node7677 = (inp[4]) ? node7683 : node7678;
														assign node7678 = (inp[12]) ? node7680 : 4'b1100;
															assign node7680 = (inp[7]) ? 4'b1011 : 4'b1110;
														assign node7683 = (inp[7]) ? 4'b1100 : node7684;
															assign node7684 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node7688 = (inp[7]) ? node7696 : node7689;
													assign node7689 = (inp[4]) ? node7693 : node7690;
														assign node7690 = (inp[12]) ? 4'b1011 : 4'b1101;
														assign node7693 = (inp[12]) ? 4'b1001 : 4'b1011;
													assign node7696 = (inp[13]) ? 4'b1101 : node7697;
														assign node7697 = (inp[9]) ? 4'b1100 : node7698;
															assign node7698 = (inp[12]) ? 4'b1100 : 4'b1111;
											assign node7703 = (inp[4]) ? node7719 : node7704;
												assign node7704 = (inp[12]) ? node7712 : node7705;
													assign node7705 = (inp[13]) ? 4'b1000 : node7706;
														assign node7706 = (inp[15]) ? node7708 : 4'b1000;
															assign node7708 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node7712 = (inp[7]) ? node7716 : node7713;
														assign node7713 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node7716 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node7719 = (inp[12]) ? node7725 : node7720;
													assign node7720 = (inp[15]) ? node7722 : 4'b1011;
														assign node7722 = (inp[7]) ? 4'b1011 : 4'b1111;
													assign node7725 = (inp[15]) ? node7729 : node7726;
														assign node7726 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node7729 = (inp[13]) ? 4'b1100 : 4'b1101;
								assign node7732 = (inp[4]) ? node7938 : node7733;
									assign node7733 = (inp[12]) ? node7831 : node7734;
										assign node7734 = (inp[8]) ? node7798 : node7735;
											assign node7735 = (inp[9]) ? node7771 : node7736;
												assign node7736 = (inp[1]) ? node7756 : node7737;
													assign node7737 = (inp[13]) ? node7749 : node7738;
														assign node7738 = (inp[2]) ? node7744 : node7739;
															assign node7739 = (inp[15]) ? node7741 : 4'b1010;
																assign node7741 = (inp[7]) ? 4'b1100 : 4'b1010;
															assign node7744 = (inp[15]) ? 4'b1110 : node7745;
																assign node7745 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node7749 = (inp[15]) ? node7751 : 4'b1100;
															assign node7751 = (inp[7]) ? 4'b1100 : node7752;
																assign node7752 = (inp[2]) ? 4'b1010 : 4'b1111;
													assign node7756 = (inp[2]) ? node7764 : node7757;
														assign node7757 = (inp[13]) ? node7759 : 4'b1010;
															assign node7759 = (inp[15]) ? 4'b1111 : node7760;
																assign node7760 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node7764 = (inp[13]) ? node7766 : 4'b1111;
															assign node7766 = (inp[7]) ? node7768 : 4'b1001;
																assign node7768 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node7771 = (inp[2]) ? node7785 : node7772;
													assign node7772 = (inp[13]) ? 4'b1101 : node7773;
														assign node7773 = (inp[1]) ? node7777 : node7774;
															assign node7774 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node7777 = (inp[15]) ? node7781 : node7778;
																assign node7778 = (inp[7]) ? 4'b1011 : 4'b1001;
																assign node7781 = (inp[7]) ? 4'b1000 : 4'b1011;
													assign node7785 = (inp[13]) ? node7793 : node7786;
														assign node7786 = (inp[15]) ? node7790 : node7787;
															assign node7787 = (inp[7]) ? 4'b1111 : 4'b1101;
															assign node7790 = (inp[1]) ? 4'b1110 : 4'b1000;
														assign node7793 = (inp[15]) ? 4'b1101 : node7794;
															assign node7794 = (inp[7]) ? 4'b1010 : 4'b1000;
											assign node7798 = (inp[2]) ? node7812 : node7799;
												assign node7799 = (inp[1]) ? node7805 : node7800;
													assign node7800 = (inp[13]) ? node7802 : 4'b1000;
														assign node7802 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node7805 = (inp[13]) ? node7807 : 4'b1100;
														assign node7807 = (inp[15]) ? node7809 : 4'b1101;
															assign node7809 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node7812 = (inp[1]) ? node7818 : node7813;
													assign node7813 = (inp[7]) ? 4'b1101 : node7814;
														assign node7814 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node7818 = (inp[9]) ? node7824 : node7819;
														assign node7819 = (inp[13]) ? node7821 : 4'b1001;
															assign node7821 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node7824 = (inp[7]) ? 4'b1000 : node7825;
															assign node7825 = (inp[15]) ? node7827 : 4'b1000;
																assign node7827 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node7831 = (inp[8]) ? node7887 : node7832;
											assign node7832 = (inp[2]) ? node7868 : node7833;
												assign node7833 = (inp[13]) ? node7857 : node7834;
													assign node7834 = (inp[15]) ? node7844 : node7835;
														assign node7835 = (inp[7]) ? node7837 : 4'b1011;
															assign node7837 = (inp[9]) ? node7841 : node7838;
																assign node7838 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node7841 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node7844 = (inp[7]) ? node7852 : node7845;
															assign node7845 = (inp[9]) ? node7849 : node7846;
																assign node7846 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node7849 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node7852 = (inp[9]) ? node7854 : 4'b1010;
																assign node7854 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node7857 = (inp[9]) ? node7861 : node7858;
														assign node7858 = (inp[1]) ? 4'b1111 : 4'b1001;
														assign node7861 = (inp[1]) ? 4'b1010 : node7862;
															assign node7862 = (inp[7]) ? node7864 : 4'b1111;
																assign node7864 = (inp[15]) ? 4'b1111 : 4'b1000;
												assign node7868 = (inp[13]) ? node7876 : node7869;
													assign node7869 = (inp[15]) ? node7873 : node7870;
														assign node7870 = (inp[7]) ? 4'b1000 : 4'b1110;
														assign node7873 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node7876 = (inp[9]) ? 4'b1100 : node7877;
														assign node7877 = (inp[1]) ? node7881 : node7878;
															assign node7878 = (inp[7]) ? 4'b1101 : 4'b1011;
															assign node7881 = (inp[7]) ? node7883 : 4'b1101;
																assign node7883 = (inp[15]) ? 4'b1010 : 4'b1100;
											assign node7887 = (inp[1]) ? node7907 : node7888;
												assign node7888 = (inp[13]) ? node7898 : node7889;
													assign node7889 = (inp[7]) ? 4'b1111 : node7890;
														assign node7890 = (inp[2]) ? node7894 : node7891;
															assign node7891 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node7894 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node7898 = (inp[15]) ? node7902 : node7899;
														assign node7899 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node7902 = (inp[2]) ? node7904 : 4'b1011;
															assign node7904 = (inp[7]) ? 4'b1111 : 4'b1011;
												assign node7907 = (inp[13]) ? node7923 : node7908;
													assign node7908 = (inp[9]) ? node7916 : node7909;
														assign node7909 = (inp[15]) ? node7911 : 4'b1010;
															assign node7911 = (inp[7]) ? node7913 : 4'b1111;
																assign node7913 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node7916 = (inp[15]) ? 4'b1010 : node7917;
															assign node7917 = (inp[7]) ? 4'b1010 : node7918;
																assign node7918 = (inp[2]) ? 4'b1010 : 4'b1111;
													assign node7923 = (inp[7]) ? node7931 : node7924;
														assign node7924 = (inp[9]) ? node7926 : 4'b1110;
															assign node7926 = (inp[15]) ? node7928 : 4'b1011;
																assign node7928 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node7931 = (inp[2]) ? node7935 : node7932;
															assign node7932 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node7935 = (inp[15]) ? 4'b1011 : 4'b1111;
									assign node7938 = (inp[12]) ? node8026 : node7939;
										assign node7939 = (inp[7]) ? node7979 : node7940;
											assign node7940 = (inp[8]) ? node7962 : node7941;
												assign node7941 = (inp[1]) ? node7949 : node7942;
													assign node7942 = (inp[2]) ? node7946 : node7943;
														assign node7943 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node7946 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node7949 = (inp[2]) ? node7951 : 4'b1000;
														assign node7951 = (inp[13]) ? node7959 : node7952;
															assign node7952 = (inp[15]) ? node7956 : node7953;
																assign node7953 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node7956 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node7959 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node7962 = (inp[1]) ? node7968 : node7963;
													assign node7963 = (inp[15]) ? 4'b1110 : node7964;
														assign node7964 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node7968 = (inp[2]) ? node7972 : node7969;
														assign node7969 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node7972 = (inp[15]) ? node7976 : node7973;
															assign node7973 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node7976 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node7979 = (inp[1]) ? node8001 : node7980;
												assign node7980 = (inp[2]) ? node7990 : node7981;
													assign node7981 = (inp[8]) ? node7985 : node7982;
														assign node7982 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node7985 = (inp[13]) ? node7987 : 4'b1011;
															assign node7987 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node7990 = (inp[8]) ? 4'b1110 : node7991;
														assign node7991 = (inp[13]) ? node7997 : node7992;
															assign node7992 = (inp[9]) ? node7994 : 4'b1110;
																assign node7994 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node7997 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node8001 = (inp[13]) ? node8021 : node8002;
													assign node8002 = (inp[15]) ? node8012 : node8003;
														assign node8003 = (inp[8]) ? node8009 : node8004;
															assign node8004 = (inp[2]) ? 4'b1111 : node8005;
																assign node8005 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node8009 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node8012 = (inp[8]) ? node8018 : node8013;
															assign node8013 = (inp[2]) ? node8015 : 4'b1010;
																assign node8015 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node8018 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node8021 = (inp[2]) ? node8023 : 4'b1111;
														assign node8023 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node8026 = (inp[7]) ? node8074 : node8027;
											assign node8027 = (inp[8]) ? node8057 : node8028;
												assign node8028 = (inp[1]) ? node8038 : node8029;
													assign node8029 = (inp[9]) ? node8031 : 4'b1010;
														assign node8031 = (inp[13]) ? 4'b1111 : node8032;
															assign node8032 = (inp[15]) ? node8034 : 4'b1011;
																assign node8034 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node8038 = (inp[2]) ? node8044 : node8039;
														assign node8039 = (inp[9]) ? 4'b1110 : node8040;
															assign node8040 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node8044 = (inp[9]) ? node8052 : node8045;
															assign node8045 = (inp[15]) ? node8049 : node8046;
																assign node8046 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node8049 = (inp[13]) ? 4'b1111 : 4'b1010;
															assign node8052 = (inp[13]) ? 4'b1110 : node8053;
																assign node8053 = (inp[15]) ? 4'b1011 : 4'b1110;
												assign node8057 = (inp[2]) ? node8067 : node8058;
													assign node8058 = (inp[1]) ? node8064 : node8059;
														assign node8059 = (inp[15]) ? node8061 : 4'b1001;
															assign node8061 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node8064 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node8067 = (inp[15]) ? node8071 : node8068;
														assign node8068 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node8071 = (inp[1]) ? 4'b1100 : 4'b1000;
											assign node8074 = (inp[8]) ? node8104 : node8075;
												assign node8075 = (inp[9]) ? node8089 : node8076;
													assign node8076 = (inp[15]) ? node8082 : node8077;
														assign node8077 = (inp[1]) ? 4'b1101 : node8078;
															assign node8078 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node8082 = (inp[2]) ? node8086 : node8083;
															assign node8083 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node8086 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node8089 = (inp[13]) ? node8099 : node8090;
														assign node8090 = (inp[2]) ? node8094 : node8091;
															assign node8091 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node8094 = (inp[15]) ? node8096 : 4'b1100;
																assign node8096 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node8099 = (inp[15]) ? 4'b1001 : node8100;
															assign node8100 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node8104 = (inp[9]) ? node8106 : 4'b1101;
													assign node8106 = (inp[2]) ? node8112 : node8107;
														assign node8107 = (inp[1]) ? 4'b1100 : node8108;
															assign node8108 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node8112 = (inp[1]) ? 4'b1001 : 4'b1101;
							assign node8115 = (inp[9]) ? node8515 : node8116;
								assign node8116 = (inp[8]) ? node8320 : node8117;
									assign node8117 = (inp[4]) ? node8209 : node8118;
										assign node8118 = (inp[15]) ? node8160 : node8119;
											assign node8119 = (inp[13]) ? node8139 : node8120;
												assign node8120 = (inp[12]) ? node8128 : node8121;
													assign node8121 = (inp[2]) ? node8125 : node8122;
														assign node8122 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node8125 = (inp[7]) ? 4'b1111 : 4'b1101;
													assign node8128 = (inp[7]) ? node8134 : node8129;
														assign node8129 = (inp[2]) ? node8131 : 4'b1110;
															assign node8131 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node8134 = (inp[2]) ? node8136 : 4'b1100;
															assign node8136 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node8139 = (inp[2]) ? node8151 : node8140;
													assign node8140 = (inp[12]) ? node8144 : node8141;
														assign node8141 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node8144 = (inp[7]) ? node8148 : node8145;
															assign node8145 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node8148 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node8151 = (inp[12]) ? node8155 : node8152;
														assign node8152 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node8155 = (inp[1]) ? node8157 : 4'b1010;
															assign node8157 = (inp[11]) ? 4'b1101 : 4'b1111;
											assign node8160 = (inp[1]) ? node8184 : node8161;
												assign node8161 = (inp[2]) ? node8169 : node8162;
													assign node8162 = (inp[13]) ? node8164 : 4'b1101;
														assign node8164 = (inp[7]) ? node8166 : 4'b1000;
															assign node8166 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node8169 = (inp[13]) ? node8177 : node8170;
														assign node8170 = (inp[11]) ? node8174 : node8171;
															assign node8171 = (inp[12]) ? 4'b1111 : 4'b1110;
															assign node8174 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node8177 = (inp[7]) ? node8181 : node8178;
															assign node8178 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node8181 = (inp[12]) ? 4'b1010 : 4'b1101;
												assign node8184 = (inp[13]) ? node8200 : node8185;
													assign node8185 = (inp[2]) ? node8193 : node8186;
														assign node8186 = (inp[12]) ? node8190 : node8187;
															assign node8187 = (inp[7]) ? 4'b1000 : 4'b1010;
															assign node8190 = (inp[7]) ? 4'b1011 : 4'b1100;
														assign node8193 = (inp[12]) ? node8197 : node8194;
															assign node8194 = (inp[11]) ? 4'b1110 : 4'b1101;
															assign node8197 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8200 = (inp[12]) ? node8202 : 4'b1101;
														assign node8202 = (inp[7]) ? 4'b1110 : node8203;
															assign node8203 = (inp[2]) ? node8205 : 4'b1000;
																assign node8205 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node8209 = (inp[15]) ? node8263 : node8210;
											assign node8210 = (inp[2]) ? node8240 : node8211;
												assign node8211 = (inp[13]) ? node8221 : node8212;
													assign node8212 = (inp[1]) ? node8214 : 4'b1011;
														assign node8214 = (inp[7]) ? node8218 : node8215;
															assign node8215 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node8218 = (inp[12]) ? 4'b1001 : 4'b1011;
													assign node8221 = (inp[11]) ? node8229 : node8222;
														assign node8222 = (inp[12]) ? node8226 : node8223;
															assign node8223 = (inp[7]) ? 4'b1111 : 4'b1101;
															assign node8226 = (inp[7]) ? 4'b1101 : 4'b1111;
														assign node8229 = (inp[1]) ? node8235 : node8230;
															assign node8230 = (inp[12]) ? 4'b1011 : node8231;
																assign node8231 = (inp[7]) ? 4'b1111 : 4'b1101;
															assign node8235 = (inp[7]) ? node8237 : 4'b1110;
																assign node8237 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node8240 = (inp[13]) ? node8256 : node8241;
													assign node8241 = (inp[11]) ? node8249 : node8242;
														assign node8242 = (inp[1]) ? node8244 : 4'b1101;
															assign node8244 = (inp[7]) ? node8246 : 4'b1110;
																assign node8246 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node8249 = (inp[12]) ? node8253 : node8250;
															assign node8250 = (inp[1]) ? 4'b1110 : 4'b1100;
															assign node8253 = (inp[1]) ? 4'b1100 : 4'b1011;
													assign node8256 = (inp[12]) ? node8260 : node8257;
														assign node8257 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node8260 = (inp[7]) ? 4'b1000 : 4'b1111;
											assign node8263 = (inp[13]) ? node8289 : node8264;
												assign node8264 = (inp[1]) ? node8278 : node8265;
													assign node8265 = (inp[2]) ? node8271 : node8266;
														assign node8266 = (inp[7]) ? node8268 : 4'b1010;
															assign node8268 = (inp[11]) ? 4'b1011 : 4'b1001;
														assign node8271 = (inp[7]) ? node8275 : node8272;
															assign node8272 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node8275 = (inp[11]) ? 4'b1100 : 4'b1111;
													assign node8278 = (inp[7]) ? node8282 : node8279;
														assign node8279 = (inp[11]) ? 4'b1101 : 4'b1111;
														assign node8282 = (inp[2]) ? node8284 : 4'b1010;
															assign node8284 = (inp[11]) ? 4'b1111 : node8285;
																assign node8285 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node8289 = (inp[1]) ? node8309 : node8290;
													assign node8290 = (inp[2]) ? node8302 : node8291;
														assign node8291 = (inp[11]) ? node8297 : node8292;
															assign node8292 = (inp[12]) ? 4'b1100 : node8293;
																assign node8293 = (inp[7]) ? 4'b1111 : 4'b1001;
															assign node8297 = (inp[12]) ? node8299 : 4'b1110;
																assign node8299 = (inp[7]) ? 4'b1101 : 4'b1110;
														assign node8302 = (inp[12]) ? node8304 : 4'b1100;
															assign node8304 = (inp[7]) ? 4'b1001 : node8305;
																assign node8305 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node8309 = (inp[7]) ? node8315 : node8310;
														assign node8310 = (inp[12]) ? node8312 : 4'b1001;
															assign node8312 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node8315 = (inp[2]) ? node8317 : 4'b1101;
															assign node8317 = (inp[12]) ? 4'b1001 : 4'b1011;
									assign node8320 = (inp[11]) ? node8406 : node8321;
										assign node8321 = (inp[2]) ? node8361 : node8322;
											assign node8322 = (inp[1]) ? node8344 : node8323;
												assign node8323 = (inp[4]) ? node8333 : node8324;
													assign node8324 = (inp[12]) ? node8326 : 4'b1000;
														assign node8326 = (inp[15]) ? node8330 : node8327;
															assign node8327 = (inp[7]) ? 4'b1110 : 4'b1010;
															assign node8330 = (inp[7]) ? 4'b1010 : 4'b1111;
													assign node8333 = (inp[12]) ? node8337 : node8334;
														assign node8334 = (inp[7]) ? 4'b1010 : 4'b1111;
														assign node8337 = (inp[7]) ? 4'b1001 : node8338;
															assign node8338 = (inp[15]) ? 4'b1100 : node8339;
																assign node8339 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node8344 = (inp[12]) ? node8350 : node8345;
													assign node8345 = (inp[4]) ? node8347 : 4'b1100;
														assign node8347 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node8350 = (inp[4]) ? node8354 : node8351;
														assign node8351 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node8354 = (inp[7]) ? node8356 : 4'b1000;
															assign node8356 = (inp[15]) ? node8358 : 4'b1100;
																assign node8358 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node8361 = (inp[1]) ? node8385 : node8362;
												assign node8362 = (inp[4]) ? node8378 : node8363;
													assign node8363 = (inp[12]) ? node8373 : node8364;
														assign node8364 = (inp[7]) ? node8366 : 4'b1100;
															assign node8366 = (inp[13]) ? node8370 : node8367;
																assign node8367 = (inp[15]) ? 4'b1101 : 4'b1100;
																assign node8370 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node8373 = (inp[13]) ? 4'b1010 : node8374;
															assign node8374 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node8378 = (inp[12]) ? 4'b1100 : node8379;
														assign node8379 = (inp[15]) ? node8381 : 4'b1110;
															assign node8381 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node8385 = (inp[4]) ? node8391 : node8386;
													assign node8386 = (inp[12]) ? node8388 : 4'b1001;
														assign node8388 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node8391 = (inp[12]) ? node8399 : node8392;
														assign node8392 = (inp[7]) ? node8396 : node8393;
															assign node8393 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node8396 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node8399 = (inp[15]) ? node8401 : 4'b1000;
															assign node8401 = (inp[7]) ? 4'b1001 : node8402;
																assign node8402 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node8406 = (inp[13]) ? node8464 : node8407;
											assign node8407 = (inp[15]) ? node8433 : node8408;
												assign node8408 = (inp[1]) ? node8424 : node8409;
													assign node8409 = (inp[2]) ? node8419 : node8410;
														assign node8410 = (inp[12]) ? node8414 : node8411;
															assign node8411 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node8414 = (inp[4]) ? 4'b1000 : node8415;
																assign node8415 = (inp[7]) ? 4'b1110 : 4'b1011;
														assign node8419 = (inp[4]) ? node8421 : 4'b1011;
															assign node8421 = (inp[12]) ? 4'b1100 : 4'b1111;
													assign node8424 = (inp[2]) ? node8430 : node8425;
														assign node8425 = (inp[4]) ? node8427 : 4'b1101;
															assign node8427 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node8430 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node8433 = (inp[2]) ? node8447 : node8434;
													assign node8434 = (inp[1]) ? node8442 : node8435;
														assign node8435 = (inp[12]) ? node8437 : 4'b1001;
															assign node8437 = (inp[7]) ? node8439 : 4'b1100;
																assign node8439 = (inp[4]) ? 4'b1001 : 4'b1010;
														assign node8442 = (inp[7]) ? 4'b1100 : node8443;
															assign node8443 = (inp[4]) ? 4'b1010 : 4'b1100;
													assign node8447 = (inp[1]) ? node8455 : node8448;
														assign node8448 = (inp[4]) ? node8452 : node8449;
															assign node8449 = (inp[7]) ? 4'b1100 : 4'b1010;
															assign node8452 = (inp[7]) ? 4'b1111 : 4'b1011;
														assign node8455 = (inp[12]) ? node8457 : 4'b1001;
															assign node8457 = (inp[7]) ? node8461 : node8458;
																assign node8458 = (inp[4]) ? 4'b1101 : 4'b1110;
																assign node8461 = (inp[4]) ? 4'b1000 : 4'b1011;
											assign node8464 = (inp[15]) ? node8492 : node8465;
												assign node8465 = (inp[12]) ? node8477 : node8466;
													assign node8466 = (inp[4]) ? node8472 : node8467;
														assign node8467 = (inp[1]) ? node8469 : 4'b1100;
															assign node8469 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node8472 = (inp[2]) ? 4'b1010 : node8473;
															assign node8473 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node8477 = (inp[4]) ? node8487 : node8478;
														assign node8478 = (inp[2]) ? 4'b1110 : node8479;
															assign node8479 = (inp[7]) ? node8483 : node8480;
																assign node8480 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node8483 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node8487 = (inp[1]) ? node8489 : 4'b1001;
															assign node8489 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node8492 = (inp[7]) ? node8506 : node8493;
													assign node8493 = (inp[2]) ? node8501 : node8494;
														assign node8494 = (inp[1]) ? 4'b1001 : node8495;
															assign node8495 = (inp[4]) ? node8497 : 4'b1001;
																assign node8497 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node8501 = (inp[12]) ? node8503 : 4'b1101;
															assign node8503 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node8506 = (inp[12]) ? node8510 : node8507;
														assign node8507 = (inp[4]) ? 4'b1010 : 4'b1001;
														assign node8510 = (inp[4]) ? node8512 : 4'b1110;
															assign node8512 = (inp[2]) ? 4'b1000 : 4'b1100;
								assign node8515 = (inp[4]) ? node8715 : node8516;
									assign node8516 = (inp[12]) ? node8594 : node8517;
										assign node8517 = (inp[8]) ? node8555 : node8518;
											assign node8518 = (inp[2]) ? node8536 : node8519;
												assign node8519 = (inp[13]) ? node8531 : node8520;
													assign node8520 = (inp[15]) ? node8524 : node8521;
														assign node8521 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node8524 = (inp[1]) ? node8528 : node8525;
															assign node8525 = (inp[7]) ? 4'b1100 : 4'b1010;
															assign node8528 = (inp[7]) ? 4'b1001 : 4'b1011;
													assign node8531 = (inp[15]) ? 4'b1111 : node8532;
														assign node8532 = (inp[7]) ? 4'b1110 : 4'b1100;
												assign node8536 = (inp[13]) ? node8548 : node8537;
													assign node8537 = (inp[15]) ? node8543 : node8538;
														assign node8538 = (inp[7]) ? node8540 : 4'b1101;
															assign node8540 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node8543 = (inp[7]) ? node8545 : 4'b1111;
															assign node8545 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node8548 = (inp[15]) ? node8552 : node8549;
														assign node8549 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node8552 = (inp[11]) ? 4'b1001 : 4'b1100;
											assign node8555 = (inp[2]) ? node8575 : node8556;
												assign node8556 = (inp[1]) ? node8562 : node8557;
													assign node8557 = (inp[15]) ? node8559 : 4'b1000;
														assign node8559 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8562 = (inp[13]) ? node8570 : node8563;
														assign node8563 = (inp[7]) ? node8565 : 4'b1100;
															assign node8565 = (inp[11]) ? node8567 : 4'b1101;
																assign node8567 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node8570 = (inp[7]) ? 4'b1100 : node8571;
															assign node8571 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node8575 = (inp[1]) ? 4'b1001 : node8576;
													assign node8576 = (inp[13]) ? node8584 : node8577;
														assign node8577 = (inp[7]) ? node8579 : 4'b1100;
															assign node8579 = (inp[11]) ? 4'b1100 : node8580;
																assign node8580 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node8584 = (inp[15]) ? node8588 : node8585;
															assign node8585 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node8588 = (inp[11]) ? node8590 : 4'b1100;
																assign node8590 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node8594 = (inp[8]) ? node8650 : node8595;
											assign node8595 = (inp[1]) ? node8617 : node8596;
												assign node8596 = (inp[7]) ? node8608 : node8597;
													assign node8597 = (inp[15]) ? 4'b1100 : node8598;
														assign node8598 = (inp[2]) ? node8602 : node8599;
															assign node8599 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node8602 = (inp[13]) ? 4'b1011 : node8603;
																assign node8603 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node8608 = (inp[15]) ? node8612 : node8609;
														assign node8609 = (inp[2]) ? 4'b1000 : 4'b1101;
														assign node8612 = (inp[2]) ? 4'b1011 : node8613;
															assign node8613 = (inp[13]) ? 4'b1110 : 4'b1011;
												assign node8617 = (inp[15]) ? node8635 : node8618;
													assign node8618 = (inp[7]) ? node8624 : node8619;
														assign node8619 = (inp[11]) ? 4'b1010 : node8620;
															assign node8620 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node8624 = (inp[13]) ? node8632 : node8625;
															assign node8625 = (inp[2]) ? node8629 : node8626;
																assign node8626 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node8629 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node8632 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node8635 = (inp[7]) ? node8645 : node8636;
														assign node8636 = (inp[2]) ? node8640 : node8637;
															assign node8637 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node8640 = (inp[13]) ? node8642 : 4'b1000;
																assign node8642 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node8645 = (inp[11]) ? node8647 : 4'b1011;
															assign node8647 = (inp[2]) ? 4'b1111 : 4'b1010;
											assign node8650 = (inp[15]) ? node8686 : node8651;
												assign node8651 = (inp[11]) ? node8669 : node8652;
													assign node8652 = (inp[13]) ? node8664 : node8653;
														assign node8653 = (inp[7]) ? node8657 : node8654;
															assign node8654 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node8657 = (inp[2]) ? node8661 : node8658;
																assign node8658 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node8661 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node8664 = (inp[1]) ? node8666 : 4'b1010;
															assign node8666 = (inp[2]) ? 4'b1111 : 4'b1010;
													assign node8669 = (inp[2]) ? node8675 : node8670;
														assign node8670 = (inp[13]) ? node8672 : 4'b1011;
															assign node8672 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node8675 = (inp[13]) ? node8681 : node8676;
															assign node8676 = (inp[1]) ? node8678 : 4'b1110;
																assign node8678 = (inp[7]) ? 4'b1110 : 4'b1011;
															assign node8681 = (inp[1]) ? node8683 : 4'b1011;
																assign node8683 = (inp[7]) ? 4'b1110 : 4'b1010;
												assign node8686 = (inp[1]) ? node8700 : node8687;
													assign node8687 = (inp[11]) ? 4'b1111 : node8688;
														assign node8688 = (inp[7]) ? node8694 : node8689;
															assign node8689 = (inp[2]) ? 4'b1010 : node8690;
																assign node8690 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node8694 = (inp[2]) ? 4'b1111 : node8695;
																assign node8695 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node8700 = (inp[13]) ? node8710 : node8701;
														assign node8701 = (inp[11]) ? node8705 : node8702;
															assign node8702 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node8705 = (inp[2]) ? 4'b1011 : node8706;
																assign node8706 = (inp[7]) ? 4'b1110 : 4'b1011;
														assign node8710 = (inp[11]) ? node8712 : 4'b1011;
															assign node8712 = (inp[2]) ? 4'b1111 : 4'b1011;
									assign node8715 = (inp[12]) ? node8797 : node8716;
										assign node8716 = (inp[7]) ? node8760 : node8717;
											assign node8717 = (inp[8]) ? node8739 : node8718;
												assign node8718 = (inp[15]) ? node8730 : node8719;
													assign node8719 = (inp[1]) ? node8725 : node8720;
														assign node8720 = (inp[2]) ? 4'b1000 : node8721;
															assign node8721 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node8725 = (inp[13]) ? 4'b1000 : node8726;
															assign node8726 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node8730 = (inp[1]) ? node8734 : node8731;
														assign node8731 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node8734 = (inp[2]) ? 4'b1000 : node8735;
															assign node8735 = (inp[13]) ? 4'b1000 : 4'b1101;
												assign node8739 = (inp[11]) ? node8751 : node8740;
													assign node8740 = (inp[15]) ? node8742 : 4'b1010;
														assign node8742 = (inp[2]) ? node8746 : node8743;
															assign node8743 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node8746 = (inp[1]) ? 4'b1110 : node8747;
																assign node8747 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node8751 = (inp[13]) ? node8755 : node8752;
														assign node8752 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node8755 = (inp[2]) ? 4'b1011 : node8756;
															assign node8756 = (inp[15]) ? 4'b1010 : 4'b1110;
											assign node8760 = (inp[13]) ? node8786 : node8761;
												assign node8761 = (inp[2]) ? node8775 : node8762;
													assign node8762 = (inp[8]) ? node8768 : node8763;
														assign node8763 = (inp[15]) ? node8765 : 4'b1010;
															assign node8765 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node8768 = (inp[1]) ? node8770 : 4'b1010;
															assign node8770 = (inp[15]) ? 4'b1111 : node8771;
																assign node8771 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node8775 = (inp[8]) ? node8781 : node8776;
														assign node8776 = (inp[15]) ? 4'b1110 : node8777;
															assign node8777 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node8781 = (inp[1]) ? node8783 : 4'b1111;
															assign node8783 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node8786 = (inp[2]) ? node8792 : node8787;
													assign node8787 = (inp[8]) ? node8789 : 4'b1110;
														assign node8789 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node8792 = (inp[1]) ? 4'b1010 : node8793;
														assign node8793 = (inp[8]) ? 4'b1111 : 4'b1010;
										assign node8797 = (inp[8]) ? node8851 : node8798;
											assign node8798 = (inp[7]) ? node8830 : node8799;
												assign node8799 = (inp[11]) ? node8821 : node8800;
													assign node8800 = (inp[1]) ? node8810 : node8801;
														assign node8801 = (inp[2]) ? node8807 : node8802;
															assign node8802 = (inp[15]) ? node8804 : 4'b1011;
																assign node8804 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node8807 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node8810 = (inp[15]) ? node8816 : node8811;
															assign node8811 = (inp[13]) ? node8813 : 4'b1111;
																assign node8813 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node8816 = (inp[13]) ? 4'b1010 : node8817;
																assign node8817 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node8821 = (inp[15]) ? node8827 : node8822;
														assign node8822 = (inp[2]) ? node8824 : 4'b1011;
															assign node8824 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node8827 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node8830 = (inp[1]) ? node8842 : node8831;
													assign node8831 = (inp[11]) ? node8837 : node8832;
														assign node8832 = (inp[15]) ? node8834 : 4'b1001;
															assign node8834 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node8837 = (inp[13]) ? node8839 : 4'b1101;
															assign node8839 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node8842 = (inp[13]) ? node8848 : node8843;
														assign node8843 = (inp[15]) ? 4'b1001 : node8844;
															assign node8844 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node8848 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node8851 = (inp[15]) ? node8871 : node8852;
												assign node8852 = (inp[13]) ? node8864 : node8853;
													assign node8853 = (inp[1]) ? node8859 : node8854;
														assign node8854 = (inp[2]) ? 4'b1100 : node8855;
															assign node8855 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8859 = (inp[2]) ? 4'b1001 : node8860;
															assign node8860 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node8864 = (inp[1]) ? node8868 : node8865;
														assign node8865 = (inp[2]) ? 4'b1100 : 4'b1001;
														assign node8868 = (inp[2]) ? 4'b1001 : 4'b1100;
												assign node8871 = (inp[2]) ? node8881 : node8872;
													assign node8872 = (inp[7]) ? node8876 : node8873;
														assign node8873 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node8876 = (inp[11]) ? node8878 : 4'b1001;
															assign node8878 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node8881 = (inp[7]) ? node8889 : node8882;
														assign node8882 = (inp[1]) ? 4'b1101 : node8883;
															assign node8883 = (inp[13]) ? node8885 : 4'b1000;
																assign node8885 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node8889 = (inp[1]) ? 4'b1000 : node8890;
															assign node8890 = (inp[11]) ? 4'b1100 : node8891;
																assign node8891 = (inp[13]) ? 4'b1100 : 4'b1101;
					assign node8896 = (inp[0]) ? node10466 : node8897;
						assign node8897 = (inp[10]) ? node9701 : node8898;
							assign node8898 = (inp[7]) ? node9308 : node8899;
								assign node8899 = (inp[12]) ? node9123 : node8900;
									assign node8900 = (inp[4]) ? node9010 : node8901;
										assign node8901 = (inp[15]) ? node8967 : node8902;
											assign node8902 = (inp[9]) ? node8926 : node8903;
												assign node8903 = (inp[13]) ? node8911 : node8904;
													assign node8904 = (inp[2]) ? node8908 : node8905;
														assign node8905 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node8908 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node8911 = (inp[2]) ? node8919 : node8912;
														assign node8912 = (inp[1]) ? node8916 : node8913;
															assign node8913 = (inp[8]) ? 4'b1100 : 4'b1000;
															assign node8916 = (inp[8]) ? 4'b1001 : 4'b1100;
														assign node8919 = (inp[1]) ? 4'b1001 : node8920;
															assign node8920 = (inp[8]) ? 4'b1001 : node8921;
																assign node8921 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node8926 = (inp[8]) ? node8952 : node8927;
													assign node8927 = (inp[2]) ? node8943 : node8928;
														assign node8928 = (inp[11]) ? node8936 : node8929;
															assign node8929 = (inp[1]) ? node8933 : node8930;
																assign node8930 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node8933 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node8936 = (inp[1]) ? node8940 : node8937;
																assign node8937 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node8940 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node8943 = (inp[1]) ? node8949 : node8944;
															assign node8944 = (inp[11]) ? node8946 : 4'b1100;
																assign node8946 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node8949 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node8952 = (inp[2]) ? node8958 : node8953;
														assign node8953 = (inp[1]) ? 4'b1000 : node8954;
															assign node8954 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node8958 = (inp[1]) ? node8962 : node8959;
															assign node8959 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node8962 = (inp[13]) ? 4'b1101 : node8963;
																assign node8963 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node8967 = (inp[8]) ? node8989 : node8968;
												assign node8968 = (inp[2]) ? node8984 : node8969;
													assign node8969 = (inp[11]) ? node8977 : node8970;
														assign node8970 = (inp[9]) ? node8972 : 4'b1110;
															assign node8972 = (inp[13]) ? node8974 : 4'b1010;
																assign node8974 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node8977 = (inp[1]) ? node8981 : node8978;
															assign node8978 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node8981 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node8984 = (inp[9]) ? 4'b1110 : node8985;
														assign node8985 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node8989 = (inp[1]) ? node9001 : node8990;
													assign node8990 = (inp[2]) ? node8996 : node8991;
														assign node8991 = (inp[13]) ? node8993 : 4'b1000;
															assign node8993 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node8996 = (inp[13]) ? 4'b1100 : node8997;
															assign node8997 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node9001 = (inp[2]) ? node9005 : node9002;
														assign node9002 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node9005 = (inp[11]) ? 4'b1001 : node9006;
															assign node9006 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node9010 = (inp[8]) ? node9064 : node9011;
											assign node9011 = (inp[9]) ? node9043 : node9012;
												assign node9012 = (inp[15]) ? node9024 : node9013;
													assign node9013 = (inp[11]) ? node9017 : node9014;
														assign node9014 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node9017 = (inp[13]) ? 4'b1000 : node9018;
															assign node9018 = (inp[2]) ? node9020 : 4'b1100;
																assign node9020 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node9024 = (inp[13]) ? node9034 : node9025;
														assign node9025 = (inp[1]) ? node9031 : node9026;
															assign node9026 = (inp[2]) ? 4'b1100 : node9027;
																assign node9027 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9031 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node9034 = (inp[1]) ? 4'b1100 : node9035;
															assign node9035 = (inp[2]) ? node9039 : node9036;
																assign node9036 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node9039 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node9043 = (inp[15]) ? node9055 : node9044;
													assign node9044 = (inp[11]) ? node9046 : 4'b1101;
														assign node9046 = (inp[2]) ? node9048 : 4'b1101;
															assign node9048 = (inp[1]) ? node9052 : node9049;
																assign node9049 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node9052 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node9055 = (inp[11]) ? node9061 : node9056;
														assign node9056 = (inp[2]) ? 4'b1101 : node9057;
															assign node9057 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node9061 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node9064 = (inp[11]) ? node9090 : node9065;
												assign node9065 = (inp[1]) ? node9083 : node9066;
													assign node9066 = (inp[9]) ? node9078 : node9067;
														assign node9067 = (inp[15]) ? node9073 : node9068;
															assign node9068 = (inp[2]) ? 4'b1011 : node9069;
																assign node9069 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node9073 = (inp[13]) ? node9075 : 4'b1011;
																assign node9075 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node9078 = (inp[13]) ? node9080 : 4'b1110;
															assign node9080 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node9083 = (inp[15]) ? node9087 : node9084;
														assign node9084 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node9087 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node9090 = (inp[15]) ? node9104 : node9091;
													assign node9091 = (inp[13]) ? node9099 : node9092;
														assign node9092 = (inp[9]) ? 4'b1010 : node9093;
															assign node9093 = (inp[2]) ? 4'b1110 : node9094;
																assign node9094 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node9099 = (inp[2]) ? node9101 : 4'b1110;
															assign node9101 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node9104 = (inp[9]) ? node9112 : node9105;
														assign node9105 = (inp[2]) ? node9109 : node9106;
															assign node9106 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node9109 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node9112 = (inp[13]) ? node9118 : node9113;
															assign node9113 = (inp[1]) ? node9115 : 4'b1110;
																assign node9115 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node9118 = (inp[1]) ? 4'b1010 : node9119;
																assign node9119 = (inp[2]) ? 4'b1111 : 4'b1010;
									assign node9123 = (inp[15]) ? node9225 : node9124;
										assign node9124 = (inp[8]) ? node9184 : node9125;
											assign node9125 = (inp[11]) ? node9161 : node9126;
												assign node9126 = (inp[9]) ? node9146 : node9127;
													assign node9127 = (inp[1]) ? node9137 : node9128;
														assign node9128 = (inp[4]) ? node9130 : 4'b1111;
															assign node9130 = (inp[2]) ? node9134 : node9131;
																assign node9131 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node9134 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node9137 = (inp[4]) ? node9141 : node9138;
															assign node9138 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node9141 = (inp[13]) ? node9143 : 4'b1110;
																assign node9143 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node9146 = (inp[1]) ? node9154 : node9147;
														assign node9147 = (inp[2]) ? 4'b1010 : node9148;
															assign node9148 = (inp[4]) ? 4'b1110 : node9149;
																assign node9149 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node9154 = (inp[13]) ? 4'b1011 : node9155;
															assign node9155 = (inp[4]) ? node9157 : 4'b1111;
																assign node9157 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node9161 = (inp[1]) ? node9175 : node9162;
													assign node9162 = (inp[2]) ? node9170 : node9163;
														assign node9163 = (inp[4]) ? node9167 : node9164;
															assign node9164 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node9167 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node9170 = (inp[13]) ? node9172 : 4'b1010;
															assign node9172 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node9175 = (inp[9]) ? node9181 : node9176;
														assign node9176 = (inp[13]) ? 4'b1111 : node9177;
															assign node9177 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node9181 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node9184 = (inp[4]) ? node9206 : node9185;
												assign node9185 = (inp[13]) ? node9195 : node9186;
													assign node9186 = (inp[2]) ? node9190 : node9187;
														assign node9187 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node9190 = (inp[1]) ? 4'b1010 : node9191;
															assign node9191 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node9195 = (inp[2]) ? node9203 : node9196;
														assign node9196 = (inp[1]) ? node9200 : node9197;
															assign node9197 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node9200 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node9203 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node9206 = (inp[1]) ? node9216 : node9207;
													assign node9207 = (inp[2]) ? node9213 : node9208;
														assign node9208 = (inp[13]) ? 4'b1101 : node9209;
															assign node9209 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node9213 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9216 = (inp[2]) ? node9222 : node9217;
														assign node9217 = (inp[13]) ? node9219 : 4'b1000;
															assign node9219 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9222 = (inp[13]) ? 4'b1100 : 4'b1101;
										assign node9225 = (inp[4]) ? node9269 : node9226;
											assign node9226 = (inp[8]) ? node9254 : node9227;
												assign node9227 = (inp[9]) ? node9239 : node9228;
													assign node9228 = (inp[13]) ? 4'b1101 : node9229;
														assign node9229 = (inp[1]) ? node9233 : node9230;
															assign node9230 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node9233 = (inp[2]) ? 4'b1001 : node9234;
																assign node9234 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9239 = (inp[1]) ? node9245 : node9240;
														assign node9240 = (inp[13]) ? node9242 : 4'b1001;
															assign node9242 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node9245 = (inp[11]) ? 4'b1000 : node9246;
															assign node9246 = (inp[2]) ? node9250 : node9247;
																assign node9247 = (inp[13]) ? 4'b1000 : 4'b1101;
																assign node9250 = (inp[13]) ? 4'b1101 : 4'b1000;
												assign node9254 = (inp[11]) ? node9262 : node9255;
													assign node9255 = (inp[13]) ? node9259 : node9256;
														assign node9256 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node9259 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node9262 = (inp[1]) ? node9266 : node9263;
														assign node9263 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node9266 = (inp[2]) ? 4'b1010 : 4'b1111;
											assign node9269 = (inp[8]) ? node9291 : node9270;
												assign node9270 = (inp[9]) ? node9280 : node9271;
													assign node9271 = (inp[13]) ? node9277 : node9272;
														assign node9272 = (inp[2]) ? node9274 : 4'b1011;
															assign node9274 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node9277 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node9280 = (inp[2]) ? node9288 : node9281;
														assign node9281 = (inp[13]) ? node9285 : node9282;
															assign node9282 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node9285 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node9288 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node9291 = (inp[11]) ? node9303 : node9292;
													assign node9292 = (inp[13]) ? node9296 : node9293;
														assign node9293 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node9296 = (inp[2]) ? node9300 : node9297;
															assign node9297 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node9300 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node9303 = (inp[1]) ? node9305 : 4'b1100;
														assign node9305 = (inp[2]) ? 4'b1000 : 4'b1100;
								assign node9308 = (inp[12]) ? node9490 : node9309;
									assign node9309 = (inp[4]) ? node9395 : node9310;
										assign node9310 = (inp[15]) ? node9354 : node9311;
											assign node9311 = (inp[8]) ? node9343 : node9312;
												assign node9312 = (inp[9]) ? node9328 : node9313;
													assign node9313 = (inp[2]) ? node9319 : node9314;
														assign node9314 = (inp[1]) ? node9316 : 4'b1011;
															assign node9316 = (inp[11]) ? 4'b1111 : 4'b1011;
														assign node9319 = (inp[13]) ? node9325 : node9320;
															assign node9320 = (inp[11]) ? node9322 : 4'b1010;
																assign node9322 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node9325 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node9328 = (inp[2]) ? node9336 : node9329;
														assign node9329 = (inp[11]) ? node9331 : 4'b1010;
															assign node9331 = (inp[1]) ? node9333 : 4'b1111;
																assign node9333 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node9336 = (inp[1]) ? node9338 : 4'b1110;
															assign node9338 = (inp[13]) ? 4'b1011 : node9339;
																assign node9339 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node9343 = (inp[2]) ? node9349 : node9344;
													assign node9344 = (inp[1]) ? node9346 : 4'b1001;
														assign node9346 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9349 = (inp[1]) ? 4'b1000 : node9350;
														assign node9350 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node9354 = (inp[1]) ? node9370 : node9355;
												assign node9355 = (inp[2]) ? node9361 : node9356;
													assign node9356 = (inp[8]) ? 4'b1101 : node9357;
														assign node9357 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node9361 = (inp[13]) ? node9363 : 4'b1000;
														assign node9363 = (inp[8]) ? node9367 : node9364;
															assign node9364 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node9367 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node9370 = (inp[2]) ? node9378 : node9371;
													assign node9371 = (inp[11]) ? node9373 : 4'b1000;
														assign node9373 = (inp[13]) ? node9375 : 4'b1000;
															assign node9375 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node9378 = (inp[13]) ? node9388 : node9379;
														assign node9379 = (inp[8]) ? node9385 : node9380;
															assign node9380 = (inp[9]) ? node9382 : 4'b1001;
																assign node9382 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node9385 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node9388 = (inp[8]) ? 4'b1100 : node9389;
															assign node9389 = (inp[11]) ? node9391 : 4'b1100;
																assign node9391 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node9395 = (inp[9]) ? node9445 : node9396;
											assign node9396 = (inp[15]) ? node9420 : node9397;
												assign node9397 = (inp[11]) ? node9405 : node9398;
													assign node9398 = (inp[2]) ? node9402 : node9399;
														assign node9399 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node9402 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node9405 = (inp[8]) ? node9417 : node9406;
														assign node9406 = (inp[2]) ? node9412 : node9407;
															assign node9407 = (inp[1]) ? 4'b1111 : node9408;
																assign node9408 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node9412 = (inp[13]) ? node9414 : 4'b1011;
																assign node9414 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node9417 = (inp[2]) ? 4'b1111 : 4'b1010;
												assign node9420 = (inp[8]) ? node9434 : node9421;
													assign node9421 = (inp[2]) ? node9427 : node9422;
														assign node9422 = (inp[13]) ? node9424 : 4'b1011;
															assign node9424 = (inp[11]) ? 4'b1011 : 4'b1110;
														assign node9427 = (inp[13]) ? node9429 : 4'b1110;
															assign node9429 = (inp[1]) ? node9431 : 4'b1110;
																assign node9431 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node9434 = (inp[11]) ? node9440 : node9435;
														assign node9435 = (inp[13]) ? 4'b1111 : node9436;
															assign node9436 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node9440 = (inp[2]) ? 4'b1010 : node9441;
															assign node9441 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node9445 = (inp[15]) ? node9467 : node9446;
												assign node9446 = (inp[13]) ? node9454 : node9447;
													assign node9447 = (inp[8]) ? node9449 : 4'b1010;
														assign node9449 = (inp[11]) ? 4'b1111 : node9450;
															assign node9450 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node9454 = (inp[11]) ? node9460 : node9455;
														assign node9455 = (inp[1]) ? 4'b1111 : node9456;
															assign node9456 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node9460 = (inp[2]) ? node9464 : node9461;
															assign node9461 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node9464 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node9467 = (inp[1]) ? node9477 : node9468;
													assign node9468 = (inp[2]) ? node9474 : node9469;
														assign node9469 = (inp[11]) ? node9471 : 4'b1010;
															assign node9471 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node9474 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node9477 = (inp[2]) ? node9487 : node9478;
														assign node9478 = (inp[8]) ? node9484 : node9479;
															assign node9479 = (inp[13]) ? 4'b1110 : node9480;
																assign node9480 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node9484 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node9487 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node9490 = (inp[4]) ? node9592 : node9491;
										assign node9491 = (inp[8]) ? node9551 : node9492;
											assign node9492 = (inp[15]) ? node9522 : node9493;
												assign node9493 = (inp[9]) ? node9507 : node9494;
													assign node9494 = (inp[2]) ? node9502 : node9495;
														assign node9495 = (inp[13]) ? node9499 : node9496;
															assign node9496 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node9499 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node9502 = (inp[1]) ? node9504 : 4'b1100;
															assign node9504 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node9507 = (inp[11]) ? node9515 : node9508;
														assign node9508 = (inp[13]) ? node9510 : 4'b1101;
															assign node9510 = (inp[2]) ? node9512 : 4'b1101;
																assign node9512 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node9515 = (inp[1]) ? 4'b1000 : node9516;
															assign node9516 = (inp[2]) ? 4'b1101 : node9517;
																assign node9517 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node9522 = (inp[1]) ? node9542 : node9523;
													assign node9523 = (inp[11]) ? node9531 : node9524;
														assign node9524 = (inp[9]) ? node9526 : 4'b1011;
															assign node9526 = (inp[13]) ? node9528 : 4'b1010;
																assign node9528 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node9531 = (inp[13]) ? node9539 : node9532;
															assign node9532 = (inp[2]) ? node9536 : node9533;
																assign node9533 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node9536 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node9539 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node9542 = (inp[2]) ? node9548 : node9543;
														assign node9543 = (inp[9]) ? 4'b1011 : node9544;
															assign node9544 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node9548 = (inp[13]) ? 4'b1011 : 4'b1111;
											assign node9551 = (inp[2]) ? node9569 : node9552;
												assign node9552 = (inp[1]) ? node9562 : node9553;
													assign node9553 = (inp[11]) ? node9555 : 4'b1010;
														assign node9555 = (inp[15]) ? node9559 : node9556;
															assign node9556 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node9559 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node9562 = (inp[13]) ? 4'b1111 : node9563;
														assign node9563 = (inp[9]) ? node9565 : 4'b1111;
															assign node9565 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node9569 = (inp[1]) ? node9577 : node9570;
													assign node9570 = (inp[9]) ? node9572 : 4'b1110;
														assign node9572 = (inp[15]) ? node9574 : 4'b1110;
															assign node9574 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node9577 = (inp[13]) ? 4'b1010 : node9578;
														assign node9578 = (inp[9]) ? node9586 : node9579;
															assign node9579 = (inp[15]) ? node9583 : node9580;
																assign node9580 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node9583 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node9586 = (inp[15]) ? node9588 : 4'b1010;
																assign node9588 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node9592 = (inp[13]) ? node9656 : node9593;
											assign node9593 = (inp[15]) ? node9625 : node9594;
												assign node9594 = (inp[9]) ? node9608 : node9595;
													assign node9595 = (inp[1]) ? node9601 : node9596;
														assign node9596 = (inp[8]) ? 4'b1001 : node9597;
															assign node9597 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node9601 = (inp[2]) ? node9605 : node9602;
															assign node9602 = (inp[8]) ? 4'b1100 : 4'b1000;
															assign node9605 = (inp[8]) ? 4'b1001 : 4'b1101;
													assign node9608 = (inp[2]) ? node9618 : node9609;
														assign node9609 = (inp[11]) ? node9611 : 4'b1101;
															assign node9611 = (inp[8]) ? node9615 : node9612;
																assign node9612 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node9615 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node9618 = (inp[8]) ? node9620 : 4'b1100;
															assign node9620 = (inp[1]) ? node9622 : 4'b1100;
																assign node9622 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node9625 = (inp[9]) ? node9643 : node9626;
													assign node9626 = (inp[11]) ? node9632 : node9627;
														assign node9627 = (inp[8]) ? node9629 : 4'b1101;
															assign node9629 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node9632 = (inp[1]) ? node9638 : node9633;
															assign node9633 = (inp[8]) ? node9635 : 4'b1100;
																assign node9635 = (inp[2]) ? 4'b1100 : 4'b1001;
															assign node9638 = (inp[2]) ? 4'b1000 : node9639;
																assign node9639 = (inp[8]) ? 4'b1100 : 4'b1000;
													assign node9643 = (inp[11]) ? node9651 : node9644;
														assign node9644 = (inp[8]) ? node9648 : node9645;
															assign node9645 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node9648 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node9651 = (inp[1]) ? node9653 : 4'b1001;
															assign node9653 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node9656 = (inp[8]) ? node9684 : node9657;
												assign node9657 = (inp[1]) ? node9671 : node9658;
													assign node9658 = (inp[2]) ? node9668 : node9659;
														assign node9659 = (inp[9]) ? node9665 : node9660;
															assign node9660 = (inp[11]) ? 4'b1000 : node9661;
																assign node9661 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node9665 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node9668 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node9671 = (inp[2]) ? node9679 : node9672;
														assign node9672 = (inp[11]) ? node9676 : node9673;
															assign node9673 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node9676 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node9679 = (inp[11]) ? node9681 : 4'b1000;
															assign node9681 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node9684 = (inp[11]) ? node9692 : node9685;
													assign node9685 = (inp[1]) ? node9689 : node9686;
														assign node9686 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node9689 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node9692 = (inp[9]) ? 4'b1100 : node9693;
														assign node9693 = (inp[1]) ? node9697 : node9694;
															assign node9694 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node9697 = (inp[2]) ? 4'b1000 : 4'b1100;
							assign node9701 = (inp[8]) ? node10131 : node9702;
								assign node9702 = (inp[15]) ? node9914 : node9703;
									assign node9703 = (inp[9]) ? node9813 : node9704;
										assign node9704 = (inp[2]) ? node9766 : node9705;
											assign node9705 = (inp[7]) ? node9737 : node9706;
												assign node9706 = (inp[12]) ? node9726 : node9707;
													assign node9707 = (inp[11]) ? node9713 : node9708;
														assign node9708 = (inp[4]) ? 4'b1000 : node9709;
															assign node9709 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node9713 = (inp[4]) ? node9719 : node9714;
															assign node9714 = (inp[1]) ? 4'b1001 : node9715;
																assign node9715 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node9719 = (inp[1]) ? node9723 : node9720;
																assign node9720 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node9723 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node9726 = (inp[1]) ? 4'b1010 : node9727;
														assign node9727 = (inp[4]) ? node9731 : node9728;
															assign node9728 = (inp[11]) ? 4'b1111 : 4'b1011;
															assign node9731 = (inp[13]) ? 4'b1010 : node9732;
																assign node9732 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node9737 = (inp[12]) ? node9753 : node9738;
													assign node9738 = (inp[4]) ? node9744 : node9739;
														assign node9739 = (inp[11]) ? node9741 : 4'b1010;
															assign node9741 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node9744 = (inp[11]) ? node9748 : node9745;
															assign node9745 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node9748 = (inp[1]) ? node9750 : 4'b1110;
																assign node9750 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node9753 = (inp[4]) ? node9759 : node9754;
														assign node9754 = (inp[11]) ? 4'b1000 : node9755;
															assign node9755 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node9759 = (inp[11]) ? node9761 : 4'b1101;
															assign node9761 = (inp[1]) ? node9763 : 4'b1001;
																assign node9763 = (inp[13]) ? 4'b1100 : 4'b1000;
											assign node9766 = (inp[1]) ? node9786 : node9767;
												assign node9767 = (inp[13]) ? node9779 : node9768;
													assign node9768 = (inp[12]) ? node9774 : node9769;
														assign node9769 = (inp[11]) ? 4'b1001 : node9770;
															assign node9770 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node9774 = (inp[4]) ? node9776 : 4'b1101;
															assign node9776 = (inp[7]) ? 4'b1001 : 4'b1011;
													assign node9779 = (inp[12]) ? 4'b1001 : node9780;
														assign node9780 = (inp[11]) ? 4'b1101 : node9781;
															assign node9781 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node9786 = (inp[13]) ? node9796 : node9787;
													assign node9787 = (inp[12]) ? 4'b1110 : node9788;
														assign node9788 = (inp[7]) ? 4'b1111 : node9789;
															assign node9789 = (inp[11]) ? 4'b1101 : node9790;
																assign node9790 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node9796 = (inp[12]) ? node9802 : node9797;
														assign node9797 = (inp[7]) ? 4'b1011 : node9798;
															assign node9798 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9802 = (inp[7]) ? node9808 : node9803;
															assign node9803 = (inp[4]) ? node9805 : 4'b1011;
																assign node9805 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node9808 = (inp[4]) ? 4'b1000 : node9809;
																assign node9809 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node9813 = (inp[12]) ? node9859 : node9814;
											assign node9814 = (inp[7]) ? node9838 : node9815;
												assign node9815 = (inp[11]) ? node9827 : node9816;
													assign node9816 = (inp[4]) ? node9820 : node9817;
														assign node9817 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node9820 = (inp[2]) ? node9824 : node9821;
															assign node9821 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node9824 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node9827 = (inp[1]) ? node9833 : node9828;
														assign node9828 = (inp[13]) ? node9830 : 4'b1000;
															assign node9830 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9833 = (inp[2]) ? node9835 : 4'b1100;
															assign node9835 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node9838 = (inp[4]) ? node9850 : node9839;
													assign node9839 = (inp[13]) ? node9847 : node9840;
														assign node9840 = (inp[2]) ? node9844 : node9841;
															assign node9841 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node9844 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node9847 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node9850 = (inp[2]) ? node9854 : node9851;
														assign node9851 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node9854 = (inp[13]) ? 4'b1111 : node9855;
															assign node9855 = (inp[11]) ? 4'b1011 : 4'b1111;
											assign node9859 = (inp[7]) ? node9897 : node9860;
												assign node9860 = (inp[2]) ? node9876 : node9861;
													assign node9861 = (inp[11]) ? node9867 : node9862;
														assign node9862 = (inp[1]) ? node9864 : 4'b1110;
															assign node9864 = (inp[4]) ? 4'b1110 : 4'b1011;
														assign node9867 = (inp[1]) ? 4'b1010 : node9868;
															assign node9868 = (inp[13]) ? node9872 : node9869;
																assign node9869 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node9872 = (inp[4]) ? 4'b1011 : 4'b1110;
													assign node9876 = (inp[11]) ? node9884 : node9877;
														assign node9877 = (inp[1]) ? node9879 : 4'b1011;
															assign node9879 = (inp[13]) ? 4'b1010 : node9880;
																assign node9880 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9884 = (inp[1]) ? node9890 : node9885;
															assign node9885 = (inp[4]) ? 4'b1110 : node9886;
																assign node9886 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node9890 = (inp[4]) ? node9894 : node9891;
																assign node9891 = (inp[13]) ? 4'b1010 : 4'b1111;
																assign node9894 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node9897 = (inp[4]) ? node9907 : node9898;
													assign node9898 = (inp[11]) ? node9904 : node9899;
														assign node9899 = (inp[13]) ? node9901 : 4'b1100;
															assign node9901 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node9904 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node9907 = (inp[13]) ? 4'b1100 : node9908;
														assign node9908 = (inp[11]) ? node9910 : 4'b1000;
															assign node9910 = (inp[2]) ? 4'b1000 : 4'b1100;
									assign node9914 = (inp[9]) ? node10020 : node9915;
										assign node9915 = (inp[12]) ? node9973 : node9916;
											assign node9916 = (inp[2]) ? node9950 : node9917;
												assign node9917 = (inp[13]) ? node9931 : node9918;
													assign node9918 = (inp[1]) ? node9926 : node9919;
														assign node9919 = (inp[11]) ? node9921 : 4'b1111;
															assign node9921 = (inp[7]) ? node9923 : 4'b1001;
																assign node9923 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node9926 = (inp[4]) ? 4'b1100 : node9927;
															assign node9927 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node9931 = (inp[4]) ? node9941 : node9932;
														assign node9932 = (inp[7]) ? node9936 : node9933;
															assign node9933 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node9936 = (inp[11]) ? node9938 : 4'b1000;
																assign node9938 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node9941 = (inp[7]) ? node9945 : node9942;
															assign node9942 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node9945 = (inp[1]) ? node9947 : 4'b1010;
																assign node9947 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node9950 = (inp[1]) ? node9962 : node9951;
													assign node9951 = (inp[13]) ? node9957 : node9952;
														assign node9952 = (inp[4]) ? node9954 : 4'b1011;
															assign node9954 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node9957 = (inp[4]) ? 4'b1110 : node9958;
															assign node9958 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node9962 = (inp[13]) ? node9968 : node9963;
														assign node9963 = (inp[4]) ? 4'b1000 : node9964;
															assign node9964 = (inp[7]) ? 4'b1000 : 4'b1110;
														assign node9968 = (inp[7]) ? node9970 : 4'b1010;
															assign node9970 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node9973 = (inp[13]) ? node9997 : node9974;
												assign node9974 = (inp[11]) ? node9986 : node9975;
													assign node9975 = (inp[7]) ? node9981 : node9976;
														assign node9976 = (inp[4]) ? node9978 : 4'b1000;
															assign node9978 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node9981 = (inp[1]) ? 4'b1000 : node9982;
															assign node9982 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node9986 = (inp[1]) ? node9992 : node9987;
														assign node9987 = (inp[2]) ? 4'b1111 : node9988;
															assign node9988 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9992 = (inp[7]) ? node9994 : 4'b1001;
															assign node9994 = (inp[4]) ? 4'b1001 : 4'b1111;
												assign node9997 = (inp[4]) ? node10011 : node9998;
													assign node9998 = (inp[7]) ? node10004 : node9999;
														assign node9999 = (inp[1]) ? node10001 : 4'b1001;
															assign node10001 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node10004 = (inp[11]) ? node10006 : 4'b1111;
															assign node10006 = (inp[1]) ? node10008 : 4'b1010;
																assign node10008 = (inp[2]) ? 4'b1010 : 4'b1111;
													assign node10011 = (inp[7]) ? node10013 : 4'b1111;
														assign node10013 = (inp[2]) ? node10017 : node10014;
															assign node10014 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node10017 = (inp[11]) ? 4'b1100 : 4'b1001;
										assign node10020 = (inp[2]) ? node10072 : node10021;
											assign node10021 = (inp[7]) ? node10043 : node10022;
												assign node10022 = (inp[4]) ? node10034 : node10023;
													assign node10023 = (inp[12]) ? node10025 : 4'b1011;
														assign node10025 = (inp[13]) ? node10031 : node10026;
															assign node10026 = (inp[1]) ? node10028 : 4'b1000;
																assign node10028 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node10031 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node10034 = (inp[12]) ? 4'b1011 : node10035;
														assign node10035 = (inp[1]) ? 4'b1101 : node10036;
															assign node10036 = (inp[13]) ? 4'b1101 : node10037;
																assign node10037 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node10043 = (inp[4]) ? node10059 : node10044;
													assign node10044 = (inp[12]) ? node10050 : node10045;
														assign node10045 = (inp[13]) ? node10047 : 4'b1101;
															assign node10047 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node10050 = (inp[11]) ? node10056 : node10051;
															assign node10051 = (inp[13]) ? 4'b1111 : node10052;
																assign node10052 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node10056 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node10059 = (inp[12]) ? node10065 : node10060;
														assign node10060 = (inp[1]) ? node10062 : 4'b1011;
															assign node10062 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node10065 = (inp[1]) ? node10067 : 4'b1000;
															assign node10067 = (inp[13]) ? 4'b1101 : node10068;
																assign node10068 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node10072 = (inp[4]) ? node10112 : node10073;
												assign node10073 = (inp[13]) ? node10093 : node10074;
													assign node10074 = (inp[11]) ? node10084 : node10075;
														assign node10075 = (inp[1]) ? 4'b1001 : node10076;
															assign node10076 = (inp[12]) ? node10080 : node10077;
																assign node10077 = (inp[7]) ? 4'b1000 : 4'b1011;
																assign node10080 = (inp[7]) ? 4'b1011 : 4'b1101;
														assign node10084 = (inp[7]) ? 4'b1000 : node10085;
															assign node10085 = (inp[12]) ? node10089 : node10086;
																assign node10086 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node10089 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node10093 = (inp[11]) ? node10103 : node10094;
														assign node10094 = (inp[7]) ? node10100 : node10095;
															assign node10095 = (inp[12]) ? node10097 : 4'b1011;
																assign node10097 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node10100 = (inp[1]) ? 4'b1100 : 4'b1110;
														assign node10103 = (inp[7]) ? node10107 : node10104;
															assign node10104 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node10107 = (inp[12]) ? node10109 : 4'b1101;
																assign node10109 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node10112 = (inp[13]) ? node10122 : node10113;
													assign node10113 = (inp[12]) ? node10119 : node10114;
														assign node10114 = (inp[7]) ? 4'b1110 : node10115;
															assign node10115 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node10119 = (inp[7]) ? 4'b1100 : 4'b1110;
													assign node10122 = (inp[11]) ? node10128 : node10123;
														assign node10123 = (inp[12]) ? node10125 : 4'b1000;
															assign node10125 = (inp[1]) ? 4'b1000 : 4'b1010;
														assign node10128 = (inp[12]) ? 4'b1101 : 4'b1001;
								assign node10131 = (inp[11]) ? node10317 : node10132;
									assign node10132 = (inp[7]) ? node10218 : node10133;
										assign node10133 = (inp[15]) ? node10177 : node10134;
											assign node10134 = (inp[2]) ? node10156 : node10135;
												assign node10135 = (inp[12]) ? node10143 : node10136;
													assign node10136 = (inp[4]) ? node10138 : 4'b1101;
														assign node10138 = (inp[1]) ? 4'b1010 : node10139;
															assign node10139 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node10143 = (inp[4]) ? node10151 : node10144;
														assign node10144 = (inp[1]) ? node10148 : node10145;
															assign node10145 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node10148 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node10151 = (inp[1]) ? node10153 : 4'b1100;
															assign node10153 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node10156 = (inp[1]) ? node10166 : node10157;
													assign node10157 = (inp[4]) ? node10161 : node10158;
														assign node10158 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node10161 = (inp[12]) ? 4'b1000 : node10162;
															assign node10162 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node10166 = (inp[12]) ? node10172 : node10167;
														assign node10167 = (inp[4]) ? node10169 : 4'b1100;
															assign node10169 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node10172 = (inp[4]) ? 4'b1101 : node10173;
															assign node10173 = (inp[13]) ? 4'b1010 : 4'b1011;
											assign node10177 = (inp[13]) ? node10199 : node10178;
												assign node10178 = (inp[1]) ? node10194 : node10179;
													assign node10179 = (inp[2]) ? node10185 : node10180;
														assign node10180 = (inp[4]) ? 4'b1010 : node10181;
															assign node10181 = (inp[9]) ? 4'b1011 : 4'b1001;
														assign node10185 = (inp[9]) ? 4'b1111 : node10186;
															assign node10186 = (inp[4]) ? node10190 : node10187;
																assign node10187 = (inp[12]) ? 4'b1110 : 4'b1100;
																assign node10190 = (inp[12]) ? 4'b1100 : 4'b1111;
													assign node10194 = (inp[12]) ? 4'b1010 : node10195;
														assign node10195 = (inp[4]) ? 4'b1110 : 4'b1100;
												assign node10199 = (inp[1]) ? node10209 : node10200;
													assign node10200 = (inp[2]) ? node10206 : node10201;
														assign node10201 = (inp[12]) ? node10203 : 4'b1011;
															assign node10203 = (inp[9]) ? 4'b1000 : 4'b1011;
														assign node10206 = (inp[9]) ? 4'b1101 : 4'b1111;
													assign node10209 = (inp[2]) ? node10213 : node10210;
														assign node10210 = (inp[9]) ? 4'b1110 : 4'b1101;
														assign node10213 = (inp[9]) ? node10215 : 4'b1000;
															assign node10215 = (inp[4]) ? 4'b1001 : 4'b1011;
										assign node10218 = (inp[13]) ? node10280 : node10219;
											assign node10219 = (inp[15]) ? node10249 : node10220;
												assign node10220 = (inp[2]) ? node10234 : node10221;
													assign node10221 = (inp[1]) ? node10227 : node10222;
														assign node10222 = (inp[4]) ? 4'b1011 : node10223;
															assign node10223 = (inp[12]) ? 4'b1011 : 4'b1000;
														assign node10227 = (inp[4]) ? node10231 : node10228;
															assign node10228 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node10231 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node10234 = (inp[1]) ? node10242 : node10235;
														assign node10235 = (inp[9]) ? node10237 : 4'b1101;
															assign node10237 = (inp[12]) ? 4'b1101 : node10238;
																assign node10238 = (inp[4]) ? 4'b1110 : 4'b1101;
														assign node10242 = (inp[9]) ? 4'b1011 : node10243;
															assign node10243 = (inp[12]) ? node10245 : 4'b1001;
																assign node10245 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node10249 = (inp[12]) ? node10265 : node10250;
													assign node10250 = (inp[4]) ? node10258 : node10251;
														assign node10251 = (inp[2]) ? node10255 : node10252;
															assign node10252 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node10255 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node10258 = (inp[1]) ? node10262 : node10259;
															assign node10259 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node10262 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node10265 = (inp[4]) ? node10273 : node10266;
														assign node10266 = (inp[2]) ? node10270 : node10267;
															assign node10267 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node10270 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node10273 = (inp[9]) ? node10275 : 4'b1000;
															assign node10275 = (inp[1]) ? node10277 : 4'b1100;
																assign node10277 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node10280 = (inp[1]) ? node10306 : node10281;
												assign node10281 = (inp[2]) ? node10291 : node10282;
													assign node10282 = (inp[4]) ? node10288 : node10283;
														assign node10283 = (inp[12]) ? 4'b1011 : node10284;
															assign node10284 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node10288 = (inp[12]) ? 4'b1000 : 4'b1011;
													assign node10291 = (inp[9]) ? node10295 : node10292;
														assign node10292 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node10295 = (inp[15]) ? node10303 : node10296;
															assign node10296 = (inp[12]) ? node10300 : node10297;
																assign node10297 = (inp[4]) ? 4'b1111 : 4'b1101;
																assign node10300 = (inp[4]) ? 4'b1100 : 4'b1110;
															assign node10303 = (inp[12]) ? 4'b1111 : 4'b1110;
												assign node10306 = (inp[2]) ? node10312 : node10307;
													assign node10307 = (inp[9]) ? node10309 : 4'b1001;
														assign node10309 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node10312 = (inp[4]) ? node10314 : 4'b1011;
														assign node10314 = (inp[12]) ? 4'b1001 : 4'b1011;
									assign node10317 = (inp[4]) ? node10387 : node10318;
										assign node10318 = (inp[12]) ? node10366 : node10319;
											assign node10319 = (inp[9]) ? node10341 : node10320;
												assign node10320 = (inp[15]) ? node10332 : node10321;
													assign node10321 = (inp[13]) ? node10325 : node10322;
														assign node10322 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node10325 = (inp[2]) ? node10327 : 4'b1101;
															assign node10327 = (inp[7]) ? 4'b1001 : node10328;
																assign node10328 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node10332 = (inp[2]) ? node10336 : node10333;
														assign node10333 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node10336 = (inp[13]) ? 4'b1101 : node10337;
															assign node10337 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node10341 = (inp[7]) ? node10355 : node10342;
													assign node10342 = (inp[2]) ? node10348 : node10343;
														assign node10343 = (inp[1]) ? 4'b1001 : node10344;
															assign node10344 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node10348 = (inp[13]) ? 4'b1000 : node10349;
															assign node10349 = (inp[15]) ? node10351 : 4'b1101;
																assign node10351 = (inp[1]) ? 4'b1000 : 4'b1101;
													assign node10355 = (inp[2]) ? node10363 : node10356;
														assign node10356 = (inp[15]) ? node10360 : node10357;
															assign node10357 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node10360 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node10363 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node10366 = (inp[2]) ? node10378 : node10367;
												assign node10367 = (inp[1]) ? 4'b1110 : node10368;
													assign node10368 = (inp[15]) ? node10374 : node10369;
														assign node10369 = (inp[9]) ? 4'b1011 : node10370;
															assign node10370 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node10374 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node10378 = (inp[1]) ? node10380 : 4'b1111;
													assign node10380 = (inp[15]) ? 4'b1011 : node10381;
														assign node10381 = (inp[9]) ? 4'b1011 : node10382;
															assign node10382 = (inp[13]) ? 4'b1011 : 4'b1010;
										assign node10387 = (inp[12]) ? node10425 : node10388;
											assign node10388 = (inp[7]) ? node10412 : node10389;
												assign node10389 = (inp[1]) ? node10405 : node10390;
													assign node10390 = (inp[9]) ? node10396 : node10391;
														assign node10391 = (inp[15]) ? 4'b1011 : node10392;
															assign node10392 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node10396 = (inp[2]) ? node10400 : node10397;
															assign node10397 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node10400 = (inp[15]) ? node10402 : 4'b1011;
																assign node10402 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node10405 = (inp[13]) ? 4'b1111 : node10406;
														assign node10406 = (inp[15]) ? 4'b1010 : node10407;
															assign node10407 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node10412 = (inp[1]) ? node10418 : node10413;
													assign node10413 = (inp[2]) ? 4'b1110 : node10414;
														assign node10414 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node10418 = (inp[2]) ? 4'b1011 : node10419;
														assign node10419 = (inp[15]) ? 4'b1111 : node10420;
															assign node10420 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node10425 = (inp[13]) ? node10449 : node10426;
												assign node10426 = (inp[1]) ? node10438 : node10427;
													assign node10427 = (inp[9]) ? 4'b1101 : node10428;
														assign node10428 = (inp[2]) ? node10434 : node10429;
															assign node10429 = (inp[15]) ? 4'b1000 : node10430;
																assign node10430 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node10434 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node10438 = (inp[15]) ? node10446 : node10439;
														assign node10439 = (inp[2]) ? node10443 : node10440;
															assign node10440 = (inp[7]) ? 4'b1100 : 4'b1001;
															assign node10443 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node10446 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node10449 = (inp[9]) ? node10457 : node10450;
													assign node10450 = (inp[2]) ? node10454 : node10451;
														assign node10451 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node10454 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node10457 = (inp[15]) ? node10459 : 4'b1101;
														assign node10459 = (inp[1]) ? node10463 : node10460;
															assign node10460 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node10463 = (inp[2]) ? 4'b1001 : 4'b1101;
						assign node10466 = (inp[10]) ? node11282 : node10467;
							assign node10467 = (inp[11]) ? node10903 : node10468;
								assign node10468 = (inp[9]) ? node10666 : node10469;
									assign node10469 = (inp[1]) ? node10575 : node10470;
										assign node10470 = (inp[2]) ? node10520 : node10471;
											assign node10471 = (inp[12]) ? node10499 : node10472;
												assign node10472 = (inp[7]) ? node10490 : node10473;
													assign node10473 = (inp[15]) ? node10483 : node10474;
														assign node10474 = (inp[8]) ? node10480 : node10475;
															assign node10475 = (inp[13]) ? 4'b1001 : node10476;
																assign node10476 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node10480 = (inp[4]) ? 4'b1110 : 4'b1101;
														assign node10483 = (inp[8]) ? node10487 : node10484;
															assign node10484 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node10487 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node10490 = (inp[4]) ? node10496 : node10491;
														assign node10491 = (inp[15]) ? 4'b1100 : node10492;
															assign node10492 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node10496 = (inp[8]) ? 4'b1011 : 4'b1110;
												assign node10499 = (inp[4]) ? node10509 : node10500;
													assign node10500 = (inp[8]) ? node10506 : node10501;
														assign node10501 = (inp[7]) ? 4'b1000 : node10502;
															assign node10502 = (inp[15]) ? 4'b1100 : 4'b1111;
														assign node10506 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node10509 = (inp[8]) ? node10515 : node10510;
														assign node10510 = (inp[7]) ? node10512 : 4'b1010;
															assign node10512 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node10515 = (inp[15]) ? 4'b1000 : node10516;
															assign node10516 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node10520 = (inp[8]) ? node10544 : node10521;
												assign node10521 = (inp[7]) ? node10533 : node10522;
													assign node10522 = (inp[12]) ? node10526 : node10523;
														assign node10523 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node10526 = (inp[4]) ? node10528 : 4'b1101;
															assign node10528 = (inp[15]) ? node10530 : 4'b1111;
																assign node10530 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node10533 = (inp[13]) ? node10537 : node10534;
														assign node10534 = (inp[12]) ? 4'b1001 : 4'b1010;
														assign node10537 = (inp[15]) ? node10539 : 4'b1110;
															assign node10539 = (inp[12]) ? 4'b1100 : node10540;
																assign node10540 = (inp[4]) ? 4'b1111 : 4'b1100;
												assign node10544 = (inp[7]) ? node10558 : node10545;
													assign node10545 = (inp[15]) ? node10551 : node10546;
														assign node10546 = (inp[4]) ? 4'b1000 : node10547;
															assign node10547 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node10551 = (inp[13]) ? 4'b1111 : node10552;
															assign node10552 = (inp[12]) ? node10554 : 4'b1100;
																assign node10554 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node10558 = (inp[13]) ? node10566 : node10559;
														assign node10559 = (inp[15]) ? node10563 : node10560;
															assign node10560 = (inp[4]) ? 4'b1101 : 4'b1111;
															assign node10563 = (inp[12]) ? 4'b1110 : 4'b1111;
														assign node10566 = (inp[12]) ? node10572 : node10567;
															assign node10567 = (inp[4]) ? 4'b1110 : node10568;
																assign node10568 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node10572 = (inp[4]) ? 4'b1100 : 4'b1110;
										assign node10575 = (inp[2]) ? node10623 : node10576;
											assign node10576 = (inp[15]) ? node10602 : node10577;
												assign node10577 = (inp[7]) ? node10587 : node10578;
													assign node10578 = (inp[8]) ? node10582 : node10579;
														assign node10579 = (inp[4]) ? 4'b1001 : 4'b1110;
														assign node10582 = (inp[4]) ? node10584 : 4'b1000;
															assign node10584 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node10587 = (inp[8]) ? node10595 : node10588;
														assign node10588 = (inp[12]) ? node10590 : 4'b1110;
															assign node10590 = (inp[4]) ? node10592 : 4'b1000;
																assign node10592 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node10595 = (inp[4]) ? node10599 : node10596;
															assign node10596 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node10599 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node10602 = (inp[4]) ? node10614 : node10603;
													assign node10603 = (inp[12]) ? node10605 : 4'b1001;
														assign node10605 = (inp[7]) ? node10607 : 4'b1100;
															assign node10607 = (inp[8]) ? node10611 : node10608;
																assign node10608 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node10611 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node10614 = (inp[12]) ? node10616 : 4'b1110;
														assign node10616 = (inp[7]) ? node10618 : 4'b1101;
															assign node10618 = (inp[8]) ? 4'b1100 : node10619;
																assign node10619 = (inp[13]) ? 4'b1100 : 4'b1001;
											assign node10623 = (inp[7]) ? node10653 : node10624;
												assign node10624 = (inp[12]) ? node10640 : node10625;
													assign node10625 = (inp[15]) ? node10633 : node10626;
														assign node10626 = (inp[8]) ? node10630 : node10627;
															assign node10627 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node10630 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node10633 = (inp[4]) ? node10637 : node10634;
															assign node10634 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node10637 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node10640 = (inp[8]) ? node10648 : node10641;
														assign node10641 = (inp[13]) ? node10645 : node10642;
															assign node10642 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node10645 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node10648 = (inp[4]) ? 4'b1000 : node10649;
															assign node10649 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node10653 = (inp[4]) ? node10663 : node10654;
													assign node10654 = (inp[12]) ? node10660 : node10655;
														assign node10655 = (inp[13]) ? node10657 : 4'b1001;
															assign node10657 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node10660 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node10663 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node10666 = (inp[7]) ? node10786 : node10667;
										assign node10667 = (inp[12]) ? node10735 : node10668;
											assign node10668 = (inp[15]) ? node10700 : node10669;
												assign node10669 = (inp[8]) ? node10687 : node10670;
													assign node10670 = (inp[13]) ? node10676 : node10671;
														assign node10671 = (inp[4]) ? 4'b1000 : node10672;
															assign node10672 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node10676 = (inp[4]) ? node10682 : node10677;
															assign node10677 = (inp[2]) ? 4'b1001 : node10678;
																assign node10678 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node10682 = (inp[1]) ? node10684 : 4'b1100;
																assign node10684 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node10687 = (inp[4]) ? node10697 : node10688;
														assign node10688 = (inp[2]) ? node10694 : node10689;
															assign node10689 = (inp[1]) ? node10691 : 4'b1101;
																assign node10691 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node10694 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node10697 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node10700 = (inp[8]) ? node10718 : node10701;
													assign node10701 = (inp[4]) ? node10711 : node10702;
														assign node10702 = (inp[13]) ? 4'b1111 : node10703;
															assign node10703 = (inp[1]) ? node10707 : node10704;
																assign node10704 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node10707 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node10711 = (inp[2]) ? 4'b1001 : node10712;
															assign node10712 = (inp[1]) ? 4'b1101 : node10713;
																assign node10713 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node10718 = (inp[4]) ? node10728 : node10719;
														assign node10719 = (inp[13]) ? 4'b1000 : node10720;
															assign node10720 = (inp[1]) ? node10724 : node10721;
																assign node10721 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node10724 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node10728 = (inp[2]) ? node10732 : node10729;
															assign node10729 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node10732 = (inp[1]) ? 4'b1010 : 4'b1111;
											assign node10735 = (inp[15]) ? node10761 : node10736;
												assign node10736 = (inp[4]) ? node10756 : node10737;
													assign node10737 = (inp[2]) ? node10749 : node10738;
														assign node10738 = (inp[13]) ? node10746 : node10739;
															assign node10739 = (inp[1]) ? node10743 : node10740;
																assign node10740 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node10743 = (inp[8]) ? 4'b1110 : 4'b1011;
															assign node10746 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node10749 = (inp[8]) ? node10753 : node10750;
															assign node10750 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node10753 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node10756 = (inp[1]) ? 4'b1101 : node10757;
														assign node10757 = (inp[8]) ? 4'b1000 : 4'b1110;
												assign node10761 = (inp[4]) ? node10777 : node10762;
													assign node10762 = (inp[8]) ? 4'b1011 : node10763;
														assign node10763 = (inp[1]) ? node10769 : node10764;
															assign node10764 = (inp[2]) ? node10766 : 4'b1000;
																assign node10766 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node10769 = (inp[13]) ? node10773 : node10770;
																assign node10770 = (inp[2]) ? 4'b1000 : 4'b1101;
																assign node10773 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node10777 = (inp[8]) ? node10781 : node10778;
														assign node10778 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node10781 = (inp[13]) ? 4'b1000 : node10782;
															assign node10782 = (inp[2]) ? 4'b1000 : 4'b1100;
										assign node10786 = (inp[12]) ? node10840 : node10787;
											assign node10787 = (inp[4]) ? node10811 : node10788;
												assign node10788 = (inp[8]) ? node10800 : node10789;
													assign node10789 = (inp[15]) ? node10797 : node10790;
														assign node10790 = (inp[2]) ? 4'b1011 : node10791;
															assign node10791 = (inp[13]) ? node10793 : 4'b1110;
																assign node10793 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node10797 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node10800 = (inp[2]) ? node10802 : 4'b1001;
														assign node10802 = (inp[13]) ? node10808 : node10803;
															assign node10803 = (inp[1]) ? 4'b1001 : node10804;
																assign node10804 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node10808 = (inp[15]) ? 4'b1101 : 4'b1000;
												assign node10811 = (inp[15]) ? node10823 : node10812;
													assign node10812 = (inp[8]) ? node10820 : node10813;
														assign node10813 = (inp[1]) ? node10815 : 4'b1011;
															assign node10815 = (inp[13]) ? 4'b1011 : node10816;
																assign node10816 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node10820 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node10823 = (inp[13]) ? node10833 : node10824;
														assign node10824 = (inp[1]) ? node10828 : node10825;
															assign node10825 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node10828 = (inp[2]) ? node10830 : 4'b1010;
																assign node10830 = (inp[8]) ? 4'b1010 : 4'b1110;
														assign node10833 = (inp[1]) ? node10837 : node10834;
															assign node10834 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node10837 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node10840 = (inp[4]) ? node10872 : node10841;
												assign node10841 = (inp[2]) ? node10853 : node10842;
													assign node10842 = (inp[15]) ? node10844 : 4'b1011;
														assign node10844 = (inp[13]) ? node10850 : node10845;
															assign node10845 = (inp[1]) ? node10847 : 4'b1111;
																assign node10847 = (inp[8]) ? 4'b1111 : 4'b1011;
															assign node10850 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node10853 = (inp[1]) ? node10863 : node10854;
														assign node10854 = (inp[15]) ? node10860 : node10855;
															assign node10855 = (inp[8]) ? 4'b1110 : node10856;
																assign node10856 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node10860 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node10863 = (inp[15]) ? node10867 : node10864;
															assign node10864 = (inp[8]) ? 4'b1011 : 4'b1001;
															assign node10867 = (inp[13]) ? 4'b1011 : node10868;
																assign node10868 = (inp[8]) ? 4'b1010 : 4'b1110;
												assign node10872 = (inp[8]) ? node10884 : node10873;
													assign node10873 = (inp[2]) ? node10877 : node10874;
														assign node10874 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node10877 = (inp[13]) ? node10881 : node10878;
															assign node10878 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node10881 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node10884 = (inp[1]) ? node10894 : node10885;
														assign node10885 = (inp[2]) ? node10887 : 4'b1000;
															assign node10887 = (inp[15]) ? node10891 : node10888;
																assign node10888 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node10891 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node10894 = (inp[2]) ? node10898 : node10895;
															assign node10895 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node10898 = (inp[15]) ? node10900 : 4'b1001;
																assign node10900 = (inp[13]) ? 4'b1001 : 4'b1000;
								assign node10903 = (inp[8]) ? node11135 : node10904;
									assign node10904 = (inp[1]) ? node11024 : node10905;
										assign node10905 = (inp[4]) ? node10967 : node10906;
											assign node10906 = (inp[2]) ? node10936 : node10907;
												assign node10907 = (inp[15]) ? node10925 : node10908;
													assign node10908 = (inp[9]) ? node10916 : node10909;
														assign node10909 = (inp[13]) ? node10911 : 4'b1100;
															assign node10911 = (inp[12]) ? 4'b1100 : node10912;
																assign node10912 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node10916 = (inp[7]) ? node10922 : node10917;
															assign node10917 = (inp[12]) ? 4'b1011 : node10918;
																assign node10918 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node10922 = (inp[12]) ? 4'b1101 : 4'b1110;
													assign node10925 = (inp[7]) ? node10931 : node10926;
														assign node10926 = (inp[12]) ? 4'b1000 : node10927;
															assign node10927 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node10931 = (inp[12]) ? node10933 : 4'b1001;
															assign node10933 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node10936 = (inp[9]) ? node10952 : node10937;
													assign node10937 = (inp[15]) ? node10945 : node10938;
														assign node10938 = (inp[7]) ? node10942 : node10939;
															assign node10939 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node10942 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node10945 = (inp[13]) ? node10949 : node10946;
															assign node10946 = (inp[7]) ? 4'b1011 : 4'b1101;
															assign node10949 = (inp[7]) ? 4'b1101 : 4'b1110;
													assign node10952 = (inp[13]) ? node10960 : node10953;
														assign node10953 = (inp[7]) ? node10957 : node10954;
															assign node10954 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node10957 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node10960 = (inp[12]) ? node10962 : 4'b1111;
															assign node10962 = (inp[15]) ? 4'b1001 : node10963;
																assign node10963 = (inp[7]) ? 4'b1000 : 4'b1010;
											assign node10967 = (inp[9]) ? node11001 : node10968;
												assign node10968 = (inp[15]) ? node10982 : node10969;
													assign node10969 = (inp[12]) ? node10977 : node10970;
														assign node10970 = (inp[7]) ? 4'b1111 : node10971;
															assign node10971 = (inp[13]) ? node10973 : 4'b1100;
																assign node10973 = (inp[2]) ? 4'b1100 : 4'b1001;
														assign node10977 = (inp[13]) ? node10979 : 4'b1000;
															assign node10979 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node10982 = (inp[7]) ? node10990 : node10983;
														assign node10983 = (inp[12]) ? node10985 : 4'b1100;
															assign node10985 = (inp[13]) ? node10987 : 4'b1111;
																assign node10987 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node10990 = (inp[12]) ? node10998 : node10991;
															assign node10991 = (inp[13]) ? node10995 : node10992;
																assign node10992 = (inp[2]) ? 4'b1010 : 4'b1110;
																assign node10995 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node10998 = (inp[13]) ? 4'b1100 : 4'b1001;
												assign node11001 = (inp[2]) ? node11017 : node11002;
													assign node11002 = (inp[13]) ? node11010 : node11003;
														assign node11003 = (inp[15]) ? node11005 : 4'b1110;
															assign node11005 = (inp[7]) ? 4'b1100 : node11006;
																assign node11006 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node11010 = (inp[7]) ? node11012 : 4'b1000;
															assign node11012 = (inp[12]) ? 4'b1000 : node11013;
																assign node11013 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node11017 = (inp[13]) ? node11021 : node11018;
														assign node11018 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node11021 = (inp[7]) ? 4'b1110 : 4'b1101;
										assign node11024 = (inp[7]) ? node11076 : node11025;
											assign node11025 = (inp[12]) ? node11055 : node11026;
												assign node11026 = (inp[9]) ? node11040 : node11027;
													assign node11027 = (inp[4]) ? node11031 : node11028;
														assign node11028 = (inp[2]) ? 4'b1001 : 4'b1011;
														assign node11031 = (inp[2]) ? 4'b1001 : node11032;
															assign node11032 = (inp[13]) ? node11036 : node11033;
																assign node11033 = (inp[15]) ? 4'b1101 : 4'b1001;
																assign node11036 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node11040 = (inp[15]) ? node11048 : node11041;
														assign node11041 = (inp[13]) ? node11043 : 4'b1101;
															assign node11043 = (inp[2]) ? 4'b1000 : node11044;
																assign node11044 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node11048 = (inp[4]) ? 4'b1000 : node11049;
															assign node11049 = (inp[2]) ? node11051 : 4'b1111;
																assign node11051 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node11055 = (inp[15]) ? node11071 : node11056;
													assign node11056 = (inp[9]) ? node11068 : node11057;
														assign node11057 = (inp[4]) ? node11063 : node11058;
															assign node11058 = (inp[2]) ? 4'b1110 : node11059;
																assign node11059 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node11063 = (inp[2]) ? node11065 : 4'b1010;
																assign node11065 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node11068 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node11071 = (inp[4]) ? node11073 : 4'b1001;
														assign node11073 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node11076 = (inp[12]) ? node11106 : node11077;
												assign node11077 = (inp[4]) ? node11091 : node11078;
													assign node11078 = (inp[15]) ? node11084 : node11079;
														assign node11079 = (inp[2]) ? 4'b1110 : node11080;
															assign node11080 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11084 = (inp[13]) ? 4'b1001 : node11085;
															assign node11085 = (inp[2]) ? 4'b1000 : node11086;
																assign node11086 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node11091 = (inp[9]) ? node11099 : node11092;
														assign node11092 = (inp[15]) ? node11094 : 4'b1010;
															assign node11094 = (inp[2]) ? 4'b1110 : node11095;
																assign node11095 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node11099 = (inp[13]) ? node11103 : node11100;
															assign node11100 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node11103 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node11106 = (inp[15]) ? node11118 : node11107;
													assign node11107 = (inp[13]) ? 4'b1100 : node11108;
														assign node11108 = (inp[9]) ? 4'b1100 : node11109;
															assign node11109 = (inp[4]) ? node11113 : node11110;
																assign node11110 = (inp[2]) ? 4'b1000 : 4'b1101;
																assign node11113 = (inp[2]) ? 4'b1101 : 4'b1000;
													assign node11118 = (inp[4]) ? node11128 : node11119;
														assign node11119 = (inp[9]) ? node11125 : node11120;
															assign node11120 = (inp[13]) ? node11122 : 4'b1010;
																assign node11122 = (inp[2]) ? 4'b1010 : 4'b1111;
															assign node11125 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node11128 = (inp[9]) ? node11130 : 4'b1100;
															assign node11130 = (inp[2]) ? node11132 : 4'b1101;
																assign node11132 = (inp[13]) ? 4'b1001 : 4'b1101;
									assign node11135 = (inp[2]) ? node11223 : node11136;
										assign node11136 = (inp[1]) ? node11188 : node11137;
											assign node11137 = (inp[9]) ? node11163 : node11138;
												assign node11138 = (inp[12]) ? node11148 : node11139;
													assign node11139 = (inp[4]) ? node11141 : 4'b1101;
														assign node11141 = (inp[15]) ? node11145 : node11142;
															assign node11142 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node11145 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node11148 = (inp[4]) ? node11156 : node11149;
														assign node11149 = (inp[15]) ? node11153 : node11150;
															assign node11150 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node11153 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node11156 = (inp[7]) ? node11158 : 4'b1000;
															assign node11158 = (inp[15]) ? node11160 : 4'b1001;
																assign node11160 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node11163 = (inp[15]) ? node11173 : node11164;
													assign node11164 = (inp[7]) ? node11166 : 4'b1100;
														assign node11166 = (inp[4]) ? node11170 : node11167;
															assign node11167 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node11170 = (inp[12]) ? 4'b1001 : 4'b1010;
													assign node11173 = (inp[4]) ? node11179 : node11174;
														assign node11174 = (inp[13]) ? node11176 : 4'b1011;
															assign node11176 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node11179 = (inp[12]) ? node11185 : node11180;
															assign node11180 = (inp[13]) ? node11182 : 4'b1011;
																assign node11182 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node11185 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node11188 = (inp[15]) ? node11208 : node11189;
												assign node11189 = (inp[7]) ? node11199 : node11190;
													assign node11190 = (inp[9]) ? 4'b1001 : node11191;
														assign node11191 = (inp[13]) ? node11195 : node11192;
															assign node11192 = (inp[12]) ? 4'b1110 : 4'b1001;
															assign node11195 = (inp[12]) ? 4'b1001 : 4'b1010;
													assign node11199 = (inp[12]) ? node11203 : node11200;
														assign node11200 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node11203 = (inp[4]) ? node11205 : 4'b1110;
															assign node11205 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node11208 = (inp[4]) ? node11216 : node11209;
													assign node11209 = (inp[12]) ? 4'b1110 : node11210;
														assign node11210 = (inp[7]) ? node11212 : 4'b1101;
															assign node11212 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node11216 = (inp[12]) ? 4'b1101 : node11217;
														assign node11217 = (inp[13]) ? 4'b1111 : node11218;
															assign node11218 = (inp[7]) ? 4'b1111 : 4'b1110;
										assign node11223 = (inp[1]) ? node11253 : node11224;
											assign node11224 = (inp[12]) ? node11240 : node11225;
												assign node11225 = (inp[4]) ? node11235 : node11226;
													assign node11226 = (inp[7]) ? node11230 : node11227;
														assign node11227 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node11230 = (inp[15]) ? node11232 : 4'b1100;
															assign node11232 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node11235 = (inp[7]) ? 4'b1110 : node11236;
														assign node11236 = (inp[15]) ? 4'b1111 : 4'b1011;
												assign node11240 = (inp[4]) ? node11246 : node11241;
													assign node11241 = (inp[15]) ? 4'b1111 : node11242;
														assign node11242 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node11246 = (inp[13]) ? 4'b1101 : node11247;
														assign node11247 = (inp[15]) ? 4'b1101 : node11248;
															assign node11248 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node11253 = (inp[15]) ? node11271 : node11254;
												assign node11254 = (inp[7]) ? node11262 : node11255;
													assign node11255 = (inp[13]) ? 4'b1011 : node11256;
														assign node11256 = (inp[12]) ? 4'b1100 : node11257;
															assign node11257 = (inp[4]) ? 4'b1111 : 4'b1101;
													assign node11262 = (inp[12]) ? node11266 : node11263;
														assign node11263 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node11266 = (inp[13]) ? node11268 : 4'b1010;
															assign node11268 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node11271 = (inp[12]) ? node11279 : node11272;
													assign node11272 = (inp[4]) ? node11274 : 4'b1000;
														assign node11274 = (inp[7]) ? 4'b1011 : node11275;
															assign node11275 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node11279 = (inp[4]) ? 4'b1001 : 4'b1011;
							assign node11282 = (inp[8]) ? node11754 : node11283;
								assign node11283 = (inp[2]) ? node11539 : node11284;
									assign node11284 = (inp[11]) ? node11406 : node11285;
										assign node11285 = (inp[13]) ? node11357 : node11286;
											assign node11286 = (inp[1]) ? node11326 : node11287;
												assign node11287 = (inp[7]) ? node11303 : node11288;
													assign node11288 = (inp[12]) ? node11294 : node11289;
														assign node11289 = (inp[4]) ? 4'b1001 : node11290;
															assign node11290 = (inp[9]) ? 4'b1110 : 4'b1101;
														assign node11294 = (inp[4]) ? node11298 : node11295;
															assign node11295 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11298 = (inp[15]) ? node11300 : 4'b1111;
																assign node11300 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node11303 = (inp[12]) ? node11317 : node11304;
														assign node11304 = (inp[15]) ? node11312 : node11305;
															assign node11305 = (inp[9]) ? node11309 : node11306;
																assign node11306 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node11309 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node11312 = (inp[4]) ? 4'b1110 : node11313;
																assign node11313 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node11317 = (inp[4]) ? node11323 : node11318;
															assign node11318 = (inp[15]) ? node11320 : 4'b1001;
																assign node11320 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11323 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node11326 = (inp[12]) ? node11340 : node11327;
													assign node11327 = (inp[15]) ? node11333 : node11328;
														assign node11328 = (inp[7]) ? 4'b1011 : node11329;
															assign node11329 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node11333 = (inp[9]) ? node11335 : 4'b1101;
															assign node11335 = (inp[7]) ? node11337 : 4'b1011;
																assign node11337 = (inp[4]) ? 4'b1011 : 4'b1100;
													assign node11340 = (inp[9]) ? node11352 : node11341;
														assign node11341 = (inp[4]) ? node11349 : node11342;
															assign node11342 = (inp[15]) ? node11346 : node11343;
																assign node11343 = (inp[7]) ? 4'b1100 : 4'b1011;
																assign node11346 = (inp[7]) ? 4'b1011 : 4'b1101;
															assign node11349 = (inp[15]) ? 4'b1010 : 4'b1111;
														assign node11352 = (inp[4]) ? node11354 : 4'b1010;
															assign node11354 = (inp[15]) ? 4'b1011 : 4'b1000;
											assign node11357 = (inp[1]) ? node11383 : node11358;
												assign node11358 = (inp[15]) ? node11372 : node11359;
													assign node11359 = (inp[7]) ? node11367 : node11360;
														assign node11360 = (inp[12]) ? node11364 : node11361;
															assign node11361 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node11364 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11367 = (inp[12]) ? 4'b1001 : node11368;
															assign node11368 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node11372 = (inp[7]) ? node11376 : node11373;
														assign node11373 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node11376 = (inp[4]) ? node11380 : node11377;
															assign node11377 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node11380 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node11383 = (inp[9]) ? node11391 : node11384;
													assign node11384 = (inp[12]) ? node11388 : node11385;
														assign node11385 = (inp[7]) ? 4'b1111 : 4'b1100;
														assign node11388 = (inp[4]) ? 4'b1010 : 4'b1001;
													assign node11391 = (inp[7]) ? node11399 : node11392;
														assign node11392 = (inp[12]) ? 4'b1110 : node11393;
															assign node11393 = (inp[4]) ? 4'b1001 : node11394;
																assign node11394 = (inp[15]) ? 4'b1110 : 4'b1101;
														assign node11399 = (inp[15]) ? node11403 : node11400;
															assign node11400 = (inp[12]) ? 4'b1000 : 4'b1110;
															assign node11403 = (inp[12]) ? 4'b1100 : 4'b1000;
										assign node11406 = (inp[4]) ? node11482 : node11407;
											assign node11407 = (inp[13]) ? node11441 : node11408;
												assign node11408 = (inp[9]) ? node11432 : node11409;
													assign node11409 = (inp[1]) ? node11419 : node11410;
														assign node11410 = (inp[12]) ? node11416 : node11411;
															assign node11411 = (inp[7]) ? node11413 : 4'b1111;
																assign node11413 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node11416 = (inp[15]) ? 4'b1111 : 4'b1001;
														assign node11419 = (inp[7]) ? node11425 : node11420;
															assign node11420 = (inp[12]) ? 4'b1010 : node11421;
																assign node11421 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node11425 = (inp[15]) ? node11429 : node11426;
																assign node11426 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node11429 = (inp[12]) ? 4'b1011 : 4'b1101;
													assign node11432 = (inp[12]) ? node11438 : node11433;
														assign node11433 = (inp[7]) ? 4'b1100 : node11434;
															assign node11434 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node11438 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node11441 = (inp[1]) ? node11461 : node11442;
													assign node11442 = (inp[12]) ? node11458 : node11443;
														assign node11443 = (inp[9]) ? node11451 : node11444;
															assign node11444 = (inp[7]) ? node11448 : node11445;
																assign node11445 = (inp[15]) ? 4'b1010 : 4'b1001;
																assign node11448 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node11451 = (inp[15]) ? node11455 : node11452;
																assign node11452 = (inp[7]) ? 4'b1011 : 4'b1000;
																assign node11455 = (inp[7]) ? 4'b1001 : 4'b1011;
														assign node11458 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node11461 = (inp[15]) ? node11467 : node11462;
														assign node11462 = (inp[12]) ? 4'b1110 : node11463;
															assign node11463 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node11467 = (inp[9]) ? node11475 : node11468;
															assign node11468 = (inp[7]) ? node11472 : node11469;
																assign node11469 = (inp[12]) ? 4'b1000 : 4'b1111;
																assign node11472 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node11475 = (inp[7]) ? node11479 : node11476;
																assign node11476 = (inp[12]) ? 4'b1001 : 4'b1110;
																assign node11479 = (inp[12]) ? 4'b1111 : 4'b1001;
											assign node11482 = (inp[9]) ? node11514 : node11483;
												assign node11483 = (inp[13]) ? node11499 : node11484;
													assign node11484 = (inp[15]) ? node11492 : node11485;
														assign node11485 = (inp[12]) ? 4'b1111 : node11486;
															assign node11486 = (inp[1]) ? node11488 : 4'b1110;
																assign node11488 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node11492 = (inp[12]) ? node11496 : node11493;
															assign node11493 = (inp[7]) ? 4'b1010 : 4'b1100;
															assign node11496 = (inp[7]) ? 4'b1000 : 4'b1010;
													assign node11499 = (inp[1]) ? node11509 : node11500;
														assign node11500 = (inp[7]) ? node11504 : node11501;
															assign node11501 = (inp[15]) ? 4'b1101 : 4'b1000;
															assign node11504 = (inp[12]) ? 4'b1000 : node11505;
																assign node11505 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node11509 = (inp[7]) ? node11511 : 4'b1100;
															assign node11511 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node11514 = (inp[13]) ? node11526 : node11515;
													assign node11515 = (inp[12]) ? node11523 : node11516;
														assign node11516 = (inp[7]) ? 4'b1010 : node11517;
															assign node11517 = (inp[15]) ? 4'b1001 : node11518;
																assign node11518 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node11523 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node11526 = (inp[15]) ? node11530 : node11527;
														assign node11527 = (inp[7]) ? 4'b1110 : 4'b1010;
														assign node11530 = (inp[7]) ? node11534 : node11531;
															assign node11531 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node11534 = (inp[12]) ? node11536 : 4'b1110;
																assign node11536 = (inp[1]) ? 4'b1100 : 4'b1000;
									assign node11539 = (inp[15]) ? node11651 : node11540;
										assign node11540 = (inp[11]) ? node11602 : node11541;
											assign node11541 = (inp[9]) ? node11577 : node11542;
												assign node11542 = (inp[12]) ? node11556 : node11543;
													assign node11543 = (inp[4]) ? node11549 : node11544;
														assign node11544 = (inp[13]) ? 4'b1001 : node11545;
															assign node11545 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node11549 = (inp[1]) ? node11553 : node11550;
															assign node11550 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node11553 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node11556 = (inp[7]) ? node11566 : node11557;
														assign node11557 = (inp[13]) ? node11561 : node11558;
															assign node11558 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node11561 = (inp[4]) ? 4'b1111 : node11562;
																assign node11562 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node11566 = (inp[1]) ? node11572 : node11567;
															assign node11567 = (inp[4]) ? node11569 : 4'b1000;
																assign node11569 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node11572 = (inp[4]) ? 4'b1101 : node11573;
																assign node11573 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node11577 = (inp[1]) ? node11587 : node11578;
													assign node11578 = (inp[4]) ? node11580 : 4'b1111;
														assign node11580 = (inp[13]) ? 4'b1101 : node11581;
															assign node11581 = (inp[7]) ? node11583 : 4'b1001;
																assign node11583 = (inp[12]) ? 4'b1001 : 4'b1010;
													assign node11587 = (inp[4]) ? node11595 : node11588;
														assign node11588 = (inp[13]) ? node11590 : 4'b1000;
															assign node11590 = (inp[12]) ? 4'b1011 : node11591;
																assign node11591 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node11595 = (inp[12]) ? node11599 : node11596;
															assign node11596 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node11599 = (inp[13]) ? 4'b1000 : 4'b1010;
											assign node11602 = (inp[9]) ? node11620 : node11603;
												assign node11603 = (inp[1]) ? node11615 : node11604;
													assign node11604 = (inp[12]) ? node11608 : node11605;
														assign node11605 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node11608 = (inp[4]) ? 4'b1101 : node11609;
															assign node11609 = (inp[7]) ? 4'b1000 : node11610;
																assign node11610 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node11615 = (inp[12]) ? node11617 : 4'b1011;
														assign node11617 = (inp[13]) ? 4'b1101 : 4'b1011;
												assign node11620 = (inp[1]) ? node11644 : node11621;
													assign node11621 = (inp[13]) ? node11633 : node11622;
														assign node11622 = (inp[4]) ? node11626 : node11623;
															assign node11623 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node11626 = (inp[7]) ? node11630 : node11627;
																assign node11627 = (inp[12]) ? 4'b1011 : 4'b1000;
																assign node11630 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node11633 = (inp[12]) ? node11639 : node11634;
															assign node11634 = (inp[7]) ? 4'b1111 : node11635;
																assign node11635 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node11639 = (inp[4]) ? 4'b1111 : node11640;
																assign node11640 = (inp[7]) ? 4'b1001 : 4'b1011;
													assign node11644 = (inp[7]) ? node11646 : 4'b1110;
														assign node11646 = (inp[4]) ? 4'b1101 : node11647;
															assign node11647 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node11651 = (inp[4]) ? node11709 : node11652;
											assign node11652 = (inp[11]) ? node11678 : node11653;
												assign node11653 = (inp[7]) ? node11665 : node11654;
													assign node11654 = (inp[12]) ? 4'b1101 : node11655;
														assign node11655 = (inp[9]) ? node11657 : 4'b1111;
															assign node11657 = (inp[1]) ? node11661 : node11658;
																assign node11658 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node11661 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node11665 = (inp[12]) ? node11671 : node11666;
														assign node11666 = (inp[13]) ? 4'b1101 : node11667;
															assign node11667 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node11671 = (inp[1]) ? node11675 : node11672;
															assign node11672 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11675 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node11678 = (inp[9]) ? node11694 : node11679;
													assign node11679 = (inp[12]) ? node11689 : node11680;
														assign node11680 = (inp[7]) ? node11686 : node11681;
															assign node11681 = (inp[1]) ? node11683 : 4'b1010;
																assign node11683 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node11686 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node11689 = (inp[7]) ? node11691 : 4'b1001;
															assign node11691 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node11694 = (inp[7]) ? node11700 : node11695;
														assign node11695 = (inp[12]) ? 4'b1001 : node11696;
															assign node11696 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node11700 = (inp[12]) ? node11706 : node11701;
															assign node11701 = (inp[13]) ? node11703 : 4'b1001;
																assign node11703 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node11706 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node11709 = (inp[9]) ? node11731 : node11710;
												assign node11710 = (inp[7]) ? node11720 : node11711;
													assign node11711 = (inp[12]) ? 4'b1011 : node11712;
														assign node11712 = (inp[11]) ? 4'b1101 : node11713;
															assign node11713 = (inp[13]) ? 4'b1100 : node11714;
																assign node11714 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node11720 = (inp[12]) ? node11728 : node11721;
														assign node11721 = (inp[11]) ? 4'b1111 : node11722;
															assign node11722 = (inp[1]) ? 4'b1011 : node11723;
																assign node11723 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node11728 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node11731 = (inp[7]) ? node11737 : node11732;
													assign node11732 = (inp[12]) ? node11734 : 4'b1000;
														assign node11734 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11737 = (inp[12]) ? node11747 : node11738;
														assign node11738 = (inp[11]) ? 4'b1110 : node11739;
															assign node11739 = (inp[13]) ? node11743 : node11740;
																assign node11740 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node11743 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node11747 = (inp[13]) ? 4'b1000 : node11748;
															assign node11748 = (inp[11]) ? 4'b1100 : node11749;
																assign node11749 = (inp[1]) ? 4'b1101 : 4'b1001;
								assign node11754 = (inp[11]) ? node11934 : node11755;
									assign node11755 = (inp[7]) ? node11853 : node11756;
										assign node11756 = (inp[9]) ? node11808 : node11757;
											assign node11757 = (inp[2]) ? node11781 : node11758;
												assign node11758 = (inp[4]) ? node11770 : node11759;
													assign node11759 = (inp[12]) ? node11767 : node11760;
														assign node11760 = (inp[1]) ? node11762 : 4'b1100;
															assign node11762 = (inp[15]) ? 4'b1100 : node11763;
																assign node11763 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node11767 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node11770 = (inp[12]) ? node11776 : node11771;
														assign node11771 = (inp[15]) ? 4'b1011 : node11772;
															assign node11772 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node11776 = (inp[13]) ? node11778 : 4'b1101;
															assign node11778 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node11781 = (inp[4]) ? node11795 : node11782;
													assign node11782 = (inp[12]) ? node11790 : node11783;
														assign node11783 = (inp[15]) ? node11787 : node11784;
															assign node11784 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node11787 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node11790 = (inp[13]) ? node11792 : 4'b1010;
															assign node11792 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node11795 = (inp[12]) ? node11797 : 4'b1110;
														assign node11797 = (inp[1]) ? node11803 : node11798;
															assign node11798 = (inp[15]) ? node11800 : 4'b1001;
																assign node11800 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node11803 = (inp[15]) ? node11805 : 4'b1100;
																assign node11805 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node11808 = (inp[4]) ? node11832 : node11809;
												assign node11809 = (inp[12]) ? node11817 : node11810;
													assign node11810 = (inp[13]) ? 4'b1001 : node11811;
														assign node11811 = (inp[15]) ? 4'b1000 : node11812;
															assign node11812 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node11817 = (inp[1]) ? node11825 : node11818;
														assign node11818 = (inp[2]) ? node11820 : 4'b1010;
															assign node11820 = (inp[15]) ? node11822 : 4'b1111;
																assign node11822 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node11825 = (inp[2]) ? node11827 : 4'b1110;
															assign node11827 = (inp[15]) ? 4'b1010 : node11828;
																assign node11828 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node11832 = (inp[12]) ? node11842 : node11833;
													assign node11833 = (inp[1]) ? node11839 : node11834;
														assign node11834 = (inp[15]) ? node11836 : 4'b1011;
															assign node11836 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node11839 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node11842 = (inp[1]) ? node11844 : 4'b1001;
														assign node11844 = (inp[13]) ? node11850 : node11845;
															assign node11845 = (inp[15]) ? 4'b1001 : node11846;
																assign node11846 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node11850 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node11853 = (inp[12]) ? node11899 : node11854;
											assign node11854 = (inp[4]) ? node11882 : node11855;
												assign node11855 = (inp[13]) ? node11867 : node11856;
													assign node11856 = (inp[15]) ? node11862 : node11857;
														assign node11857 = (inp[2]) ? 4'b1100 : node11858;
															assign node11858 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node11862 = (inp[2]) ? node11864 : 4'b1000;
															assign node11864 = (inp[1]) ? 4'b1101 : 4'b1000;
													assign node11867 = (inp[15]) ? node11877 : node11868;
														assign node11868 = (inp[9]) ? node11870 : 4'b1100;
															assign node11870 = (inp[1]) ? node11874 : node11871;
																assign node11871 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node11874 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node11877 = (inp[2]) ? node11879 : 4'b1000;
															assign node11879 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node11882 = (inp[2]) ? node11888 : node11883;
													assign node11883 = (inp[1]) ? node11885 : 4'b1010;
														assign node11885 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node11888 = (inp[1]) ? node11894 : node11889;
														assign node11889 = (inp[15]) ? 4'b1111 : node11890;
															assign node11890 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node11894 = (inp[13]) ? 4'b1010 : node11895;
															assign node11895 = (inp[15]) ? 4'b1011 : 4'b1010;
											assign node11899 = (inp[4]) ? node11913 : node11900;
												assign node11900 = (inp[13]) ? node11902 : 4'b1010;
													assign node11902 = (inp[9]) ? node11904 : 4'b1111;
														assign node11904 = (inp[15]) ? node11910 : node11905;
															assign node11905 = (inp[1]) ? 4'b1010 : node11906;
																assign node11906 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node11910 = (inp[2]) ? 4'b1010 : 4'b1111;
												assign node11913 = (inp[15]) ? node11923 : node11914;
													assign node11914 = (inp[1]) ? node11920 : node11915;
														assign node11915 = (inp[2]) ? node11917 : 4'b1001;
															assign node11917 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node11920 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node11923 = (inp[2]) ? node11927 : node11924;
														assign node11924 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node11927 = (inp[1]) ? node11931 : node11928;
															assign node11928 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node11931 = (inp[13]) ? 4'b1000 : 4'b1001;
									assign node11934 = (inp[15]) ? node12024 : node11935;
										assign node11935 = (inp[7]) ? node11971 : node11936;
											assign node11936 = (inp[13]) ? node11950 : node11937;
												assign node11937 = (inp[12]) ? node11943 : node11938;
													assign node11938 = (inp[4]) ? 4'b1010 : node11939;
														assign node11939 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node11943 = (inp[4]) ? node11945 : 4'b1010;
														assign node11945 = (inp[2]) ? 4'b1101 : node11946;
															assign node11946 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node11950 = (inp[2]) ? node11964 : node11951;
													assign node11951 = (inp[9]) ? node11959 : node11952;
														assign node11952 = (inp[1]) ? 4'b1000 : node11953;
															assign node11953 = (inp[4]) ? node11955 : 4'b1010;
																assign node11955 = (inp[12]) ? 4'b1101 : 4'b1110;
														assign node11959 = (inp[1]) ? node11961 : 4'b1110;
															assign node11961 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node11964 = (inp[12]) ? node11968 : node11965;
														assign node11965 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node11968 = (inp[9]) ? 4'b1100 : 4'b1010;
											assign node11971 = (inp[2]) ? node11999 : node11972;
												assign node11972 = (inp[1]) ? node11984 : node11973;
													assign node11973 = (inp[12]) ? node11979 : node11974;
														assign node11974 = (inp[4]) ? node11976 : 4'b1001;
															assign node11976 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node11979 = (inp[4]) ? node11981 : 4'b1010;
															assign node11981 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node11984 = (inp[9]) ? node11994 : node11985;
														assign node11985 = (inp[12]) ? node11991 : node11986;
															assign node11986 = (inp[4]) ? node11988 : 4'b1101;
																assign node11988 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node11991 = (inp[4]) ? 4'b1101 : 4'b1110;
														assign node11994 = (inp[13]) ? node11996 : 4'b1101;
															assign node11996 = (inp[12]) ? 4'b1111 : 4'b1101;
												assign node11999 = (inp[1]) ? node12009 : node12000;
													assign node12000 = (inp[12]) ? node12006 : node12001;
														assign node12001 = (inp[4]) ? 4'b1111 : node12002;
															assign node12002 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node12006 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node12009 = (inp[13]) ? node12015 : node12010;
														assign node12010 = (inp[12]) ? node12012 : 4'b1000;
															assign node12012 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node12015 = (inp[9]) ? 4'b1010 : node12016;
															assign node12016 = (inp[4]) ? node12020 : node12017;
																assign node12017 = (inp[12]) ? 4'b1010 : 4'b1000;
																assign node12020 = (inp[12]) ? 4'b1000 : 4'b1010;
										assign node12024 = (inp[12]) ? node12058 : node12025;
											assign node12025 = (inp[4]) ? node12041 : node12026;
												assign node12026 = (inp[7]) ? node12032 : node12027;
													assign node12027 = (inp[1]) ? node12029 : 4'b1100;
														assign node12029 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node12032 = (inp[1]) ? 4'b1000 : node12033;
														assign node12033 = (inp[2]) ? node12037 : node12034;
															assign node12034 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node12037 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node12041 = (inp[13]) ? node12049 : node12042;
													assign node12042 = (inp[1]) ? node12046 : node12043;
														assign node12043 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node12046 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node12049 = (inp[1]) ? node12055 : node12050;
														assign node12050 = (inp[2]) ? 4'b1111 : node12051;
															assign node12051 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node12055 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node12058 = (inp[4]) ? node12068 : node12059;
												assign node12059 = (inp[2]) ? node12065 : node12060;
													assign node12060 = (inp[1]) ? 4'b1111 : node12061;
														assign node12061 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node12065 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node12068 = (inp[9]) ? node12078 : node12069;
													assign node12069 = (inp[13]) ? node12073 : node12070;
														assign node12070 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node12073 = (inp[1]) ? 4'b1000 : node12074;
															assign node12074 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node12078 = (inp[2]) ? node12080 : 4'b1100;
														assign node12080 = (inp[1]) ? 4'b1000 : 4'b1100;
			assign node12083 = (inp[8]) ? node16211 : node12084;
				assign node12084 = (inp[14]) ? node14604 : node12085;
					assign node12085 = (inp[5]) ? node13385 : node12086;
						assign node12086 = (inp[13]) ? node12720 : node12087;
							assign node12087 = (inp[12]) ? node12397 : node12088;
								assign node12088 = (inp[15]) ? node12258 : node12089;
									assign node12089 = (inp[7]) ? node12183 : node12090;
										assign node12090 = (inp[1]) ? node12140 : node12091;
											assign node12091 = (inp[0]) ? node12115 : node12092;
												assign node12092 = (inp[10]) ? node12106 : node12093;
													assign node12093 = (inp[9]) ? node12103 : node12094;
														assign node12094 = (inp[4]) ? node12098 : node12095;
															assign node12095 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node12098 = (inp[11]) ? 4'b1000 : node12099;
																assign node12099 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12103 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node12106 = (inp[2]) ? 4'b1000 : node12107;
														assign node12107 = (inp[11]) ? node12111 : node12108;
															assign node12108 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node12111 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node12115 = (inp[10]) ? node12127 : node12116;
													assign node12116 = (inp[9]) ? node12122 : node12117;
														assign node12117 = (inp[11]) ? node12119 : 4'b1000;
															assign node12119 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node12122 = (inp[11]) ? node12124 : 4'b1001;
															assign node12124 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node12127 = (inp[9]) ? node12133 : node12128;
														assign node12128 = (inp[11]) ? 4'b1001 : node12129;
															assign node12129 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12133 = (inp[4]) ? node12137 : node12134;
															assign node12134 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node12137 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node12140 = (inp[2]) ? node12166 : node12141;
												assign node12141 = (inp[4]) ? node12149 : node12142;
													assign node12142 = (inp[11]) ? node12146 : node12143;
														assign node12143 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node12146 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node12149 = (inp[10]) ? node12155 : node12150;
														assign node12150 = (inp[11]) ? 4'b1000 : node12151;
															assign node12151 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node12155 = (inp[0]) ? node12161 : node12156;
															assign node12156 = (inp[9]) ? node12158 : 4'b1001;
																assign node12158 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node12161 = (inp[11]) ? node12163 : 4'b1000;
																assign node12163 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node12166 = (inp[9]) ? node12176 : node12167;
													assign node12167 = (inp[11]) ? node12169 : 4'b1001;
														assign node12169 = (inp[0]) ? node12173 : node12170;
															assign node12170 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node12173 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node12176 = (inp[11]) ? 4'b1001 : node12177;
														assign node12177 = (inp[4]) ? node12179 : 4'b1001;
															assign node12179 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node12183 = (inp[2]) ? node12219 : node12184;
											assign node12184 = (inp[10]) ? node12198 : node12185;
												assign node12185 = (inp[0]) ? node12193 : node12186;
													assign node12186 = (inp[11]) ? node12190 : node12187;
														assign node12187 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node12190 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12193 = (inp[11]) ? 4'b1011 : node12194;
														assign node12194 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node12198 = (inp[0]) ? node12212 : node12199;
													assign node12199 = (inp[1]) ? node12207 : node12200;
														assign node12200 = (inp[4]) ? node12202 : 4'b1010;
															assign node12202 = (inp[11]) ? node12204 : 4'b1011;
																assign node12204 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node12207 = (inp[9]) ? node12209 : 4'b1011;
															assign node12209 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12212 = (inp[1]) ? 4'b1010 : node12213;
														assign node12213 = (inp[4]) ? node12215 : 4'b1011;
															assign node12215 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node12219 = (inp[10]) ? node12237 : node12220;
												assign node12220 = (inp[0]) ? node12228 : node12221;
													assign node12221 = (inp[1]) ? 4'b1010 : node12222;
														assign node12222 = (inp[4]) ? 4'b1010 : node12223;
															assign node12223 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12228 = (inp[9]) ? node12230 : 4'b1011;
														assign node12230 = (inp[1]) ? 4'b1010 : node12231;
															assign node12231 = (inp[4]) ? 4'b1011 : node12232;
																assign node12232 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node12237 = (inp[9]) ? node12247 : node12238;
													assign node12238 = (inp[4]) ? 4'b1011 : node12239;
														assign node12239 = (inp[11]) ? node12243 : node12240;
															assign node12240 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12243 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12247 = (inp[11]) ? node12253 : node12248;
														assign node12248 = (inp[4]) ? 4'b1010 : node12249;
															assign node12249 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12253 = (inp[1]) ? node12255 : 4'b1011;
															assign node12255 = (inp[4]) ? 4'b1010 : 4'b1011;
									assign node12258 = (inp[7]) ? node12330 : node12259;
										assign node12259 = (inp[1]) ? node12301 : node12260;
											assign node12260 = (inp[9]) ? node12282 : node12261;
												assign node12261 = (inp[11]) ? node12267 : node12262;
													assign node12262 = (inp[2]) ? node12264 : 4'b1010;
														assign node12264 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12267 = (inp[2]) ? node12269 : 4'b1011;
														assign node12269 = (inp[10]) ? node12275 : node12270;
															assign node12270 = (inp[4]) ? node12272 : 4'b1011;
																assign node12272 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12275 = (inp[4]) ? node12279 : node12276;
																assign node12276 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node12279 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node12282 = (inp[11]) ? node12290 : node12283;
													assign node12283 = (inp[2]) ? node12285 : 4'b1011;
														assign node12285 = (inp[0]) ? 4'b1011 : node12286;
															assign node12286 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node12290 = (inp[2]) ? node12292 : 4'b1010;
														assign node12292 = (inp[10]) ? 4'b1010 : node12293;
															assign node12293 = (inp[4]) ? node12297 : node12294;
																assign node12294 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node12297 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node12301 = (inp[4]) ? node12311 : node12302;
												assign node12302 = (inp[10]) ? 4'b1011 : node12303;
													assign node12303 = (inp[9]) ? node12307 : node12304;
														assign node12304 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12307 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node12311 = (inp[2]) ? node12319 : node12312;
													assign node12312 = (inp[0]) ? node12314 : 4'b1111;
														assign node12314 = (inp[11]) ? 4'b1111 : node12315;
															assign node12315 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12319 = (inp[10]) ? node12325 : node12320;
														assign node12320 = (inp[9]) ? 4'b1110 : node12321;
															assign node12321 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12325 = (inp[11]) ? 4'b1110 : node12326;
															assign node12326 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node12330 = (inp[1]) ? node12364 : node12331;
											assign node12331 = (inp[4]) ? node12347 : node12332;
												assign node12332 = (inp[2]) ? node12338 : node12333;
													assign node12333 = (inp[9]) ? node12335 : 4'b1101;
														assign node12335 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node12338 = (inp[9]) ? node12340 : 4'b1100;
														assign node12340 = (inp[0]) ? node12344 : node12341;
															assign node12341 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12344 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node12347 = (inp[9]) ? node12353 : node12348;
													assign node12348 = (inp[2]) ? 4'b1000 : node12349;
														assign node12349 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node12353 = (inp[11]) ? node12359 : node12354;
														assign node12354 = (inp[0]) ? node12356 : 4'b1001;
															assign node12356 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node12359 = (inp[2]) ? 4'b1000 : node12360;
															assign node12360 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node12364 = (inp[2]) ? node12380 : node12365;
												assign node12365 = (inp[4]) ? node12373 : node12366;
													assign node12366 = (inp[10]) ? 4'b1001 : node12367;
														assign node12367 = (inp[0]) ? 4'b1000 : node12368;
															assign node12368 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12373 = (inp[0]) ? 4'b1000 : node12374;
														assign node12374 = (inp[11]) ? node12376 : 4'b1000;
															assign node12376 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node12380 = (inp[0]) ? node12388 : node12381;
													assign node12381 = (inp[4]) ? 4'b1001 : node12382;
														assign node12382 = (inp[11]) ? 4'b1001 : node12383;
															assign node12383 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node12388 = (inp[9]) ? node12390 : 4'b1000;
														assign node12390 = (inp[11]) ? node12394 : node12391;
															assign node12391 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node12394 = (inp[4]) ? 4'b1001 : 4'b1000;
								assign node12397 = (inp[15]) ? node12571 : node12398;
									assign node12398 = (inp[7]) ? node12492 : node12399;
										assign node12399 = (inp[10]) ? node12449 : node12400;
											assign node12400 = (inp[11]) ? node12422 : node12401;
												assign node12401 = (inp[4]) ? node12417 : node12402;
													assign node12402 = (inp[1]) ? node12414 : node12403;
														assign node12403 = (inp[9]) ? node12409 : node12404;
															assign node12404 = (inp[2]) ? node12406 : 4'b1000;
																assign node12406 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node12409 = (inp[2]) ? node12411 : 4'b1001;
																assign node12411 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node12414 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node12417 = (inp[1]) ? node12419 : 4'b1101;
														assign node12419 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node12422 = (inp[0]) ? node12432 : node12423;
													assign node12423 = (inp[4]) ? node12429 : node12424;
														assign node12424 = (inp[1]) ? node12426 : 4'b1000;
															assign node12426 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node12429 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node12432 = (inp[2]) ? node12442 : node12433;
														assign node12433 = (inp[9]) ? node12439 : node12434;
															assign node12434 = (inp[4]) ? node12436 : 4'b1100;
																assign node12436 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node12439 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node12442 = (inp[1]) ? 4'b1101 : node12443;
															assign node12443 = (inp[4]) ? 4'b1101 : node12444;
																assign node12444 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node12449 = (inp[1]) ? node12463 : node12450;
												assign node12450 = (inp[4]) ? node12454 : node12451;
													assign node12451 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node12454 = (inp[0]) ? node12456 : 4'b1100;
														assign node12456 = (inp[9]) ? node12460 : node12457;
															assign node12457 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node12460 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node12463 = (inp[4]) ? node12481 : node12464;
													assign node12464 = (inp[2]) ? node12470 : node12465;
														assign node12465 = (inp[11]) ? 4'b1101 : node12466;
															assign node12466 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node12470 = (inp[9]) ? node12476 : node12471;
															assign node12471 = (inp[0]) ? node12473 : 4'b1100;
																assign node12473 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node12476 = (inp[11]) ? node12478 : 4'b1101;
																assign node12478 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node12481 = (inp[9]) ? node12483 : 4'b1000;
														assign node12483 = (inp[11]) ? node12487 : node12484;
															assign node12484 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node12487 = (inp[0]) ? node12489 : 4'b1001;
																assign node12489 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node12492 = (inp[4]) ? node12526 : node12493;
											assign node12493 = (inp[1]) ? node12509 : node12494;
												assign node12494 = (inp[2]) ? node12502 : node12495;
													assign node12495 = (inp[11]) ? 4'b1011 : node12496;
														assign node12496 = (inp[9]) ? node12498 : 4'b1011;
															assign node12498 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12502 = (inp[9]) ? node12506 : node12503;
														assign node12503 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12506 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node12509 = (inp[9]) ? node12515 : node12510;
													assign node12510 = (inp[11]) ? 4'b1111 : node12511;
														assign node12511 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node12515 = (inp[11]) ? node12521 : node12516;
														assign node12516 = (inp[0]) ? 4'b1111 : node12517;
															assign node12517 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node12521 = (inp[2]) ? 4'b1110 : node12522;
															assign node12522 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node12526 = (inp[1]) ? node12560 : node12527;
												assign node12527 = (inp[0]) ? node12545 : node12528;
													assign node12528 = (inp[10]) ? node12540 : node12529;
														assign node12529 = (inp[2]) ? node12535 : node12530;
															assign node12530 = (inp[11]) ? node12532 : 4'b1110;
																assign node12532 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12535 = (inp[9]) ? 4'b1111 : node12536;
																assign node12536 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12540 = (inp[11]) ? node12542 : 4'b1110;
															assign node12542 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12545 = (inp[2]) ? node12553 : node12546;
														assign node12546 = (inp[9]) ? node12550 : node12547;
															assign node12547 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node12550 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12553 = (inp[9]) ? node12557 : node12554;
															assign node12554 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12557 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12560 = (inp[9]) ? node12566 : node12561;
													assign node12561 = (inp[11]) ? node12563 : 4'b1010;
														assign node12563 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12566 = (inp[11]) ? node12568 : 4'b1011;
														assign node12568 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node12571 = (inp[7]) ? node12649 : node12572;
										assign node12572 = (inp[4]) ? node12604 : node12573;
											assign node12573 = (inp[1]) ? node12591 : node12574;
												assign node12574 = (inp[9]) ? node12586 : node12575;
													assign node12575 = (inp[11]) ? node12581 : node12576;
														assign node12576 = (inp[2]) ? node12578 : 4'b1010;
															assign node12578 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12581 = (inp[2]) ? node12583 : 4'b1011;
															assign node12583 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12586 = (inp[11]) ? 4'b1010 : node12587;
														assign node12587 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node12591 = (inp[11]) ? node12597 : node12592;
													assign node12592 = (inp[0]) ? node12594 : 4'b1110;
														assign node12594 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12597 = (inp[9]) ? node12599 : 4'b1111;
														assign node12599 = (inp[0]) ? 4'b1110 : node12600;
															assign node12600 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node12604 = (inp[9]) ? node12626 : node12605;
												assign node12605 = (inp[11]) ? node12619 : node12606;
													assign node12606 = (inp[10]) ? node12612 : node12607;
														assign node12607 = (inp[0]) ? 4'b1010 : node12608;
															assign node12608 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12612 = (inp[0]) ? 4'b1011 : node12613;
															assign node12613 = (inp[2]) ? node12615 : 4'b1010;
																assign node12615 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node12619 = (inp[0]) ? 4'b1011 : node12620;
														assign node12620 = (inp[2]) ? node12622 : 4'b1011;
															assign node12622 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node12626 = (inp[11]) ? node12638 : node12627;
													assign node12627 = (inp[1]) ? node12633 : node12628;
														assign node12628 = (inp[2]) ? 4'b1011 : node12629;
															assign node12629 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node12633 = (inp[2]) ? node12635 : 4'b1011;
															assign node12635 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12638 = (inp[10]) ? 4'b1010 : node12639;
														assign node12639 = (inp[1]) ? node12643 : node12640;
															assign node12640 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12643 = (inp[0]) ? 4'b1010 : node12644;
																assign node12644 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node12649 = (inp[1]) ? node12687 : node12650;
											assign node12650 = (inp[4]) ? node12664 : node12651;
												assign node12651 = (inp[9]) ? node12659 : node12652;
													assign node12652 = (inp[0]) ? node12654 : 4'b1001;
														assign node12654 = (inp[2]) ? node12656 : 4'b1000;
															assign node12656 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12659 = (inp[11]) ? node12661 : 4'b1000;
														assign node12661 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node12664 = (inp[2]) ? node12672 : node12665;
													assign node12665 = (inp[11]) ? node12669 : node12666;
														assign node12666 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node12669 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node12672 = (inp[10]) ? node12684 : node12673;
														assign node12673 = (inp[0]) ? node12679 : node12674;
															assign node12674 = (inp[9]) ? node12676 : 4'b1100;
																assign node12676 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12679 = (inp[9]) ? node12681 : 4'b1101;
																assign node12681 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12684 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node12687 = (inp[9]) ? node12703 : node12688;
												assign node12688 = (inp[0]) ? node12700 : node12689;
													assign node12689 = (inp[11]) ? node12691 : 4'b1000;
														assign node12691 = (inp[10]) ? node12693 : 4'b1001;
															assign node12693 = (inp[2]) ? node12697 : node12694;
																assign node12694 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node12697 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node12700 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node12703 = (inp[11]) ? node12711 : node12704;
													assign node12704 = (inp[0]) ? 4'b1000 : node12705;
														assign node12705 = (inp[2]) ? 4'b1001 : node12706;
															assign node12706 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node12711 = (inp[0]) ? 4'b1001 : node12712;
														assign node12712 = (inp[2]) ? node12716 : node12713;
															assign node12713 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node12716 = (inp[4]) ? 4'b1000 : 4'b1001;
							assign node12720 = (inp[12]) ? node13052 : node12721;
								assign node12721 = (inp[15]) ? node12873 : node12722;
									assign node12722 = (inp[7]) ? node12790 : node12723;
										assign node12723 = (inp[10]) ? node12755 : node12724;
											assign node12724 = (inp[11]) ? node12746 : node12725;
												assign node12725 = (inp[9]) ? node12733 : node12726;
													assign node12726 = (inp[4]) ? 4'b1100 : node12727;
														assign node12727 = (inp[0]) ? node12729 : 4'b1100;
															assign node12729 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node12733 = (inp[2]) ? node12735 : 4'b1101;
														assign node12735 = (inp[1]) ? node12741 : node12736;
															assign node12736 = (inp[0]) ? 4'b1101 : node12737;
																assign node12737 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node12741 = (inp[0]) ? node12743 : 4'b1101;
																assign node12743 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node12746 = (inp[9]) ? node12752 : node12747;
													assign node12747 = (inp[2]) ? node12749 : 4'b1101;
														assign node12749 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node12752 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node12755 = (inp[11]) ? node12767 : node12756;
												assign node12756 = (inp[9]) ? node12758 : 4'b1100;
													assign node12758 = (inp[2]) ? node12760 : 4'b1101;
														assign node12760 = (inp[4]) ? node12764 : node12761;
															assign node12761 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node12764 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node12767 = (inp[9]) ? node12777 : node12768;
													assign node12768 = (inp[2]) ? node12770 : 4'b1101;
														assign node12770 = (inp[4]) ? node12774 : node12771;
															assign node12771 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node12774 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node12777 = (inp[2]) ? node12779 : 4'b1100;
														assign node12779 = (inp[1]) ? node12785 : node12780;
															assign node12780 = (inp[0]) ? 4'b1101 : node12781;
																assign node12781 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node12785 = (inp[0]) ? 4'b1100 : node12786;
																assign node12786 = (inp[4]) ? 4'b1101 : 4'b1100;
										assign node12790 = (inp[10]) ? node12832 : node12791;
											assign node12791 = (inp[2]) ? node12807 : node12792;
												assign node12792 = (inp[0]) ? node12800 : node12793;
													assign node12793 = (inp[1]) ? 4'b1110 : node12794;
														assign node12794 = (inp[11]) ? 4'b1110 : node12795;
															assign node12795 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12800 = (inp[9]) ? node12804 : node12801;
														assign node12801 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12804 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12807 = (inp[11]) ? node12819 : node12808;
													assign node12808 = (inp[1]) ? node12810 : 4'b1110;
														assign node12810 = (inp[4]) ? 4'b1111 : node12811;
															assign node12811 = (inp[9]) ? node12815 : node12812;
																assign node12812 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node12815 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node12819 = (inp[1]) ? node12821 : 4'b1111;
														assign node12821 = (inp[9]) ? node12827 : node12822;
															assign node12822 = (inp[4]) ? node12824 : 4'b1111;
																assign node12824 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12827 = (inp[0]) ? 4'b1110 : node12828;
																assign node12828 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node12832 = (inp[4]) ? node12856 : node12833;
												assign node12833 = (inp[2]) ? node12847 : node12834;
													assign node12834 = (inp[1]) ? node12842 : node12835;
														assign node12835 = (inp[9]) ? node12839 : node12836;
															assign node12836 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12839 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12842 = (inp[11]) ? node12844 : 4'b1111;
															assign node12844 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12847 = (inp[11]) ? node12849 : 4'b1110;
														assign node12849 = (inp[1]) ? node12851 : 4'b1111;
															assign node12851 = (inp[9]) ? node12853 : 4'b1110;
																assign node12853 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node12856 = (inp[9]) ? node12864 : node12857;
													assign node12857 = (inp[0]) ? 4'b1110 : node12858;
														assign node12858 = (inp[2]) ? 4'b1111 : node12859;
															assign node12859 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12864 = (inp[11]) ? node12868 : node12865;
														assign node12865 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node12868 = (inp[0]) ? 4'b1110 : node12869;
															assign node12869 = (inp[1]) ? 4'b1111 : 4'b1110;
									assign node12873 = (inp[7]) ? node12969 : node12874;
										assign node12874 = (inp[1]) ? node12920 : node12875;
											assign node12875 = (inp[2]) ? node12889 : node12876;
												assign node12876 = (inp[0]) ? node12884 : node12877;
													assign node12877 = (inp[9]) ? node12881 : node12878;
														assign node12878 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12881 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12884 = (inp[10]) ? 4'b1111 : node12885;
														assign node12885 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node12889 = (inp[9]) ? node12907 : node12890;
													assign node12890 = (inp[0]) ? node12900 : node12891;
														assign node12891 = (inp[10]) ? node12895 : node12892;
															assign node12892 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node12895 = (inp[11]) ? 4'b1111 : node12896;
																assign node12896 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node12900 = (inp[11]) ? node12904 : node12901;
															assign node12901 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node12904 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node12907 = (inp[4]) ? node12913 : node12908;
														assign node12908 = (inp[11]) ? 4'b1110 : node12909;
															assign node12909 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node12913 = (inp[11]) ? node12917 : node12914;
															assign node12914 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12917 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node12920 = (inp[4]) ? node12948 : node12921;
												assign node12921 = (inp[10]) ? node12939 : node12922;
													assign node12922 = (inp[2]) ? node12934 : node12923;
														assign node12923 = (inp[9]) ? node12929 : node12924;
															assign node12924 = (inp[11]) ? 4'b1111 : node12925;
																assign node12925 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12929 = (inp[0]) ? node12931 : 4'b1110;
																assign node12931 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12934 = (inp[9]) ? 4'b1111 : node12935;
															assign node12935 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12939 = (inp[0]) ? node12941 : 4'b1110;
														assign node12941 = (inp[9]) ? node12945 : node12942;
															assign node12942 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12945 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12948 = (inp[9]) ? node12960 : node12949;
													assign node12949 = (inp[11]) ? node12955 : node12950;
														assign node12950 = (inp[0]) ? 4'b1010 : node12951;
															assign node12951 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12955 = (inp[0]) ? 4'b1011 : node12956;
															assign node12956 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node12960 = (inp[11]) ? node12964 : node12961;
														assign node12961 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node12964 = (inp[0]) ? 4'b1010 : node12965;
															assign node12965 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node12969 = (inp[4]) ? node13019 : node12970;
											assign node12970 = (inp[1]) ? node12986 : node12971;
												assign node12971 = (inp[2]) ? node12979 : node12972;
													assign node12972 = (inp[11]) ? node12974 : 4'b1001;
														assign node12974 = (inp[9]) ? node12976 : 4'b1001;
															assign node12976 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node12979 = (inp[9]) ? node12983 : node12980;
														assign node12980 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12983 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node12986 = (inp[10]) ? node12998 : node12987;
													assign node12987 = (inp[2]) ? 4'b1100 : node12988;
														assign node12988 = (inp[0]) ? 4'b1100 : node12989;
															assign node12989 = (inp[11]) ? node12993 : node12990;
																assign node12990 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node12993 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node12998 = (inp[0]) ? node13004 : node12999;
														assign node12999 = (inp[11]) ? node13001 : 4'b1101;
															assign node13001 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node13004 = (inp[11]) ? node13012 : node13005;
															assign node13005 = (inp[9]) ? node13009 : node13006;
																assign node13006 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node13009 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node13012 = (inp[2]) ? node13016 : node13013;
																assign node13013 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node13016 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node13019 = (inp[0]) ? node13029 : node13020;
												assign node13020 = (inp[9]) ? node13026 : node13021;
													assign node13021 = (inp[11]) ? node13023 : 4'b1101;
														assign node13023 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node13026 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node13029 = (inp[11]) ? node13039 : node13030;
													assign node13030 = (inp[1]) ? 4'b1100 : node13031;
														assign node13031 = (inp[9]) ? node13035 : node13032;
															assign node13032 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13035 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node13039 = (inp[9]) ? node13047 : node13040;
														assign node13040 = (inp[10]) ? 4'b1101 : node13041;
															assign node13041 = (inp[1]) ? 4'b1101 : node13042;
																assign node13042 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node13047 = (inp[1]) ? 4'b1100 : node13048;
															assign node13048 = (inp[2]) ? 4'b1101 : 4'b1100;
								assign node13052 = (inp[15]) ? node13244 : node13053;
									assign node13053 = (inp[7]) ? node13155 : node13054;
										assign node13054 = (inp[10]) ? node13116 : node13055;
											assign node13055 = (inp[2]) ? node13087 : node13056;
												assign node13056 = (inp[1]) ? node13072 : node13057;
													assign node13057 = (inp[4]) ? node13063 : node13058;
														assign node13058 = (inp[0]) ? node13060 : 4'b1100;
															assign node13060 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node13063 = (inp[11]) ? node13065 : 4'b1000;
															assign node13065 = (inp[0]) ? node13069 : node13066;
																assign node13066 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node13069 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13072 = (inp[4]) ? node13080 : node13073;
														assign node13073 = (inp[11]) ? 4'b1001 : node13074;
															assign node13074 = (inp[9]) ? node13076 : 4'b1001;
																assign node13076 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node13080 = (inp[9]) ? node13082 : 4'b1100;
															assign node13082 = (inp[0]) ? node13084 : 4'b1101;
																assign node13084 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node13087 = (inp[0]) ? node13105 : node13088;
													assign node13088 = (inp[4]) ? node13096 : node13089;
														assign node13089 = (inp[1]) ? 4'b1001 : node13090;
															assign node13090 = (inp[11]) ? node13092 : 4'b1101;
																assign node13092 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node13096 = (inp[1]) ? node13102 : node13097;
															assign node13097 = (inp[9]) ? 4'b1001 : node13098;
																assign node13098 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13102 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13105 = (inp[1]) ? node13111 : node13106;
														assign node13106 = (inp[9]) ? node13108 : 4'b1001;
															assign node13108 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13111 = (inp[4]) ? 4'b1101 : node13112;
															assign node13112 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node13116 = (inp[4]) ? node13138 : node13117;
												assign node13117 = (inp[1]) ? node13127 : node13118;
													assign node13118 = (inp[0]) ? 4'b1101 : node13119;
														assign node13119 = (inp[11]) ? node13123 : node13120;
															assign node13120 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node13123 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node13127 = (inp[9]) ? node13129 : 4'b1000;
														assign node13129 = (inp[0]) ? 4'b1001 : node13130;
															assign node13130 = (inp[2]) ? node13134 : node13131;
																assign node13131 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13134 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node13138 = (inp[1]) ? node13142 : node13139;
													assign node13139 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node13142 = (inp[2]) ? node13150 : node13143;
														assign node13143 = (inp[9]) ? node13147 : node13144;
															assign node13144 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13147 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13150 = (inp[9]) ? node13152 : 4'b1101;
															assign node13152 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node13155 = (inp[4]) ? node13209 : node13156;
											assign node13156 = (inp[1]) ? node13176 : node13157;
												assign node13157 = (inp[10]) ? node13165 : node13158;
													assign node13158 = (inp[9]) ? node13160 : 4'b1110;
														assign node13160 = (inp[11]) ? node13162 : 4'b1110;
															assign node13162 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node13165 = (inp[11]) ? node13173 : node13166;
														assign node13166 = (inp[9]) ? 4'b1110 : node13167;
															assign node13167 = (inp[0]) ? 4'b1111 : node13168;
																assign node13168 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node13173 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node13176 = (inp[2]) ? node13190 : node13177;
													assign node13177 = (inp[0]) ? node13185 : node13178;
														assign node13178 = (inp[11]) ? node13182 : node13179;
															assign node13179 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node13182 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node13185 = (inp[10]) ? node13187 : 4'b1010;
															assign node13187 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13190 = (inp[11]) ? node13204 : node13191;
														assign node13191 = (inp[10]) ? node13197 : node13192;
															assign node13192 = (inp[9]) ? node13194 : 4'b1010;
																assign node13194 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node13197 = (inp[0]) ? node13201 : node13198;
																assign node13198 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node13201 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node13204 = (inp[0]) ? node13206 : 4'b1011;
															assign node13206 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node13209 = (inp[1]) ? node13225 : node13210;
												assign node13210 = (inp[9]) ? node13218 : node13211;
													assign node13211 = (inp[11]) ? node13213 : 4'b1011;
														assign node13213 = (inp[0]) ? 4'b1010 : node13214;
															assign node13214 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node13218 = (inp[11]) ? node13220 : 4'b1010;
														assign node13220 = (inp[0]) ? 4'b1011 : node13221;
															assign node13221 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node13225 = (inp[9]) ? node13235 : node13226;
													assign node13226 = (inp[0]) ? 4'b1111 : node13227;
														assign node13227 = (inp[10]) ? node13229 : 4'b1111;
															assign node13229 = (inp[11]) ? node13231 : 4'b1110;
																assign node13231 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node13235 = (inp[0]) ? 4'b1110 : node13236;
														assign node13236 = (inp[2]) ? node13240 : node13237;
															assign node13237 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13240 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node13244 = (inp[7]) ? node13312 : node13245;
										assign node13245 = (inp[4]) ? node13287 : node13246;
											assign node13246 = (inp[1]) ? node13274 : node13247;
												assign node13247 = (inp[10]) ? node13257 : node13248;
													assign node13248 = (inp[11]) ? 4'b1111 : node13249;
														assign node13249 = (inp[2]) ? node13253 : node13250;
															assign node13250 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node13253 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node13257 = (inp[11]) ? node13269 : node13258;
														assign node13258 = (inp[9]) ? node13264 : node13259;
															assign node13259 = (inp[2]) ? node13261 : 4'b1111;
																assign node13261 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node13264 = (inp[0]) ? node13266 : 4'b1110;
																assign node13266 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node13269 = (inp[9]) ? node13271 : 4'b1110;
															assign node13271 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node13274 = (inp[10]) ? node13284 : node13275;
													assign node13275 = (inp[9]) ? node13277 : 4'b1010;
														assign node13277 = (inp[11]) ? node13279 : 4'b1010;
															assign node13279 = (inp[0]) ? node13281 : 4'b1011;
																assign node13281 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node13284 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node13287 = (inp[11]) ? node13301 : node13288;
												assign node13288 = (inp[9]) ? node13294 : node13289;
													assign node13289 = (inp[2]) ? node13291 : 4'b1111;
														assign node13291 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node13294 = (inp[1]) ? node13296 : 4'b1111;
														assign node13296 = (inp[0]) ? 4'b1110 : node13297;
															assign node13297 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node13301 = (inp[9]) ? node13309 : node13302;
													assign node13302 = (inp[10]) ? node13304 : 4'b1110;
														assign node13304 = (inp[2]) ? node13306 : 4'b1110;
															assign node13306 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node13309 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node13312 = (inp[1]) ? node13356 : node13313;
											assign node13313 = (inp[4]) ? node13337 : node13314;
												assign node13314 = (inp[10]) ? node13326 : node13315;
													assign node13315 = (inp[2]) ? node13321 : node13316;
														assign node13316 = (inp[11]) ? node13318 : 4'b1101;
															assign node13318 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node13321 = (inp[11]) ? node13323 : 4'b1100;
															assign node13323 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13326 = (inp[9]) ? 4'b1101 : node13327;
														assign node13327 = (inp[0]) ? node13329 : 4'b1100;
															assign node13329 = (inp[11]) ? node13333 : node13330;
																assign node13330 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node13333 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node13337 = (inp[9]) ? node13347 : node13338;
													assign node13338 = (inp[11]) ? node13344 : node13339;
														assign node13339 = (inp[2]) ? 4'b1000 : node13340;
															assign node13340 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node13344 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node13347 = (inp[10]) ? node13349 : 4'b1001;
														assign node13349 = (inp[2]) ? node13353 : node13350;
															assign node13350 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13353 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node13356 = (inp[11]) ? node13376 : node13357;
												assign node13357 = (inp[9]) ? node13369 : node13358;
													assign node13358 = (inp[0]) ? 4'b1100 : node13359;
														assign node13359 = (inp[10]) ? node13361 : 4'b1101;
															assign node13361 = (inp[4]) ? node13365 : node13362;
																assign node13362 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node13365 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node13369 = (inp[0]) ? 4'b1101 : node13370;
														assign node13370 = (inp[2]) ? 4'b1100 : node13371;
															assign node13371 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node13376 = (inp[9]) ? node13380 : node13377;
													assign node13377 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13380 = (inp[0]) ? 4'b1100 : node13381;
														assign node13381 = (inp[4]) ? 4'b1101 : 4'b1100;
						assign node13385 = (inp[13]) ? node13965 : node13386;
							assign node13386 = (inp[12]) ? node13656 : node13387;
								assign node13387 = (inp[15]) ? node13519 : node13388;
									assign node13388 = (inp[7]) ? node13454 : node13389;
										assign node13389 = (inp[1]) ? node13421 : node13390;
											assign node13390 = (inp[0]) ? node13416 : node13391;
												assign node13391 = (inp[2]) ? node13403 : node13392;
													assign node13392 = (inp[4]) ? node13398 : node13393;
														assign node13393 = (inp[11]) ? 4'b1101 : node13394;
															assign node13394 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node13398 = (inp[9]) ? 4'b1100 : node13399;
															assign node13399 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13403 = (inp[4]) ? 4'b1101 : node13404;
														assign node13404 = (inp[10]) ? node13410 : node13405;
															assign node13405 = (inp[9]) ? node13407 : 4'b1101;
																assign node13407 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13410 = (inp[11]) ? 4'b1101 : node13411;
																assign node13411 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node13416 = (inp[2]) ? node13418 : 4'b1101;
													assign node13418 = (inp[4]) ? 4'b1100 : 4'b1101;
											assign node13421 = (inp[9]) ? node13437 : node13422;
												assign node13422 = (inp[4]) ? node13432 : node13423;
													assign node13423 = (inp[0]) ? node13425 : 4'b1101;
														assign node13425 = (inp[2]) ? node13429 : node13426;
															assign node13426 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13429 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13432 = (inp[0]) ? node13434 : 4'b1100;
														assign node13434 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node13437 = (inp[2]) ? node13447 : node13438;
													assign node13438 = (inp[4]) ? node13440 : 4'b1100;
														assign node13440 = (inp[11]) ? node13444 : node13441;
															assign node13441 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13444 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13447 = (inp[10]) ? node13449 : 4'b1100;
														assign node13449 = (inp[4]) ? 4'b1100 : node13450;
															assign node13450 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node13454 = (inp[10]) ? node13490 : node13455;
											assign node13455 = (inp[1]) ? node13469 : node13456;
												assign node13456 = (inp[0]) ? node13464 : node13457;
													assign node13457 = (inp[9]) ? node13461 : node13458;
														assign node13458 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node13461 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node13464 = (inp[9]) ? 4'b1110 : node13465;
														assign node13465 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node13469 = (inp[9]) ? node13481 : node13470;
													assign node13470 = (inp[2]) ? 4'b1111 : node13471;
														assign node13471 = (inp[11]) ? node13477 : node13472;
															assign node13472 = (inp[0]) ? node13474 : 4'b1111;
																assign node13474 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node13477 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node13481 = (inp[11]) ? node13483 : 4'b1110;
														assign node13483 = (inp[0]) ? node13485 : 4'b1111;
															assign node13485 = (inp[4]) ? 4'b1110 : node13486;
																assign node13486 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node13490 = (inp[2]) ? node13500 : node13491;
												assign node13491 = (inp[9]) ? 4'b1110 : node13492;
													assign node13492 = (inp[11]) ? node13494 : 4'b1111;
														assign node13494 = (inp[0]) ? node13496 : 4'b1110;
															assign node13496 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node13500 = (inp[9]) ? node13510 : node13501;
													assign node13501 = (inp[11]) ? node13505 : node13502;
														assign node13502 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node13505 = (inp[4]) ? 4'b1110 : node13506;
															assign node13506 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node13510 = (inp[11]) ? node13514 : node13511;
														assign node13511 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node13514 = (inp[0]) ? node13516 : 4'b1111;
															assign node13516 = (inp[4]) ? 4'b1111 : 4'b1110;
									assign node13519 = (inp[7]) ? node13595 : node13520;
										assign node13520 = (inp[1]) ? node13552 : node13521;
											assign node13521 = (inp[10]) ? node13537 : node13522;
												assign node13522 = (inp[11]) ? node13524 : 4'b1111;
													assign node13524 = (inp[9]) ? node13530 : node13525;
														assign node13525 = (inp[2]) ? node13527 : 4'b1111;
															assign node13527 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13530 = (inp[4]) ? node13532 : 4'b1110;
															assign node13532 = (inp[2]) ? 4'b1110 : node13533;
																assign node13533 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node13537 = (inp[0]) ? node13545 : node13538;
													assign node13538 = (inp[2]) ? 4'b1111 : node13539;
														assign node13539 = (inp[11]) ? 4'b1110 : node13540;
															assign node13540 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node13545 = (inp[2]) ? 4'b1110 : node13546;
														assign node13546 = (inp[9]) ? 4'b1110 : node13547;
															assign node13547 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node13552 = (inp[4]) ? node13568 : node13553;
												assign node13553 = (inp[9]) ? node13557 : node13554;
													assign node13554 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node13557 = (inp[2]) ? 4'b1110 : node13558;
														assign node13558 = (inp[10]) ? node13560 : 4'b1111;
															assign node13560 = (inp[0]) ? node13564 : node13561;
																assign node13561 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node13564 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node13568 = (inp[2]) ? node13584 : node13569;
													assign node13569 = (inp[11]) ? node13571 : 4'b1010;
														assign node13571 = (inp[10]) ? node13579 : node13572;
															assign node13572 = (inp[9]) ? node13576 : node13573;
																assign node13573 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node13576 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node13579 = (inp[9]) ? 4'b1010 : node13580;
																assign node13580 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node13584 = (inp[0]) ? node13590 : node13585;
														assign node13585 = (inp[9]) ? node13587 : 4'b1011;
															assign node13587 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node13590 = (inp[9]) ? node13592 : 4'b1010;
															assign node13592 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node13595 = (inp[4]) ? node13627 : node13596;
											assign node13596 = (inp[1]) ? node13614 : node13597;
												assign node13597 = (inp[11]) ? node13603 : node13598;
													assign node13598 = (inp[9]) ? node13600 : 4'b1000;
														assign node13600 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node13603 = (inp[9]) ? node13609 : node13604;
														assign node13604 = (inp[2]) ? 4'b1001 : node13605;
															assign node13605 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node13609 = (inp[2]) ? 4'b1000 : node13610;
															assign node13610 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node13614 = (inp[2]) ? node13622 : node13615;
													assign node13615 = (inp[11]) ? node13619 : node13616;
														assign node13616 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node13619 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13622 = (inp[9]) ? 4'b1100 : node13623;
														assign node13623 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node13627 = (inp[0]) ? node13647 : node13628;
												assign node13628 = (inp[9]) ? node13640 : node13629;
													assign node13629 = (inp[2]) ? node13631 : 4'b1100;
														assign node13631 = (inp[10]) ? node13637 : node13632;
															assign node13632 = (inp[11]) ? 4'b1100 : node13633;
																assign node13633 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node13637 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13640 = (inp[11]) ? node13644 : node13641;
														assign node13641 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node13644 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node13647 = (inp[1]) ? 4'b1101 : node13648;
													assign node13648 = (inp[9]) ? node13652 : node13649;
														assign node13649 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13652 = (inp[11]) ? 4'b1100 : 4'b1101;
								assign node13656 = (inp[15]) ? node13790 : node13657;
									assign node13657 = (inp[7]) ? node13735 : node13658;
										assign node13658 = (inp[4]) ? node13692 : node13659;
											assign node13659 = (inp[1]) ? node13675 : node13660;
												assign node13660 = (inp[10]) ? node13670 : node13661;
													assign node13661 = (inp[11]) ? node13663 : 4'b1101;
														assign node13663 = (inp[2]) ? node13665 : 4'b1100;
															assign node13665 = (inp[0]) ? node13667 : 4'b1101;
																assign node13667 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node13670 = (inp[0]) ? 4'b1100 : node13671;
														assign node13671 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node13675 = (inp[9]) ? node13687 : node13676;
													assign node13676 = (inp[11]) ? node13682 : node13677;
														assign node13677 = (inp[2]) ? 4'b1000 : node13678;
															assign node13678 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node13682 = (inp[0]) ? 4'b1001 : node13683;
															assign node13683 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node13687 = (inp[11]) ? node13689 : 4'b1001;
														assign node13689 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node13692 = (inp[1]) ? node13716 : node13693;
												assign node13693 = (inp[10]) ? node13705 : node13694;
													assign node13694 = (inp[11]) ? 4'b1000 : node13695;
														assign node13695 = (inp[0]) ? 4'b1000 : node13696;
															assign node13696 = (inp[2]) ? node13700 : node13697;
																assign node13697 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node13700 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13705 = (inp[9]) ? node13713 : node13706;
														assign node13706 = (inp[11]) ? node13708 : 4'b1001;
															assign node13708 = (inp[2]) ? node13710 : 4'b1000;
																assign node13710 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node13713 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node13716 = (inp[11]) ? node13724 : node13717;
													assign node13717 = (inp[9]) ? node13719 : 4'b1100;
														assign node13719 = (inp[0]) ? 4'b1101 : node13720;
															assign node13720 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node13724 = (inp[10]) ? 4'b1101 : node13725;
														assign node13725 = (inp[9]) ? node13731 : node13726;
															assign node13726 = (inp[2]) ? node13728 : 4'b1101;
																assign node13728 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node13731 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node13735 = (inp[4]) ? node13763 : node13736;
											assign node13736 = (inp[1]) ? node13746 : node13737;
												assign node13737 = (inp[9]) ? 4'b1110 : node13738;
													assign node13738 = (inp[11]) ? node13740 : 4'b1110;
														assign node13740 = (inp[2]) ? 4'b1111 : node13741;
															assign node13741 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node13746 = (inp[11]) ? node13758 : node13747;
													assign node13747 = (inp[9]) ? node13753 : node13748;
														assign node13748 = (inp[10]) ? node13750 : 4'b1011;
															assign node13750 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node13753 = (inp[2]) ? node13755 : 4'b1010;
															assign node13755 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node13758 = (inp[9]) ? node13760 : 4'b1010;
														assign node13760 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node13763 = (inp[1]) ? node13773 : node13764;
												assign node13764 = (inp[11]) ? node13766 : 4'b1011;
													assign node13766 = (inp[2]) ? 4'b1010 : node13767;
														assign node13767 = (inp[0]) ? 4'b1011 : node13768;
															assign node13768 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node13773 = (inp[9]) ? node13779 : node13774;
													assign node13774 = (inp[11]) ? 4'b1110 : node13775;
														assign node13775 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node13779 = (inp[11]) ? node13785 : node13780;
														assign node13780 = (inp[0]) ? node13782 : 4'b1110;
															assign node13782 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node13785 = (inp[2]) ? 4'b1111 : node13786;
															assign node13786 = (inp[10]) ? 4'b1110 : 4'b1111;
									assign node13790 = (inp[7]) ? node13874 : node13791;
										assign node13791 = (inp[1]) ? node13831 : node13792;
											assign node13792 = (inp[9]) ? node13812 : node13793;
												assign node13793 = (inp[11]) ? node13805 : node13794;
													assign node13794 = (inp[0]) ? node13802 : node13795;
														assign node13795 = (inp[10]) ? node13797 : 4'b1110;
															assign node13797 = (inp[4]) ? node13799 : 4'b1110;
																assign node13799 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node13802 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node13805 = (inp[10]) ? node13807 : 4'b1111;
														assign node13807 = (inp[2]) ? 4'b1110 : node13808;
															assign node13808 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node13812 = (inp[0]) ? node13822 : node13813;
													assign node13813 = (inp[11]) ? node13819 : node13814;
														assign node13814 = (inp[2]) ? 4'b1111 : node13815;
															assign node13815 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13819 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node13822 = (inp[11]) ? node13828 : node13823;
														assign node13823 = (inp[2]) ? 4'b1110 : node13824;
															assign node13824 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node13828 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node13831 = (inp[4]) ? node13851 : node13832;
												assign node13832 = (inp[9]) ? node13844 : node13833;
													assign node13833 = (inp[10]) ? 4'b1011 : node13834;
														assign node13834 = (inp[2]) ? node13836 : 4'b1011;
															assign node13836 = (inp[0]) ? node13840 : node13837;
																assign node13837 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node13840 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13844 = (inp[11]) ? node13846 : 4'b1011;
														assign node13846 = (inp[2]) ? node13848 : 4'b1010;
															assign node13848 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node13851 = (inp[11]) ? node13863 : node13852;
													assign node13852 = (inp[10]) ? node13856 : node13853;
														assign node13853 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node13856 = (inp[0]) ? node13858 : 4'b1110;
															assign node13858 = (inp[9]) ? 4'b1110 : node13859;
																assign node13859 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node13863 = (inp[10]) ? 4'b1111 : node13864;
														assign node13864 = (inp[2]) ? node13870 : node13865;
															assign node13865 = (inp[0]) ? node13867 : 4'b1111;
																assign node13867 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node13870 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node13874 = (inp[1]) ? node13914 : node13875;
											assign node13875 = (inp[4]) ? node13897 : node13876;
												assign node13876 = (inp[10]) ? node13892 : node13877;
													assign node13877 = (inp[0]) ? node13883 : node13878;
														assign node13878 = (inp[11]) ? node13880 : 4'b1100;
															assign node13880 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node13883 = (inp[2]) ? 4'b1101 : node13884;
															assign node13884 = (inp[11]) ? node13888 : node13885;
																assign node13885 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node13888 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13892 = (inp[0]) ? node13894 : 4'b1101;
														assign node13894 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node13897 = (inp[2]) ? node13905 : node13898;
													assign node13898 = (inp[0]) ? 4'b1001 : node13899;
														assign node13899 = (inp[11]) ? node13901 : 4'b1000;
															assign node13901 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13905 = (inp[9]) ? 4'b1000 : node13906;
														assign node13906 = (inp[11]) ? node13910 : node13907;
															assign node13907 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node13910 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node13914 = (inp[10]) ? node13932 : node13915;
												assign node13915 = (inp[2]) ? node13923 : node13916;
													assign node13916 = (inp[4]) ? 4'b1101 : node13917;
														assign node13917 = (inp[11]) ? node13919 : 4'b1101;
															assign node13919 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13923 = (inp[4]) ? node13925 : 4'b1101;
														assign node13925 = (inp[0]) ? 4'b1101 : node13926;
															assign node13926 = (inp[9]) ? 4'b1100 : node13927;
																assign node13927 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node13932 = (inp[0]) ? node13950 : node13933;
													assign node13933 = (inp[2]) ? node13943 : node13934;
														assign node13934 = (inp[11]) ? 4'b1101 : node13935;
															assign node13935 = (inp[4]) ? node13939 : node13936;
																assign node13936 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node13939 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node13943 = (inp[9]) ? node13947 : node13944;
															assign node13944 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13947 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13950 = (inp[9]) ? node13958 : node13951;
														assign node13951 = (inp[11]) ? node13955 : node13952;
															assign node13952 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node13955 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node13958 = (inp[11]) ? 4'b1100 : node13959;
															assign node13959 = (inp[2]) ? 4'b1101 : node13960;
																assign node13960 = (inp[4]) ? 4'b1100 : 4'b1101;
							assign node13965 = (inp[12]) ? node14249 : node13966;
								assign node13966 = (inp[15]) ? node14098 : node13967;
									assign node13967 = (inp[7]) ? node14045 : node13968;
										assign node13968 = (inp[1]) ? node14008 : node13969;
											assign node13969 = (inp[0]) ? node13999 : node13970;
												assign node13970 = (inp[10]) ? node13984 : node13971;
													assign node13971 = (inp[4]) ? 4'b1001 : node13972;
														assign node13972 = (inp[11]) ? node13978 : node13973;
															assign node13973 = (inp[9]) ? 4'b1000 : node13974;
																assign node13974 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node13978 = (inp[2]) ? node13980 : 4'b1001;
																assign node13980 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13984 = (inp[4]) ? node13992 : node13985;
														assign node13985 = (inp[11]) ? node13987 : 4'b1001;
															assign node13987 = (inp[2]) ? node13989 : 4'b1000;
																assign node13989 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node13992 = (inp[11]) ? node13994 : 4'b1000;
															assign node13994 = (inp[2]) ? 4'b1000 : node13995;
																assign node13995 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node13999 = (inp[10]) ? 4'b1001 : node14000;
													assign node14000 = (inp[9]) ? node14004 : node14001;
														assign node14001 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node14004 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node14008 = (inp[0]) ? node14032 : node14009;
												assign node14009 = (inp[9]) ? node14021 : node14010;
													assign node14010 = (inp[2]) ? node14012 : 4'b1001;
														assign node14012 = (inp[10]) ? node14018 : node14013;
															assign node14013 = (inp[4]) ? 4'b1001 : node14014;
																assign node14014 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node14018 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node14021 = (inp[4]) ? node14027 : node14022;
														assign node14022 = (inp[11]) ? 4'b1000 : node14023;
															assign node14023 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14027 = (inp[11]) ? 4'b1001 : node14028;
															assign node14028 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node14032 = (inp[10]) ? node14040 : node14033;
													assign node14033 = (inp[9]) ? node14037 : node14034;
														assign node14034 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node14037 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14040 = (inp[9]) ? node14042 : 4'b1000;
														assign node14042 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node14045 = (inp[9]) ? node14073 : node14046;
											assign node14046 = (inp[11]) ? node14064 : node14047;
												assign node14047 = (inp[0]) ? 4'b1010 : node14048;
													assign node14048 = (inp[1]) ? node14058 : node14049;
														assign node14049 = (inp[10]) ? node14051 : 4'b1011;
															assign node14051 = (inp[4]) ? node14055 : node14052;
																assign node14052 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node14055 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node14058 = (inp[4]) ? node14060 : 4'b1010;
															assign node14060 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node14064 = (inp[0]) ? 4'b1011 : node14065;
													assign node14065 = (inp[2]) ? node14069 : node14066;
														assign node14066 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node14069 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node14073 = (inp[11]) ? node14089 : node14074;
												assign node14074 = (inp[0]) ? 4'b1011 : node14075;
													assign node14075 = (inp[10]) ? node14083 : node14076;
														assign node14076 = (inp[4]) ? node14080 : node14077;
															assign node14077 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node14080 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14083 = (inp[2]) ? 4'b1011 : node14084;
															assign node14084 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node14089 = (inp[0]) ? 4'b1010 : node14090;
													assign node14090 = (inp[4]) ? node14094 : node14091;
														assign node14091 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14094 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node14098 = (inp[7]) ? node14186 : node14099;
										assign node14099 = (inp[4]) ? node14139 : node14100;
											assign node14100 = (inp[11]) ? node14118 : node14101;
												assign node14101 = (inp[9]) ? node14111 : node14102;
													assign node14102 = (inp[0]) ? node14106 : node14103;
														assign node14103 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14106 = (inp[1]) ? node14108 : 4'b1010;
															assign node14108 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node14111 = (inp[2]) ? node14113 : 4'b1011;
														assign node14113 = (inp[0]) ? node14115 : 4'b1011;
															assign node14115 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node14118 = (inp[9]) ? node14134 : node14119;
													assign node14119 = (inp[10]) ? node14127 : node14120;
														assign node14120 = (inp[2]) ? 4'b1010 : node14121;
															assign node14121 = (inp[1]) ? 4'b1011 : node14122;
																assign node14122 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node14127 = (inp[0]) ? node14129 : 4'b1011;
															assign node14129 = (inp[2]) ? node14131 : 4'b1011;
																assign node14131 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node14134 = (inp[2]) ? node14136 : 4'b1010;
														assign node14136 = (inp[1]) ? 4'b1011 : 4'b1010;
											assign node14139 = (inp[1]) ? node14161 : node14140;
												assign node14140 = (inp[2]) ? node14148 : node14141;
													assign node14141 = (inp[11]) ? node14145 : node14142;
														assign node14142 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14145 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node14148 = (inp[9]) ? node14154 : node14149;
														assign node14149 = (inp[11]) ? 4'b1010 : node14150;
															assign node14150 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node14154 = (inp[0]) ? node14158 : node14155;
															assign node14155 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node14158 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node14161 = (inp[0]) ? node14169 : node14162;
													assign node14162 = (inp[10]) ? 4'b1110 : node14163;
														assign node14163 = (inp[11]) ? 4'b1111 : node14164;
															assign node14164 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node14169 = (inp[2]) ? node14179 : node14170;
														assign node14170 = (inp[10]) ? 4'b1111 : node14171;
															assign node14171 = (inp[9]) ? node14175 : node14172;
																assign node14172 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node14175 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node14179 = (inp[11]) ? node14183 : node14180;
															assign node14180 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14183 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node14186 = (inp[4]) ? node14222 : node14187;
											assign node14187 = (inp[1]) ? node14205 : node14188;
												assign node14188 = (inp[2]) ? node14198 : node14189;
													assign node14189 = (inp[9]) ? node14191 : 4'b1101;
														assign node14191 = (inp[10]) ? node14193 : 4'b1100;
															assign node14193 = (inp[0]) ? 4'b1101 : node14194;
																assign node14194 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node14198 = (inp[11]) ? node14202 : node14199;
														assign node14199 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14202 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node14205 = (inp[11]) ? node14217 : node14206;
													assign node14206 = (inp[9]) ? node14212 : node14207;
														assign node14207 = (inp[0]) ? 4'b1000 : node14208;
															assign node14208 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14212 = (inp[0]) ? 4'b1001 : node14213;
															assign node14213 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node14217 = (inp[2]) ? 4'b1001 : node14218;
														assign node14218 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node14222 = (inp[2]) ? node14234 : node14223;
												assign node14223 = (inp[0]) ? node14227 : node14224;
													assign node14224 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node14227 = (inp[11]) ? node14231 : node14228;
														assign node14228 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14231 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node14234 = (inp[9]) ? node14242 : node14235;
													assign node14235 = (inp[11]) ? node14239 : node14236;
														assign node14236 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14239 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14242 = (inp[11]) ? 4'b1001 : node14243;
														assign node14243 = (inp[0]) ? node14245 : 4'b1000;
															assign node14245 = (inp[1]) ? 4'b1001 : 4'b1000;
								assign node14249 = (inp[15]) ? node14427 : node14250;
									assign node14250 = (inp[7]) ? node14340 : node14251;
										assign node14251 = (inp[11]) ? node14289 : node14252;
											assign node14252 = (inp[2]) ? node14272 : node14253;
												assign node14253 = (inp[9]) ? node14265 : node14254;
													assign node14254 = (inp[1]) ? node14258 : node14255;
														assign node14255 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node14258 = (inp[4]) ? node14262 : node14259;
															assign node14259 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node14262 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14265 = (inp[0]) ? node14267 : 4'b1100;
														assign node14267 = (inp[4]) ? node14269 : 4'b1101;
															assign node14269 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node14272 = (inp[9]) ? node14280 : node14273;
													assign node14273 = (inp[4]) ? node14277 : node14274;
														assign node14274 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node14277 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node14280 = (inp[1]) ? node14286 : node14281;
														assign node14281 = (inp[4]) ? node14283 : 4'b1000;
															assign node14283 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node14286 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node14289 = (inp[10]) ? node14321 : node14290;
												assign node14290 = (inp[0]) ? node14310 : node14291;
													assign node14291 = (inp[2]) ? node14301 : node14292;
														assign node14292 = (inp[4]) ? node14296 : node14293;
															assign node14293 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node14296 = (inp[1]) ? node14298 : 4'b1101;
																assign node14298 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node14301 = (inp[9]) ? node14307 : node14302;
															assign node14302 = (inp[4]) ? node14304 : 4'b1101;
																assign node14304 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node14307 = (inp[4]) ? 4'b1100 : 4'b1001;
													assign node14310 = (inp[9]) ? node14312 : 4'b1000;
														assign node14312 = (inp[1]) ? node14316 : node14313;
															assign node14313 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node14316 = (inp[4]) ? node14318 : 4'b1100;
																assign node14318 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node14321 = (inp[9]) ? node14325 : node14322;
													assign node14322 = (inp[0]) ? 4'b1101 : 4'b1001;
													assign node14325 = (inp[0]) ? node14335 : node14326;
														assign node14326 = (inp[4]) ? node14332 : node14327;
															assign node14327 = (inp[1]) ? 4'b1101 : node14328;
																assign node14328 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node14332 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node14335 = (inp[2]) ? node14337 : 4'b1001;
															assign node14337 = (inp[1]) ? 4'b1100 : 4'b1001;
										assign node14340 = (inp[4]) ? node14382 : node14341;
											assign node14341 = (inp[1]) ? node14363 : node14342;
												assign node14342 = (inp[10]) ? node14356 : node14343;
													assign node14343 = (inp[2]) ? 4'b1011 : node14344;
														assign node14344 = (inp[0]) ? node14350 : node14345;
															assign node14345 = (inp[11]) ? 4'b1010 : node14346;
																assign node14346 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14350 = (inp[11]) ? node14352 : 4'b1010;
																assign node14352 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node14356 = (inp[2]) ? 4'b1010 : node14357;
														assign node14357 = (inp[9]) ? node14359 : 4'b1011;
															assign node14359 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node14363 = (inp[10]) ? node14369 : node14364;
													assign node14364 = (inp[9]) ? node14366 : 4'b1110;
														assign node14366 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node14369 = (inp[2]) ? node14377 : node14370;
														assign node14370 = (inp[0]) ? node14372 : 4'b1111;
															assign node14372 = (inp[11]) ? node14374 : 4'b1110;
																assign node14374 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14377 = (inp[0]) ? node14379 : 4'b1110;
															assign node14379 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node14382 = (inp[1]) ? node14400 : node14383;
												assign node14383 = (inp[9]) ? node14389 : node14384;
													assign node14384 = (inp[11]) ? 4'b1111 : node14385;
														assign node14385 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node14389 = (inp[2]) ? 4'b1110 : node14390;
														assign node14390 = (inp[10]) ? 4'b1111 : node14391;
															assign node14391 = (inp[0]) ? node14395 : node14392;
																assign node14392 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node14395 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node14400 = (inp[10]) ? node14410 : node14401;
													assign node14401 = (inp[2]) ? node14407 : node14402;
														assign node14402 = (inp[9]) ? 4'b1011 : node14403;
															assign node14403 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node14407 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node14410 = (inp[2]) ? node14418 : node14411;
														assign node14411 = (inp[11]) ? node14415 : node14412;
															assign node14412 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14415 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node14418 = (inp[11]) ? node14420 : 4'b1011;
															assign node14420 = (inp[0]) ? node14424 : node14421;
																assign node14421 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node14424 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node14427 = (inp[7]) ? node14517 : node14428;
										assign node14428 = (inp[4]) ? node14466 : node14429;
											assign node14429 = (inp[1]) ? node14449 : node14430;
												assign node14430 = (inp[9]) ? node14438 : node14431;
													assign node14431 = (inp[11]) ? 4'b1011 : node14432;
														assign node14432 = (inp[2]) ? 4'b1010 : node14433;
															assign node14433 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node14438 = (inp[11]) ? node14444 : node14439;
														assign node14439 = (inp[10]) ? 4'b1011 : node14440;
															assign node14440 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node14444 = (inp[2]) ? 4'b1010 : node14445;
															assign node14445 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node14449 = (inp[2]) ? node14461 : node14450;
													assign node14450 = (inp[10]) ? node14458 : node14451;
														assign node14451 = (inp[0]) ? 4'b1110 : node14452;
															assign node14452 = (inp[11]) ? 4'b1110 : node14453;
																assign node14453 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node14458 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node14461 = (inp[11]) ? 4'b1111 : node14462;
														assign node14462 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node14466 = (inp[9]) ? node14494 : node14467;
												assign node14467 = (inp[10]) ? node14479 : node14468;
													assign node14468 = (inp[0]) ? node14474 : node14469;
														assign node14469 = (inp[1]) ? 4'b1010 : node14470;
															assign node14470 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node14474 = (inp[1]) ? 4'b1011 : node14475;
															assign node14475 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node14479 = (inp[0]) ? node14487 : node14480;
														assign node14480 = (inp[2]) ? node14484 : node14481;
															assign node14481 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node14484 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node14487 = (inp[2]) ? 4'b1010 : node14488;
															assign node14488 = (inp[11]) ? 4'b1010 : node14489;
																assign node14489 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node14494 = (inp[11]) ? node14504 : node14495;
													assign node14495 = (inp[2]) ? node14499 : node14496;
														assign node14496 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node14499 = (inp[1]) ? node14501 : 4'b1011;
															assign node14501 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node14504 = (inp[10]) ? node14510 : node14505;
														assign node14505 = (inp[1]) ? 4'b1010 : node14506;
															assign node14506 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14510 = (inp[1]) ? node14514 : node14511;
															assign node14511 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node14514 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node14517 = (inp[1]) ? node14557 : node14518;
											assign node14518 = (inp[4]) ? node14532 : node14519;
												assign node14519 = (inp[11]) ? node14525 : node14520;
													assign node14520 = (inp[10]) ? node14522 : 4'b1001;
														assign node14522 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node14525 = (inp[9]) ? 4'b1000 : node14526;
														assign node14526 = (inp[0]) ? 4'b1001 : node14527;
															assign node14527 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node14532 = (inp[2]) ? node14540 : node14533;
													assign node14533 = (inp[11]) ? node14537 : node14534;
														assign node14534 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node14537 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node14540 = (inp[10]) ? node14550 : node14541;
														assign node14541 = (inp[11]) ? 4'b1101 : node14542;
															assign node14542 = (inp[9]) ? node14546 : node14543;
																assign node14543 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node14546 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14550 = (inp[0]) ? node14552 : 4'b1100;
															assign node14552 = (inp[9]) ? node14554 : 4'b1101;
																assign node14554 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node14557 = (inp[9]) ? node14581 : node14558;
												assign node14558 = (inp[2]) ? node14564 : node14559;
													assign node14559 = (inp[10]) ? 4'b1001 : node14560;
														assign node14560 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node14564 = (inp[4]) ? node14570 : node14565;
														assign node14565 = (inp[11]) ? 4'b1001 : node14566;
															assign node14566 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14570 = (inp[10]) ? node14576 : node14571;
															assign node14571 = (inp[0]) ? node14573 : 4'b1000;
																assign node14573 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node14576 = (inp[11]) ? 4'b1000 : node14577;
																assign node14577 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node14581 = (inp[0]) ? node14593 : node14582;
													assign node14582 = (inp[11]) ? node14588 : node14583;
														assign node14583 = (inp[10]) ? 4'b1000 : node14584;
															assign node14584 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14588 = (inp[10]) ? 4'b1001 : node14589;
															assign node14589 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node14593 = (inp[2]) ? 4'b1000 : node14594;
														assign node14594 = (inp[10]) ? node14598 : node14595;
															assign node14595 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node14598 = (inp[11]) ? 4'b1000 : node14599;
																assign node14599 = (inp[4]) ? 4'b1001 : 4'b1000;
					assign node14604 = (inp[15]) ? node15364 : node14605;
						assign node14605 = (inp[13]) ? node14909 : node14606;
							assign node14606 = (inp[12]) ? node14696 : node14607;
								assign node14607 = (inp[9]) ? node14665 : node14608;
									assign node14608 = (inp[5]) ? node14622 : node14609;
										assign node14609 = (inp[4]) ? node14617 : node14610;
											assign node14610 = (inp[7]) ? node14614 : node14611;
												assign node14611 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node14614 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node14617 = (inp[7]) ? node14619 : 4'b0010;
												assign node14619 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node14622 = (inp[7]) ? node14634 : node14623;
											assign node14623 = (inp[4]) ? 4'b0011 : node14624;
												assign node14624 = (inp[11]) ? node14626 : 4'b0000;
													assign node14626 = (inp[2]) ? node14630 : node14627;
														assign node14627 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node14630 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node14634 = (inp[4]) ? node14662 : node14635;
												assign node14635 = (inp[10]) ? node14655 : node14636;
													assign node14636 = (inp[1]) ? node14644 : node14637;
														assign node14637 = (inp[11]) ? 4'b0011 : node14638;
															assign node14638 = (inp[2]) ? 4'b0011 : node14639;
																assign node14639 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node14644 = (inp[11]) ? node14650 : node14645;
															assign node14645 = (inp[0]) ? node14647 : 4'b0011;
																assign node14647 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node14650 = (inp[2]) ? node14652 : 4'b0010;
																assign node14652 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node14655 = (inp[0]) ? node14659 : node14656;
														assign node14656 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node14659 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node14662 = (inp[1]) ? 4'b0100 : 4'b0000;
									assign node14665 = (inp[7]) ? node14681 : node14666;
										assign node14666 = (inp[4]) ? node14678 : node14667;
											assign node14667 = (inp[2]) ? node14673 : node14668;
												assign node14668 = (inp[0]) ? node14670 : 4'b0001;
													assign node14670 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node14673 = (inp[0]) ? node14675 : 4'b0000;
													assign node14675 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node14678 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node14681 = (inp[4]) ? node14693 : node14682;
											assign node14682 = (inp[2]) ? node14688 : node14683;
												assign node14683 = (inp[0]) ? 4'b0011 : node14684;
													assign node14684 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node14688 = (inp[0]) ? 4'b0010 : node14689;
													assign node14689 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node14693 = (inp[1]) ? 4'b0101 : 4'b0001;
								assign node14696 = (inp[4]) ? node14830 : node14697;
									assign node14697 = (inp[7]) ? node14765 : node14698;
										assign node14698 = (inp[2]) ? node14740 : node14699;
											assign node14699 = (inp[0]) ? node14719 : node14700;
												assign node14700 = (inp[5]) ? node14708 : node14701;
													assign node14701 = (inp[11]) ? 4'b0100 : node14702;
														assign node14702 = (inp[9]) ? 4'b0101 : node14703;
															assign node14703 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node14708 = (inp[11]) ? node14716 : node14709;
														assign node14709 = (inp[9]) ? node14713 : node14710;
															assign node14710 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node14713 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node14716 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node14719 = (inp[5]) ? node14733 : node14720;
													assign node14720 = (inp[10]) ? node14726 : node14721;
														assign node14721 = (inp[1]) ? 4'b0101 : node14722;
															assign node14722 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node14726 = (inp[1]) ? node14730 : node14727;
															assign node14727 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node14730 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node14733 = (inp[9]) ? node14737 : node14734;
														assign node14734 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node14737 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node14740 = (inp[0]) ? node14754 : node14741;
												assign node14741 = (inp[11]) ? node14749 : node14742;
													assign node14742 = (inp[9]) ? node14746 : node14743;
														assign node14743 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node14746 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node14749 = (inp[9]) ? 4'b0101 : node14750;
														assign node14750 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node14754 = (inp[1]) ? node14760 : node14755;
													assign node14755 = (inp[5]) ? node14757 : 4'b0101;
														assign node14757 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node14760 = (inp[5]) ? node14762 : 4'b0100;
														assign node14762 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node14765 = (inp[11]) ? node14805 : node14766;
											assign node14766 = (inp[10]) ? node14782 : node14767;
												assign node14767 = (inp[0]) ? node14775 : node14768;
													assign node14768 = (inp[5]) ? node14770 : 4'b0111;
														assign node14770 = (inp[1]) ? 4'b0111 : node14771;
															assign node14771 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node14775 = (inp[5]) ? 4'b0111 : node14776;
														assign node14776 = (inp[2]) ? node14778 : 4'b0110;
															assign node14778 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node14782 = (inp[1]) ? node14792 : node14783;
													assign node14783 = (inp[9]) ? node14787 : node14784;
														assign node14784 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node14787 = (inp[2]) ? 4'b0110 : node14788;
															assign node14788 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node14792 = (inp[5]) ? node14800 : node14793;
														assign node14793 = (inp[2]) ? 4'b0110 : node14794;
															assign node14794 = (inp[9]) ? 4'b0111 : node14795;
																assign node14795 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node14800 = (inp[9]) ? node14802 : 4'b0111;
															assign node14802 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node14805 = (inp[1]) ? node14821 : node14806;
												assign node14806 = (inp[5]) ? node14812 : node14807;
													assign node14807 = (inp[9]) ? 4'b0111 : node14808;
														assign node14808 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node14812 = (inp[0]) ? node14818 : node14813;
														assign node14813 = (inp[10]) ? 4'b0110 : node14814;
															assign node14814 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node14818 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node14821 = (inp[10]) ? node14823 : 4'b0110;
													assign node14823 = (inp[5]) ? node14827 : node14824;
														assign node14824 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node14827 = (inp[2]) ? 4'b0110 : 4'b0111;
									assign node14830 = (inp[7]) ? node14902 : node14831;
										assign node14831 = (inp[10]) ? node14857 : node14832;
											assign node14832 = (inp[0]) ? node14846 : node14833;
												assign node14833 = (inp[9]) ? node14839 : node14834;
													assign node14834 = (inp[1]) ? node14836 : 4'b0011;
														assign node14836 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node14839 = (inp[1]) ? node14843 : node14840;
														assign node14840 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node14843 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node14846 = (inp[5]) ? 4'b0011 : node14847;
													assign node14847 = (inp[11]) ? node14849 : 4'b0010;
														assign node14849 = (inp[1]) ? node14853 : node14850;
															assign node14850 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node14853 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node14857 = (inp[11]) ? node14881 : node14858;
												assign node14858 = (inp[2]) ? node14872 : node14859;
													assign node14859 = (inp[5]) ? node14865 : node14860;
														assign node14860 = (inp[9]) ? node14862 : 4'b0010;
															assign node14862 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node14865 = (inp[0]) ? 4'b0010 : node14866;
															assign node14866 = (inp[1]) ? 4'b0011 : node14867;
																assign node14867 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node14872 = (inp[1]) ? 4'b0011 : node14873;
														assign node14873 = (inp[9]) ? node14877 : node14874;
															assign node14874 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node14877 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node14881 = (inp[9]) ? node14889 : node14882;
													assign node14882 = (inp[1]) ? 4'b0011 : node14883;
														assign node14883 = (inp[5]) ? 4'b0010 : node14884;
															assign node14884 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node14889 = (inp[1]) ? 4'b0010 : node14890;
														assign node14890 = (inp[2]) ? node14896 : node14891;
															assign node14891 = (inp[0]) ? 4'b0010 : node14892;
																assign node14892 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node14896 = (inp[0]) ? node14898 : 4'b0010;
																assign node14898 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node14902 = (inp[1]) ? node14906 : node14903;
											assign node14903 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node14906 = (inp[9]) ? 4'b0101 : 4'b0100;
							assign node14909 = (inp[12]) ? node15091 : node14910;
								assign node14910 = (inp[7]) ? node15022 : node14911;
									assign node14911 = (inp[4]) ? node14977 : node14912;
										assign node14912 = (inp[10]) ? node14958 : node14913;
											assign node14913 = (inp[11]) ? node14933 : node14914;
												assign node14914 = (inp[9]) ? node14926 : node14915;
													assign node14915 = (inp[2]) ? node14921 : node14916;
														assign node14916 = (inp[0]) ? node14918 : 4'b0100;
															assign node14918 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node14921 = (inp[5]) ? node14923 : 4'b0101;
															assign node14923 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node14926 = (inp[2]) ? node14928 : 4'b0101;
														assign node14928 = (inp[5]) ? node14930 : 4'b0100;
															assign node14930 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node14933 = (inp[0]) ? node14947 : node14934;
													assign node14934 = (inp[1]) ? node14942 : node14935;
														assign node14935 = (inp[9]) ? node14939 : node14936;
															assign node14936 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node14939 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node14942 = (inp[2]) ? node14944 : 4'b0101;
															assign node14944 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node14947 = (inp[2]) ? 4'b0100 : node14948;
														assign node14948 = (inp[1]) ? 4'b0100 : node14949;
															assign node14949 = (inp[9]) ? node14953 : node14950;
																assign node14950 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node14953 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node14958 = (inp[2]) ? node14970 : node14959;
												assign node14959 = (inp[9]) ? node14965 : node14960;
													assign node14960 = (inp[0]) ? node14962 : 4'b0100;
														assign node14962 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node14965 = (inp[5]) ? node14967 : 4'b0101;
														assign node14967 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node14970 = (inp[9]) ? node14972 : 4'b0101;
													assign node14972 = (inp[0]) ? node14974 : 4'b0100;
														assign node14974 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node14977 = (inp[0]) ? node15001 : node14978;
											assign node14978 = (inp[11]) ? node14994 : node14979;
												assign node14979 = (inp[10]) ? node14987 : node14980;
													assign node14980 = (inp[9]) ? node14984 : node14981;
														assign node14981 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node14984 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node14987 = (inp[5]) ? node14991 : node14988;
														assign node14988 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node14991 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node14994 = (inp[5]) ? node14998 : node14995;
													assign node14995 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node14998 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node15001 = (inp[1]) ? node15015 : node15002;
												assign node15002 = (inp[2]) ? node15008 : node15003;
													assign node15003 = (inp[9]) ? node15005 : 4'b0111;
														assign node15005 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node15008 = (inp[9]) ? node15012 : node15009;
														assign node15009 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node15012 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node15015 = (inp[9]) ? node15019 : node15016;
													assign node15016 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node15019 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node15022 = (inp[4]) ? node15064 : node15023;
										assign node15023 = (inp[5]) ? node15029 : node15024;
											assign node15024 = (inp[2]) ? 4'b0110 : node15025;
												assign node15025 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node15029 = (inp[10]) ? node15051 : node15030;
												assign node15030 = (inp[2]) ? node15040 : node15031;
													assign node15031 = (inp[1]) ? 4'b0111 : node15032;
														assign node15032 = (inp[0]) ? node15036 : node15033;
															assign node15033 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node15036 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node15040 = (inp[1]) ? node15046 : node15041;
														assign node15041 = (inp[0]) ? 4'b0111 : node15042;
															assign node15042 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node15046 = (inp[9]) ? 4'b0110 : node15047;
															assign node15047 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node15051 = (inp[9]) ? node15059 : node15052;
													assign node15052 = (inp[2]) ? node15056 : node15053;
														assign node15053 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node15056 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node15059 = (inp[2]) ? node15061 : 4'b0110;
														assign node15061 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node15064 = (inp[1]) ? node15068 : node15065;
											assign node15065 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node15068 = (inp[2]) ? node15082 : node15069;
												assign node15069 = (inp[10]) ? node15075 : node15070;
													assign node15070 = (inp[0]) ? node15072 : 4'b0001;
														assign node15072 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15075 = (inp[9]) ? node15079 : node15076;
														assign node15076 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node15079 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node15082 = (inp[10]) ? node15084 : 4'b0000;
													assign node15084 = (inp[0]) ? node15088 : node15085;
														assign node15085 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node15088 = (inp[9]) ? 4'b0000 : 4'b0001;
								assign node15091 = (inp[4]) ? node15263 : node15092;
									assign node15092 = (inp[7]) ? node15184 : node15093;
										assign node15093 = (inp[11]) ? node15149 : node15094;
											assign node15094 = (inp[2]) ? node15124 : node15095;
												assign node15095 = (inp[10]) ? node15111 : node15096;
													assign node15096 = (inp[9]) ? node15106 : node15097;
														assign node15097 = (inp[0]) ? 4'b0001 : node15098;
															assign node15098 = (inp[5]) ? node15102 : node15099;
																assign node15099 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node15102 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node15106 = (inp[1]) ? 4'b0001 : node15107;
															assign node15107 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node15111 = (inp[9]) ? node15119 : node15112;
														assign node15112 = (inp[0]) ? node15116 : node15113;
															assign node15113 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node15116 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node15119 = (inp[0]) ? node15121 : 4'b0000;
															assign node15121 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node15124 = (inp[10]) ? node15130 : node15125;
													assign node15125 = (inp[0]) ? 4'b0000 : node15126;
														assign node15126 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15130 = (inp[0]) ? node15142 : node15131;
														assign node15131 = (inp[5]) ? node15137 : node15132;
															assign node15132 = (inp[9]) ? 4'b0000 : node15133;
																assign node15133 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node15137 = (inp[9]) ? 4'b0001 : node15138;
																assign node15138 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node15142 = (inp[1]) ? node15146 : node15143;
															assign node15143 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node15146 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node15149 = (inp[2]) ? node15173 : node15150;
												assign node15150 = (inp[5]) ? node15166 : node15151;
													assign node15151 = (inp[10]) ? node15163 : node15152;
														assign node15152 = (inp[0]) ? node15158 : node15153;
															assign node15153 = (inp[9]) ? 4'b0000 : node15154;
																assign node15154 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node15158 = (inp[9]) ? 4'b0001 : node15159;
																assign node15159 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node15163 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node15166 = (inp[9]) ? node15170 : node15167;
														assign node15167 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node15170 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node15173 = (inp[10]) ? node15175 : 4'b0001;
													assign node15175 = (inp[1]) ? node15181 : node15176;
														assign node15176 = (inp[9]) ? 4'b0001 : node15177;
															assign node15177 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node15181 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node15184 = (inp[1]) ? node15228 : node15185;
											assign node15185 = (inp[5]) ? node15199 : node15186;
												assign node15186 = (inp[0]) ? node15192 : node15187;
													assign node15187 = (inp[10]) ? node15189 : 4'b0011;
														assign node15189 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node15192 = (inp[2]) ? node15196 : node15193;
														assign node15193 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node15196 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node15199 = (inp[2]) ? node15217 : node15200;
													assign node15200 = (inp[11]) ? node15212 : node15201;
														assign node15201 = (inp[10]) ? node15207 : node15202;
															assign node15202 = (inp[9]) ? 4'b0010 : node15203;
																assign node15203 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node15207 = (inp[9]) ? 4'b0011 : node15208;
																assign node15208 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node15212 = (inp[0]) ? node15214 : 4'b0011;
															assign node15214 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node15217 = (inp[11]) ? node15219 : 4'b0011;
														assign node15219 = (inp[10]) ? 4'b0011 : node15220;
															assign node15220 = (inp[9]) ? node15224 : node15221;
																assign node15221 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node15224 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node15228 = (inp[0]) ? node15250 : node15229;
												assign node15229 = (inp[11]) ? node15235 : node15230;
													assign node15230 = (inp[9]) ? 4'b0010 : node15231;
														assign node15231 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node15235 = (inp[10]) ? node15241 : node15236;
														assign node15236 = (inp[2]) ? 4'b0011 : node15237;
															assign node15237 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node15241 = (inp[9]) ? node15243 : 4'b0010;
															assign node15243 = (inp[2]) ? node15247 : node15244;
																assign node15244 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node15247 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node15250 = (inp[5]) ? node15256 : node15251;
													assign node15251 = (inp[9]) ? 4'b0011 : node15252;
														assign node15252 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node15256 = (inp[2]) ? node15260 : node15257;
														assign node15257 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node15260 = (inp[9]) ? 4'b0010 : 4'b0011;
									assign node15263 = (inp[7]) ? node15331 : node15264;
										assign node15264 = (inp[0]) ? node15304 : node15265;
											assign node15265 = (inp[5]) ? node15281 : node15266;
												assign node15266 = (inp[11]) ? node15274 : node15267;
													assign node15267 = (inp[9]) ? node15271 : node15268;
														assign node15268 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node15271 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node15274 = (inp[2]) ? node15276 : 4'b0110;
														assign node15276 = (inp[10]) ? node15278 : 4'b0110;
															assign node15278 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node15281 = (inp[11]) ? node15289 : node15282;
													assign node15282 = (inp[1]) ? node15286 : node15283;
														assign node15283 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node15286 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node15289 = (inp[10]) ? node15295 : node15290;
														assign node15290 = (inp[9]) ? 4'b0110 : node15291;
															assign node15291 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node15295 = (inp[2]) ? node15297 : 4'b0111;
															assign node15297 = (inp[1]) ? node15301 : node15298;
																assign node15298 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node15301 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node15304 = (inp[5]) ? node15312 : node15305;
												assign node15305 = (inp[9]) ? node15309 : node15306;
													assign node15306 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node15309 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node15312 = (inp[11]) ? node15320 : node15313;
													assign node15313 = (inp[1]) ? node15317 : node15314;
														assign node15314 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node15317 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node15320 = (inp[2]) ? node15326 : node15321;
														assign node15321 = (inp[9]) ? 4'b0110 : node15322;
															assign node15322 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node15326 = (inp[9]) ? node15328 : 4'b0110;
															assign node15328 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node15331 = (inp[1]) ? node15335 : node15332;
											assign node15332 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node15335 = (inp[11]) ? node15357 : node15336;
												assign node15336 = (inp[10]) ? node15350 : node15337;
													assign node15337 = (inp[2]) ? node15345 : node15338;
														assign node15338 = (inp[9]) ? node15342 : node15339;
															assign node15339 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node15342 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node15345 = (inp[0]) ? 4'b0001 : node15346;
															assign node15346 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15350 = (inp[0]) ? node15354 : node15351;
														assign node15351 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node15354 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node15357 = (inp[9]) ? node15361 : node15358;
													assign node15358 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15361 = (inp[0]) ? 4'b0000 : 4'b0001;
						assign node15364 = (inp[13]) ? node15782 : node15365;
							assign node15365 = (inp[4]) ? node15623 : node15366;
								assign node15366 = (inp[7]) ? node15468 : node15367;
									assign node15367 = (inp[1]) ? node15425 : node15368;
										assign node15368 = (inp[12]) ? node15388 : node15369;
											assign node15369 = (inp[2]) ? node15381 : node15370;
												assign node15370 = (inp[9]) ? node15376 : node15371;
													assign node15371 = (inp[5]) ? node15373 : 4'b0000;
														assign node15373 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15376 = (inp[5]) ? node15378 : 4'b0001;
														assign node15378 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node15381 = (inp[9]) ? 4'b0000 : node15382;
													assign node15382 = (inp[5]) ? node15384 : 4'b0001;
														assign node15384 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node15388 = (inp[5]) ? node15398 : node15389;
												assign node15389 = (inp[0]) ? node15391 : 4'b0100;
													assign node15391 = (inp[10]) ? 4'b0100 : node15392;
														assign node15392 = (inp[2]) ? 4'b0101 : node15393;
															assign node15393 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node15398 = (inp[11]) ? node15412 : node15399;
													assign node15399 = (inp[0]) ? node15407 : node15400;
														assign node15400 = (inp[10]) ? 4'b0101 : node15401;
															assign node15401 = (inp[9]) ? 4'b0100 : node15402;
																assign node15402 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node15407 = (inp[10]) ? 4'b0100 : node15408;
															assign node15408 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node15412 = (inp[2]) ? node15414 : 4'b0101;
														assign node15414 = (inp[10]) ? node15420 : node15415;
															assign node15415 = (inp[9]) ? node15417 : 4'b0101;
																assign node15417 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node15420 = (inp[9]) ? node15422 : 4'b0100;
																assign node15422 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node15425 = (inp[12]) ? node15449 : node15426;
											assign node15426 = (inp[2]) ? node15438 : node15427;
												assign node15427 = (inp[9]) ? node15433 : node15428;
													assign node15428 = (inp[0]) ? 4'b0101 : node15429;
														assign node15429 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node15433 = (inp[0]) ? 4'b0100 : node15434;
														assign node15434 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node15438 = (inp[9]) ? node15444 : node15439;
													assign node15439 = (inp[5]) ? 4'b0100 : node15440;
														assign node15440 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node15444 = (inp[5]) ? 4'b0101 : node15445;
														assign node15445 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node15449 = (inp[9]) ? node15461 : node15450;
												assign node15450 = (inp[2]) ? node15456 : node15451;
													assign node15451 = (inp[5]) ? node15453 : 4'b0000;
														assign node15453 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15456 = (inp[0]) ? node15458 : 4'b0001;
														assign node15458 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node15461 = (inp[2]) ? 4'b0000 : node15462;
													assign node15462 = (inp[0]) ? node15464 : 4'b0001;
														assign node15464 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node15468 = (inp[5]) ? node15540 : node15469;
										assign node15469 = (inp[12]) ? node15493 : node15470;
											assign node15470 = (inp[1]) ? node15486 : node15471;
												assign node15471 = (inp[11]) ? node15479 : node15472;
													assign node15472 = (inp[9]) ? node15476 : node15473;
														assign node15473 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node15476 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node15479 = (inp[2]) ? node15483 : node15480;
														assign node15480 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node15483 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node15486 = (inp[2]) ? node15490 : node15487;
													assign node15487 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node15490 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node15493 = (inp[1]) ? node15517 : node15494;
												assign node15494 = (inp[11]) ? node15508 : node15495;
													assign node15495 = (inp[0]) ? node15503 : node15496;
														assign node15496 = (inp[10]) ? node15498 : 4'b0011;
															assign node15498 = (inp[2]) ? 4'b0010 : node15499;
																assign node15499 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node15503 = (inp[2]) ? node15505 : 4'b0010;
															assign node15505 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node15508 = (inp[0]) ? node15510 : 4'b0010;
														assign node15510 = (inp[2]) ? node15514 : node15511;
															assign node15511 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node15514 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node15517 = (inp[11]) ? node15525 : node15518;
													assign node15518 = (inp[2]) ? 4'b0111 : node15519;
														assign node15519 = (inp[0]) ? 4'b0110 : node15520;
															assign node15520 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node15525 = (inp[2]) ? node15535 : node15526;
														assign node15526 = (inp[10]) ? node15528 : 4'b0111;
															assign node15528 = (inp[9]) ? node15532 : node15529;
																assign node15529 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node15532 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node15535 = (inp[0]) ? node15537 : 4'b0110;
															assign node15537 = (inp[9]) ? 4'b0111 : 4'b0110;
										assign node15540 = (inp[11]) ? node15578 : node15541;
											assign node15541 = (inp[9]) ? node15555 : node15542;
												assign node15542 = (inp[2]) ? node15548 : node15543;
													assign node15543 = (inp[0]) ? 4'b0110 : node15544;
														assign node15544 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node15548 = (inp[12]) ? node15550 : 4'b0111;
														assign node15550 = (inp[0]) ? 4'b0010 : node15551;
															assign node15551 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node15555 = (inp[2]) ? node15567 : node15556;
													assign node15556 = (inp[1]) ? node15564 : node15557;
														assign node15557 = (inp[12]) ? node15561 : node15558;
															assign node15558 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node15561 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node15564 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node15567 = (inp[0]) ? node15573 : node15568;
														assign node15568 = (inp[1]) ? node15570 : 4'b0111;
															assign node15570 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node15573 = (inp[12]) ? node15575 : 4'b0011;
															assign node15575 = (inp[1]) ? 4'b0110 : 4'b0011;
											assign node15578 = (inp[10]) ? node15594 : node15579;
												assign node15579 = (inp[9]) ? node15585 : node15580;
													assign node15580 = (inp[0]) ? node15582 : 4'b0011;
														assign node15582 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node15585 = (inp[2]) ? node15587 : 4'b0011;
														assign node15587 = (inp[1]) ? 4'b0110 : node15588;
															assign node15588 = (inp[12]) ? 4'b0011 : node15589;
																assign node15589 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node15594 = (inp[1]) ? node15612 : node15595;
													assign node15595 = (inp[12]) ? node15601 : node15596;
														assign node15596 = (inp[0]) ? node15598 : 4'b0110;
															assign node15598 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node15601 = (inp[0]) ? node15607 : node15602;
															assign node15602 = (inp[9]) ? node15604 : 4'b0011;
																assign node15604 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node15607 = (inp[2]) ? node15609 : 4'b0010;
																assign node15609 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node15612 = (inp[12]) ? node15616 : node15613;
														assign node15613 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node15616 = (inp[2]) ? node15620 : node15617;
															assign node15617 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node15620 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node15623 = (inp[7]) ? node15725 : node15624;
									assign node15624 = (inp[0]) ? node15632 : node15625;
										assign node15625 = (inp[9]) ? node15629 : node15626;
											assign node15626 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node15629 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node15632 = (inp[11]) ? node15678 : node15633;
											assign node15633 = (inp[9]) ? node15653 : node15634;
												assign node15634 = (inp[5]) ? node15640 : node15635;
													assign node15635 = (inp[12]) ? node15637 : 4'b0110;
														assign node15637 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node15640 = (inp[2]) ? node15646 : node15641;
														assign node15641 = (inp[1]) ? 4'b0110 : node15642;
															assign node15642 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node15646 = (inp[1]) ? node15650 : node15647;
															assign node15647 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node15650 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node15653 = (inp[5]) ? node15663 : node15654;
													assign node15654 = (inp[2]) ? 4'b0111 : node15655;
														assign node15655 = (inp[10]) ? 4'b0111 : node15656;
															assign node15656 = (inp[1]) ? node15658 : 4'b0110;
																assign node15658 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node15663 = (inp[10]) ? node15671 : node15664;
														assign node15664 = (inp[1]) ? node15668 : node15665;
															assign node15665 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node15668 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node15671 = (inp[1]) ? node15675 : node15672;
															assign node15672 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node15675 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node15678 = (inp[10]) ? node15702 : node15679;
												assign node15679 = (inp[12]) ? node15689 : node15680;
													assign node15680 = (inp[1]) ? node15682 : 4'b0111;
														assign node15682 = (inp[9]) ? node15686 : node15683;
															assign node15683 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node15686 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node15689 = (inp[1]) ? node15697 : node15690;
														assign node15690 = (inp[9]) ? node15694 : node15691;
															assign node15691 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node15694 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node15697 = (inp[5]) ? node15699 : 4'b0111;
															assign node15699 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node15702 = (inp[5]) ? node15712 : node15703;
													assign node15703 = (inp[1]) ? 4'b0111 : node15704;
														assign node15704 = (inp[12]) ? node15708 : node15705;
															assign node15705 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node15708 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node15712 = (inp[9]) ? node15718 : node15713;
														assign node15713 = (inp[1]) ? node15715 : 4'b0110;
															assign node15715 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node15718 = (inp[1]) ? node15722 : node15719;
															assign node15719 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node15722 = (inp[12]) ? 4'b0110 : 4'b0111;
									assign node15725 = (inp[1]) ? node15779 : node15726;
										assign node15726 = (inp[10]) ? node15750 : node15727;
											assign node15727 = (inp[11]) ? node15743 : node15728;
												assign node15728 = (inp[12]) ? node15732 : node15729;
													assign node15729 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15732 = (inp[2]) ? 4'b0001 : node15733;
														assign node15733 = (inp[5]) ? 4'b0000 : node15734;
															assign node15734 = (inp[9]) ? node15738 : node15735;
																assign node15735 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node15738 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node15743 = (inp[9]) ? 4'b0000 : node15744;
													assign node15744 = (inp[12]) ? 4'b0000 : node15745;
														assign node15745 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node15750 = (inp[9]) ? node15760 : node15751;
												assign node15751 = (inp[11]) ? node15753 : 4'b0001;
													assign node15753 = (inp[12]) ? node15757 : node15754;
														assign node15754 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node15757 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node15760 = (inp[11]) ? node15772 : node15761;
													assign node15761 = (inp[5]) ? node15767 : node15762;
														assign node15762 = (inp[12]) ? node15764 : 4'b0000;
															assign node15764 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node15767 = (inp[0]) ? 4'b0000 : node15768;
															assign node15768 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node15772 = (inp[2]) ? 4'b0001 : node15773;
														assign node15773 = (inp[0]) ? node15775 : 4'b0000;
															assign node15775 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node15779 = (inp[9]) ? 4'b0100 : 4'b0101;
							assign node15782 = (inp[1]) ? node16038 : node15783;
								assign node15783 = (inp[7]) ? node15897 : node15784;
									assign node15784 = (inp[4]) ? node15852 : node15785;
										assign node15785 = (inp[12]) ? node15829 : node15786;
											assign node15786 = (inp[0]) ? node15816 : node15787;
												assign node15787 = (inp[5]) ? node15803 : node15788;
													assign node15788 = (inp[11]) ? node15796 : node15789;
														assign node15789 = (inp[2]) ? node15793 : node15790;
															assign node15790 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node15793 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node15796 = (inp[2]) ? node15800 : node15797;
															assign node15797 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node15800 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node15803 = (inp[11]) ? node15809 : node15804;
														assign node15804 = (inp[9]) ? node15806 : 4'b0101;
															assign node15806 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node15809 = (inp[10]) ? node15811 : 4'b0101;
															assign node15811 = (inp[9]) ? 4'b0101 : node15812;
																assign node15812 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node15816 = (inp[9]) ? node15822 : node15817;
													assign node15817 = (inp[2]) ? 4'b0100 : node15818;
														assign node15818 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node15822 = (inp[5]) ? node15826 : node15823;
														assign node15823 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node15826 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node15829 = (inp[9]) ? node15841 : node15830;
												assign node15830 = (inp[2]) ? node15836 : node15831;
													assign node15831 = (inp[5]) ? 4'b0000 : node15832;
														assign node15832 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node15836 = (inp[5]) ? 4'b0001 : node15837;
														assign node15837 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node15841 = (inp[2]) ? node15847 : node15842;
													assign node15842 = (inp[0]) ? 4'b0001 : node15843;
														assign node15843 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15847 = (inp[5]) ? 4'b0000 : node15848;
														assign node15848 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node15852 = (inp[0]) ? node15882 : node15853;
											assign node15853 = (inp[5]) ? node15865 : node15854;
												assign node15854 = (inp[2]) ? node15860 : node15855;
													assign node15855 = (inp[12]) ? 4'b0010 : node15856;
														assign node15856 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node15860 = (inp[12]) ? node15862 : 4'b0010;
														assign node15862 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node15865 = (inp[2]) ? node15875 : node15866;
													assign node15866 = (inp[11]) ? node15872 : node15867;
														assign node15867 = (inp[12]) ? 4'b0010 : node15868;
															assign node15868 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node15872 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node15875 = (inp[9]) ? node15879 : node15876;
														assign node15876 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node15879 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node15882 = (inp[10]) ? node15892 : node15883;
												assign node15883 = (inp[2]) ? 4'b0011 : node15884;
													assign node15884 = (inp[9]) ? node15888 : node15885;
														assign node15885 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node15888 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node15892 = (inp[9]) ? node15894 : 4'b0010;
													assign node15894 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node15897 = (inp[4]) ? node15955 : node15898;
										assign node15898 = (inp[12]) ? node15930 : node15899;
											assign node15899 = (inp[11]) ? node15915 : node15900;
												assign node15900 = (inp[0]) ? node15908 : node15901;
													assign node15901 = (inp[2]) ? node15905 : node15902;
														assign node15902 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node15905 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node15908 = (inp[5]) ? 4'b0010 : node15909;
														assign node15909 = (inp[9]) ? node15911 : 4'b0010;
															assign node15911 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node15915 = (inp[2]) ? node15921 : node15916;
													assign node15916 = (inp[9]) ? node15918 : 4'b0011;
														assign node15918 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node15921 = (inp[9]) ? node15927 : node15922;
														assign node15922 = (inp[0]) ? node15924 : 4'b0010;
															assign node15924 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node15927 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node15930 = (inp[0]) ? node15948 : node15931;
												assign node15931 = (inp[10]) ? node15939 : node15932;
													assign node15932 = (inp[9]) ? node15934 : 4'b0110;
														assign node15934 = (inp[5]) ? 4'b0110 : node15935;
															assign node15935 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node15939 = (inp[5]) ? node15941 : 4'b0110;
														assign node15941 = (inp[2]) ? node15945 : node15942;
															assign node15942 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node15945 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node15948 = (inp[9]) ? node15952 : node15949;
													assign node15949 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node15952 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node15955 = (inp[10]) ? node16005 : node15956;
											assign node15956 = (inp[2]) ? node15988 : node15957;
												assign node15957 = (inp[11]) ? node15971 : node15958;
													assign node15958 = (inp[0]) ? node15966 : node15959;
														assign node15959 = (inp[12]) ? node15963 : node15960;
															assign node15960 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node15963 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node15966 = (inp[5]) ? node15968 : 4'b0101;
															assign node15968 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node15971 = (inp[0]) ? node15979 : node15972;
														assign node15972 = (inp[12]) ? node15976 : node15973;
															assign node15973 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node15976 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node15979 = (inp[5]) ? node15985 : node15980;
															assign node15980 = (inp[9]) ? node15982 : 4'b0100;
																assign node15982 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node15985 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node15988 = (inp[12]) ? node15996 : node15989;
													assign node15989 = (inp[0]) ? node15993 : node15990;
														assign node15990 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node15993 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node15996 = (inp[11]) ? 4'b0101 : node15997;
														assign node15997 = (inp[9]) ? node16001 : node15998;
															assign node15998 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node16001 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node16005 = (inp[5]) ? node16023 : node16006;
												assign node16006 = (inp[12]) ? node16014 : node16007;
													assign node16007 = (inp[0]) ? node16011 : node16008;
														assign node16008 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node16011 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node16014 = (inp[2]) ? node16016 : 4'b0100;
														assign node16016 = (inp[9]) ? node16020 : node16017;
															assign node16017 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node16020 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node16023 = (inp[9]) ? node16031 : node16024;
													assign node16024 = (inp[0]) ? node16028 : node16025;
														assign node16025 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node16028 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node16031 = (inp[0]) ? node16035 : node16032;
														assign node16032 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node16035 = (inp[12]) ? 4'b0100 : 4'b0101;
								assign node16038 = (inp[4]) ? node16180 : node16039;
									assign node16039 = (inp[7]) ? node16107 : node16040;
										assign node16040 = (inp[12]) ? node16062 : node16041;
											assign node16041 = (inp[9]) ? node16053 : node16042;
												assign node16042 = (inp[2]) ? node16048 : node16043;
													assign node16043 = (inp[5]) ? node16045 : 4'b0000;
														assign node16045 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node16048 = (inp[5]) ? node16050 : 4'b0001;
														assign node16050 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node16053 = (inp[2]) ? node16059 : node16054;
													assign node16054 = (inp[0]) ? node16056 : 4'b0001;
														assign node16056 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node16059 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node16062 = (inp[0]) ? node16084 : node16063;
												assign node16063 = (inp[11]) ? node16073 : node16064;
													assign node16064 = (inp[10]) ? node16066 : 4'b0101;
														assign node16066 = (inp[9]) ? node16070 : node16067;
															assign node16067 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node16070 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node16073 = (inp[5]) ? node16079 : node16074;
														assign node16074 = (inp[2]) ? 4'b0101 : node16075;
															assign node16075 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node16079 = (inp[9]) ? node16081 : 4'b0100;
															assign node16081 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node16084 = (inp[5]) ? node16092 : node16085;
													assign node16085 = (inp[2]) ? node16089 : node16086;
														assign node16086 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node16089 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node16092 = (inp[10]) ? node16100 : node16093;
														assign node16093 = (inp[11]) ? node16095 : 4'b0100;
															assign node16095 = (inp[9]) ? 4'b0100 : node16096;
																assign node16096 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node16100 = (inp[2]) ? node16104 : node16101;
															assign node16101 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node16104 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node16107 = (inp[12]) ? node16151 : node16108;
											assign node16108 = (inp[11]) ? node16134 : node16109;
												assign node16109 = (inp[10]) ? node16121 : node16110;
													assign node16110 = (inp[0]) ? node16112 : 4'b0110;
														assign node16112 = (inp[5]) ? node16118 : node16113;
															assign node16113 = (inp[2]) ? node16115 : 4'b0111;
																assign node16115 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node16118 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node16121 = (inp[0]) ? node16129 : node16122;
														assign node16122 = (inp[2]) ? 4'b0111 : node16123;
															assign node16123 = (inp[9]) ? node16125 : 4'b0111;
																assign node16125 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node16129 = (inp[9]) ? node16131 : 4'b0110;
															assign node16131 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node16134 = (inp[2]) ? node16144 : node16135;
													assign node16135 = (inp[0]) ? node16141 : node16136;
														assign node16136 = (inp[9]) ? 4'b0110 : node16137;
															assign node16137 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node16141 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node16144 = (inp[9]) ? 4'b0110 : node16145;
														assign node16145 = (inp[0]) ? 4'b0111 : node16146;
															assign node16146 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node16151 = (inp[0]) ? node16173 : node16152;
												assign node16152 = (inp[5]) ? node16164 : node16153;
													assign node16153 = (inp[10]) ? node16159 : node16154;
														assign node16154 = (inp[2]) ? 4'b0011 : node16155;
															assign node16155 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node16159 = (inp[9]) ? node16161 : 4'b0011;
															assign node16161 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node16164 = (inp[10]) ? node16170 : node16165;
														assign node16165 = (inp[2]) ? node16167 : 4'b0010;
															assign node16167 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node16170 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node16173 = (inp[2]) ? node16177 : node16174;
													assign node16174 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node16177 = (inp[9]) ? 4'b0010 : 4'b0011;
									assign node16180 = (inp[7]) ? node16204 : node16181;
										assign node16181 = (inp[9]) ? node16193 : node16182;
											assign node16182 = (inp[5]) ? node16188 : node16183;
												assign node16183 = (inp[12]) ? node16185 : 4'b0010;
													assign node16185 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node16188 = (inp[12]) ? node16190 : 4'b0011;
													assign node16190 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node16193 = (inp[5]) ? node16199 : node16194;
												assign node16194 = (inp[0]) ? 4'b0011 : node16195;
													assign node16195 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node16199 = (inp[0]) ? 4'b0010 : node16200;
													assign node16200 = (inp[12]) ? 4'b0011 : 4'b0010;
										assign node16204 = (inp[9]) ? node16208 : node16205;
											assign node16205 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node16208 = (inp[0]) ? 4'b0000 : 4'b0001;
				assign node16211 = (inp[4]) ? node17925 : node16212;
					assign node16212 = (inp[14]) ? node17012 : node16213;
						assign node16213 = (inp[15]) ? node16661 : node16214;
							assign node16214 = (inp[12]) ? node16414 : node16215;
								assign node16215 = (inp[1]) ? node16305 : node16216;
									assign node16216 = (inp[5]) ? node16238 : node16217;
										assign node16217 = (inp[11]) ? node16229 : node16218;
											assign node16218 = (inp[0]) ? node16224 : node16219;
												assign node16219 = (inp[2]) ? node16221 : 4'b0000;
													assign node16221 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node16224 = (inp[2]) ? node16226 : 4'b0001;
													assign node16226 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node16229 = (inp[0]) ? node16233 : node16230;
												assign node16230 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node16233 = (inp[13]) ? node16235 : 4'b0000;
													assign node16235 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node16238 = (inp[10]) ? node16270 : node16239;
											assign node16239 = (inp[7]) ? node16259 : node16240;
												assign node16240 = (inp[13]) ? node16252 : node16241;
													assign node16241 = (inp[2]) ? 4'b0100 : node16242;
														assign node16242 = (inp[9]) ? node16244 : 4'b0101;
															assign node16244 = (inp[0]) ? node16248 : node16245;
																assign node16245 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node16248 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node16252 = (inp[2]) ? 4'b0101 : node16253;
														assign node16253 = (inp[11]) ? 4'b0100 : node16254;
															assign node16254 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node16259 = (inp[0]) ? 4'b0101 : node16260;
													assign node16260 = (inp[11]) ? node16266 : node16261;
														assign node16261 = (inp[13]) ? node16263 : 4'b0101;
															assign node16263 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node16266 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node16270 = (inp[0]) ? node16286 : node16271;
												assign node16271 = (inp[11]) ? node16279 : node16272;
													assign node16272 = (inp[7]) ? 4'b0101 : node16273;
														assign node16273 = (inp[13]) ? node16275 : 4'b0100;
															assign node16275 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node16279 = (inp[7]) ? 4'b0100 : node16280;
														assign node16280 = (inp[13]) ? node16282 : 4'b0101;
															assign node16282 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node16286 = (inp[13]) ? node16294 : node16287;
													assign node16287 = (inp[9]) ? node16289 : 4'b0100;
														assign node16289 = (inp[7]) ? node16291 : 4'b0101;
															assign node16291 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node16294 = (inp[11]) ? node16302 : node16295;
														assign node16295 = (inp[7]) ? node16299 : node16296;
															assign node16296 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node16299 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node16302 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node16305 = (inp[5]) ? node16361 : node16306;
										assign node16306 = (inp[2]) ? node16322 : node16307;
											assign node16307 = (inp[7]) ? node16315 : node16308;
												assign node16308 = (inp[0]) ? node16312 : node16309;
													assign node16309 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node16312 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node16315 = (inp[11]) ? node16319 : node16316;
													assign node16316 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node16319 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node16322 = (inp[11]) ? node16344 : node16323;
												assign node16323 = (inp[10]) ? node16331 : node16324;
													assign node16324 = (inp[0]) ? node16328 : node16325;
														assign node16325 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node16328 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node16331 = (inp[9]) ? node16333 : 4'b0100;
														assign node16333 = (inp[7]) ? node16339 : node16334;
															assign node16334 = (inp[13]) ? 4'b0100 : node16335;
																assign node16335 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node16339 = (inp[13]) ? node16341 : 4'b0101;
																assign node16341 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node16344 = (inp[10]) ? node16350 : node16345;
													assign node16345 = (inp[13]) ? 4'b0100 : node16346;
														assign node16346 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node16350 = (inp[9]) ? node16356 : node16351;
														assign node16351 = (inp[0]) ? 4'b0100 : node16352;
															assign node16352 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node16356 = (inp[0]) ? 4'b0101 : node16357;
															assign node16357 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node16361 = (inp[0]) ? node16391 : node16362;
											assign node16362 = (inp[13]) ? node16376 : node16363;
												assign node16363 = (inp[7]) ? node16369 : node16364;
													assign node16364 = (inp[11]) ? 4'b0000 : node16365;
														assign node16365 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node16369 = (inp[2]) ? node16373 : node16370;
														assign node16370 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node16373 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node16376 = (inp[2]) ? node16384 : node16377;
													assign node16377 = (inp[7]) ? node16381 : node16378;
														assign node16378 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node16381 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16384 = (inp[11]) ? node16388 : node16385;
														assign node16385 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16388 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node16391 = (inp[2]) ? node16407 : node16392;
												assign node16392 = (inp[11]) ? node16400 : node16393;
													assign node16393 = (inp[13]) ? node16397 : node16394;
														assign node16394 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16397 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node16400 = (inp[9]) ? 4'b0001 : node16401;
														assign node16401 = (inp[7]) ? node16403 : 4'b0001;
															assign node16403 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node16407 = (inp[7]) ? node16411 : node16408;
													assign node16408 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16411 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node16414 = (inp[11]) ? node16538 : node16415;
									assign node16415 = (inp[1]) ? node16463 : node16416;
										assign node16416 = (inp[0]) ? node16438 : node16417;
											assign node16417 = (inp[13]) ? node16421 : node16418;
												assign node16418 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node16421 = (inp[2]) ? node16425 : node16422;
													assign node16422 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node16425 = (inp[10]) ? node16427 : 4'b0101;
														assign node16427 = (inp[9]) ? node16433 : node16428;
															assign node16428 = (inp[7]) ? 4'b0101 : node16429;
																assign node16429 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node16433 = (inp[5]) ? node16435 : 4'b0101;
																assign node16435 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node16438 = (inp[13]) ? node16452 : node16439;
												assign node16439 = (inp[2]) ? node16447 : node16440;
													assign node16440 = (inp[5]) ? node16444 : node16441;
														assign node16441 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node16444 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node16447 = (inp[10]) ? 4'b0001 : node16448;
														assign node16448 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node16452 = (inp[7]) ? node16460 : node16453;
													assign node16453 = (inp[5]) ? node16457 : node16454;
														assign node16454 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node16457 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node16460 = (inp[5]) ? 4'b0000 : 4'b0100;
										assign node16463 = (inp[2]) ? node16499 : node16464;
											assign node16464 = (inp[9]) ? node16482 : node16465;
												assign node16465 = (inp[5]) ? node16473 : node16466;
													assign node16466 = (inp[7]) ? node16470 : node16467;
														assign node16467 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node16470 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node16473 = (inp[7]) ? 4'b0101 : node16474;
														assign node16474 = (inp[13]) ? node16478 : node16475;
															assign node16475 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node16478 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node16482 = (inp[0]) ? node16490 : node16483;
													assign node16483 = (inp[7]) ? node16487 : node16484;
														assign node16484 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node16487 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node16490 = (inp[13]) ? 4'b0001 : node16491;
														assign node16491 = (inp[10]) ? 4'b0100 : node16492;
															assign node16492 = (inp[5]) ? node16494 : 4'b0001;
																assign node16494 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node16499 = (inp[13]) ? node16525 : node16500;
												assign node16500 = (inp[0]) ? node16510 : node16501;
													assign node16501 = (inp[9]) ? 4'b0101 : node16502;
														assign node16502 = (inp[10]) ? 4'b0101 : node16503;
															assign node16503 = (inp[5]) ? node16505 : 4'b0000;
																assign node16505 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node16510 = (inp[10]) ? 4'b0100 : node16511;
														assign node16511 = (inp[9]) ? node16517 : node16512;
															assign node16512 = (inp[7]) ? 4'b0100 : node16513;
																assign node16513 = (inp[5]) ? 4'b0001 : 4'b0100;
															assign node16517 = (inp[5]) ? node16521 : node16518;
																assign node16518 = (inp[7]) ? 4'b0001 : 4'b0100;
																assign node16521 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node16525 = (inp[0]) ? node16533 : node16526;
													assign node16526 = (inp[5]) ? node16530 : node16527;
														assign node16527 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node16530 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node16533 = (inp[5]) ? node16535 : 4'b0101;
														assign node16535 = (inp[7]) ? 4'b0101 : 4'b0001;
									assign node16538 = (inp[0]) ? node16612 : node16539;
										assign node16539 = (inp[7]) ? node16589 : node16540;
											assign node16540 = (inp[9]) ? node16566 : node16541;
												assign node16541 = (inp[10]) ? node16553 : node16542;
													assign node16542 = (inp[5]) ? node16548 : node16543;
														assign node16543 = (inp[1]) ? 4'b0101 : node16544;
															assign node16544 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node16548 = (inp[2]) ? 4'b0001 : node16549;
															assign node16549 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node16553 = (inp[1]) ? node16559 : node16554;
														assign node16554 = (inp[5]) ? 4'b0101 : node16555;
															assign node16555 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node16559 = (inp[5]) ? node16561 : 4'b0101;
															assign node16561 = (inp[13]) ? 4'b0001 : node16562;
																assign node16562 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node16566 = (inp[10]) ? node16576 : node16567;
													assign node16567 = (inp[13]) ? node16571 : node16568;
														assign node16568 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node16571 = (inp[1]) ? node16573 : 4'b0000;
															assign node16573 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node16576 = (inp[13]) ? node16582 : node16577;
														assign node16577 = (inp[1]) ? node16579 : 4'b0001;
															assign node16579 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node16582 = (inp[2]) ? node16584 : 4'b0100;
															assign node16584 = (inp[1]) ? 4'b0001 : node16585;
																assign node16585 = (inp[5]) ? 4'b0100 : 4'b0000;
											assign node16589 = (inp[2]) ? node16599 : node16590;
												assign node16590 = (inp[1]) ? node16596 : node16591;
													assign node16591 = (inp[5]) ? 4'b0001 : node16592;
														assign node16592 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node16596 = (inp[5]) ? 4'b0100 : 4'b0001;
												assign node16599 = (inp[5]) ? node16605 : node16600;
													assign node16600 = (inp[1]) ? node16602 : 4'b0100;
														assign node16602 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node16605 = (inp[1]) ? node16609 : node16606;
														assign node16606 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node16609 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node16612 = (inp[2]) ? node16632 : node16613;
											assign node16613 = (inp[1]) ? node16623 : node16614;
												assign node16614 = (inp[5]) ? node16620 : node16615;
													assign node16615 = (inp[7]) ? node16617 : 4'b0000;
														assign node16617 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node16620 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node16623 = (inp[5]) ? node16627 : node16624;
													assign node16624 = (inp[7]) ? 4'b0000 : 4'b0101;
													assign node16627 = (inp[7]) ? 4'b0101 : node16628;
														assign node16628 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node16632 = (inp[7]) ? node16648 : node16633;
												assign node16633 = (inp[13]) ? node16641 : node16634;
													assign node16634 = (inp[5]) ? node16638 : node16635;
														assign node16635 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node16638 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node16641 = (inp[1]) ? node16645 : node16642;
														assign node16642 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node16645 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node16648 = (inp[5]) ? node16654 : node16649;
													assign node16649 = (inp[1]) ? node16651 : 4'b0101;
														assign node16651 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node16654 = (inp[1]) ? node16658 : node16655;
														assign node16655 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node16658 = (inp[13]) ? 4'b0100 : 4'b0101;
							assign node16661 = (inp[0]) ? node16845 : node16662;
								assign node16662 = (inp[11]) ? node16738 : node16663;
									assign node16663 = (inp[13]) ? node16695 : node16664;
										assign node16664 = (inp[1]) ? node16678 : node16665;
											assign node16665 = (inp[5]) ? node16671 : node16666;
												assign node16666 = (inp[7]) ? node16668 : 4'b0010;
													assign node16668 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node16671 = (inp[12]) ? 4'b0110 : node16672;
													assign node16672 = (inp[7]) ? node16674 : 4'b0110;
														assign node16674 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node16678 = (inp[5]) ? node16690 : node16679;
												assign node16679 = (inp[12]) ? node16685 : node16680;
													assign node16680 = (inp[7]) ? 4'b0011 : node16681;
														assign node16681 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node16685 = (inp[2]) ? node16687 : 4'b0110;
														assign node16687 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node16690 = (inp[12]) ? 4'b0010 : node16691;
													assign node16691 = (inp[7]) ? 4'b0110 : 4'b0011;
										assign node16695 = (inp[2]) ? node16715 : node16696;
											assign node16696 = (inp[5]) ? node16706 : node16697;
												assign node16697 = (inp[1]) ? node16703 : node16698;
													assign node16698 = (inp[7]) ? node16700 : 4'b0011;
														assign node16700 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node16703 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node16706 = (inp[1]) ? node16712 : node16707;
													assign node16707 = (inp[12]) ? 4'b0111 : node16708;
														assign node16708 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node16712 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node16715 = (inp[1]) ? node16727 : node16716;
												assign node16716 = (inp[5]) ? node16722 : node16717;
													assign node16717 = (inp[7]) ? node16719 : 4'b0010;
														assign node16719 = (inp[12]) ? 4'b0011 : 4'b0110;
													assign node16722 = (inp[12]) ? 4'b0110 : node16723;
														assign node16723 = (inp[7]) ? 4'b0011 : 4'b0110;
												assign node16727 = (inp[5]) ? node16733 : node16728;
													assign node16728 = (inp[12]) ? node16730 : 4'b0110;
														assign node16730 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node16733 = (inp[7]) ? node16735 : 4'b0011;
														assign node16735 = (inp[12]) ? 4'b0010 : 4'b0110;
									assign node16738 = (inp[13]) ? node16776 : node16739;
										assign node16739 = (inp[12]) ? node16765 : node16740;
											assign node16740 = (inp[1]) ? node16750 : node16741;
												assign node16741 = (inp[5]) ? node16745 : node16742;
													assign node16742 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node16745 = (inp[7]) ? node16747 : 4'b0111;
														assign node16747 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node16750 = (inp[2]) ? node16758 : node16751;
													assign node16751 = (inp[5]) ? node16755 : node16752;
														assign node16752 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node16755 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node16758 = (inp[5]) ? node16762 : node16759;
														assign node16759 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node16762 = (inp[7]) ? 4'b0111 : 4'b0010;
											assign node16765 = (inp[5]) ? node16773 : node16766;
												assign node16766 = (inp[1]) ? node16770 : node16767;
													assign node16767 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node16770 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node16773 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node16776 = (inp[2]) ? node16800 : node16777;
											assign node16777 = (inp[5]) ? node16789 : node16778;
												assign node16778 = (inp[1]) ? node16784 : node16779;
													assign node16779 = (inp[12]) ? 4'b0011 : node16780;
														assign node16780 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node16784 = (inp[7]) ? 4'b0111 : node16785;
														assign node16785 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node16789 = (inp[1]) ? node16795 : node16790;
													assign node16790 = (inp[7]) ? node16792 : 4'b0110;
														assign node16792 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node16795 = (inp[12]) ? 4'b0010 : node16796;
														assign node16796 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node16800 = (inp[10]) ? node16826 : node16801;
												assign node16801 = (inp[5]) ? node16817 : node16802;
													assign node16802 = (inp[1]) ? node16810 : node16803;
														assign node16803 = (inp[12]) ? node16807 : node16804;
															assign node16804 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node16807 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node16810 = (inp[12]) ? node16814 : node16811;
															assign node16811 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node16814 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node16817 = (inp[12]) ? 4'b0011 : node16818;
														assign node16818 = (inp[7]) ? node16822 : node16819;
															assign node16819 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node16822 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node16826 = (inp[12]) ? node16840 : node16827;
													assign node16827 = (inp[7]) ? node16833 : node16828;
														assign node16828 = (inp[5]) ? 4'b0111 : node16829;
															assign node16829 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node16833 = (inp[5]) ? node16837 : node16834;
															assign node16834 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node16837 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node16840 = (inp[7]) ? 4'b0111 : node16841;
														assign node16841 = (inp[5]) ? 4'b0111 : 4'b0110;
								assign node16845 = (inp[11]) ? node16931 : node16846;
									assign node16846 = (inp[13]) ? node16878 : node16847;
										assign node16847 = (inp[5]) ? node16865 : node16848;
											assign node16848 = (inp[1]) ? node16854 : node16849;
												assign node16849 = (inp[7]) ? node16851 : 4'b0011;
													assign node16851 = (inp[12]) ? 4'b0010 : 4'b0111;
												assign node16854 = (inp[12]) ? node16858 : node16855;
													assign node16855 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node16858 = (inp[10]) ? node16860 : 4'b0110;
														assign node16860 = (inp[9]) ? 4'b0111 : node16861;
															assign node16861 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node16865 = (inp[1]) ? node16873 : node16866;
												assign node16866 = (inp[7]) ? node16868 : 4'b0111;
													assign node16868 = (inp[12]) ? 4'b0111 : node16869;
														assign node16869 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node16873 = (inp[12]) ? 4'b0011 : node16874;
													assign node16874 = (inp[7]) ? 4'b0111 : 4'b0010;
										assign node16878 = (inp[2]) ? node16906 : node16879;
											assign node16879 = (inp[5]) ? node16895 : node16880;
												assign node16880 = (inp[1]) ? node16888 : node16881;
													assign node16881 = (inp[12]) ? node16885 : node16882;
														assign node16882 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node16885 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node16888 = (inp[12]) ? node16892 : node16889;
														assign node16889 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node16892 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node16895 = (inp[1]) ? node16901 : node16896;
													assign node16896 = (inp[12]) ? 4'b0110 : node16897;
														assign node16897 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node16901 = (inp[12]) ? 4'b0010 : node16902;
														assign node16902 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node16906 = (inp[1]) ? node16918 : node16907;
												assign node16907 = (inp[5]) ? node16913 : node16908;
													assign node16908 = (inp[7]) ? node16910 : 4'b0011;
														assign node16910 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node16913 = (inp[12]) ? 4'b0111 : node16914;
														assign node16914 = (inp[7]) ? 4'b0010 : 4'b0111;
												assign node16918 = (inp[5]) ? node16926 : node16919;
													assign node16919 = (inp[7]) ? node16923 : node16920;
														assign node16920 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node16923 = (inp[12]) ? 4'b0111 : 4'b0010;
													assign node16926 = (inp[12]) ? 4'b0011 : node16927;
														assign node16927 = (inp[7]) ? 4'b0111 : 4'b0010;
									assign node16931 = (inp[1]) ? node16969 : node16932;
										assign node16932 = (inp[5]) ? node16950 : node16933;
											assign node16933 = (inp[7]) ? node16939 : node16934;
												assign node16934 = (inp[13]) ? node16936 : 4'b0010;
													assign node16936 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node16939 = (inp[12]) ? node16945 : node16940;
													assign node16940 = (inp[13]) ? node16942 : 4'b0110;
														assign node16942 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node16945 = (inp[13]) ? node16947 : 4'b0011;
														assign node16947 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node16950 = (inp[13]) ? node16958 : node16951;
												assign node16951 = (inp[7]) ? node16953 : 4'b0110;
													assign node16953 = (inp[12]) ? 4'b0110 : node16954;
														assign node16954 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node16958 = (inp[2]) ? node16964 : node16959;
													assign node16959 = (inp[12]) ? 4'b0111 : node16960;
														assign node16960 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node16964 = (inp[7]) ? node16966 : 4'b0110;
														assign node16966 = (inp[12]) ? 4'b0110 : 4'b0011;
										assign node16969 = (inp[5]) ? node16991 : node16970;
											assign node16970 = (inp[7]) ? node16982 : node16971;
												assign node16971 = (inp[12]) ? node16977 : node16972;
													assign node16972 = (inp[13]) ? 4'b0110 : node16973;
														assign node16973 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node16977 = (inp[13]) ? 4'b0111 : node16978;
														assign node16978 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node16982 = (inp[12]) ? node16988 : node16983;
													assign node16983 = (inp[2]) ? 4'b0011 : node16984;
														assign node16984 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node16988 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node16991 = (inp[7]) ? node17003 : node16992;
												assign node16992 = (inp[12]) ? node16998 : node16993;
													assign node16993 = (inp[13]) ? node16995 : 4'b0011;
														assign node16995 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node16998 = (inp[2]) ? 4'b0010 : node16999;
														assign node16999 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node17003 = (inp[12]) ? node17009 : node17004;
													assign node17004 = (inp[2]) ? 4'b0110 : node17005;
														assign node17005 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node17009 = (inp[2]) ? 4'b0010 : 4'b0011;
						assign node17012 = (inp[10]) ? node17438 : node17013;
							assign node17013 = (inp[5]) ? node17199 : node17014;
								assign node17014 = (inp[2]) ? node17100 : node17015;
									assign node17015 = (inp[0]) ? node17061 : node17016;
										assign node17016 = (inp[12]) ? node17032 : node17017;
											assign node17017 = (inp[1]) ? node17025 : node17018;
												assign node17018 = (inp[13]) ? node17020 : 4'b0010;
													assign node17020 = (inp[7]) ? 4'b0010 : node17021;
														assign node17021 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node17025 = (inp[15]) ? node17027 : 4'b0110;
													assign node17027 = (inp[7]) ? node17029 : 4'b0110;
														assign node17029 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node17032 = (inp[1]) ? node17046 : node17033;
												assign node17033 = (inp[13]) ? node17039 : node17034;
													assign node17034 = (inp[7]) ? node17036 : 4'b0110;
														assign node17036 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node17039 = (inp[15]) ? node17043 : node17040;
														assign node17040 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17043 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node17046 = (inp[15]) ? node17052 : node17047;
													assign node17047 = (inp[13]) ? 4'b0010 : node17048;
														assign node17048 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17052 = (inp[9]) ? node17054 : 4'b0011;
														assign node17054 = (inp[11]) ? 4'b0011 : node17055;
															assign node17055 = (inp[7]) ? node17057 : 4'b0010;
																assign node17057 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node17061 = (inp[12]) ? node17077 : node17062;
											assign node17062 = (inp[1]) ? node17070 : node17063;
												assign node17063 = (inp[13]) ? node17065 : 4'b0011;
													assign node17065 = (inp[9]) ? 4'b0011 : node17066;
														assign node17066 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node17070 = (inp[13]) ? 4'b0111 : node17071;
													assign node17071 = (inp[7]) ? node17073 : 4'b0111;
														assign node17073 = (inp[15]) ? 4'b0110 : 4'b0111;
											assign node17077 = (inp[1]) ? node17089 : node17078;
												assign node17078 = (inp[13]) ? node17084 : node17079;
													assign node17079 = (inp[7]) ? node17081 : 4'b0111;
														assign node17081 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node17084 = (inp[15]) ? node17086 : 4'b0110;
														assign node17086 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node17089 = (inp[15]) ? node17093 : node17090;
													assign node17090 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node17093 = (inp[13]) ? node17097 : node17094;
														assign node17094 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17097 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node17100 = (inp[0]) ? node17146 : node17101;
										assign node17101 = (inp[15]) ? node17117 : node17102;
											assign node17102 = (inp[12]) ? node17106 : node17103;
												assign node17103 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node17106 = (inp[1]) ? node17112 : node17107;
													assign node17107 = (inp[7]) ? node17109 : 4'b0111;
														assign node17109 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node17112 = (inp[13]) ? 4'b0011 : node17113;
														assign node17113 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node17117 = (inp[13]) ? node17135 : node17118;
												assign node17118 = (inp[7]) ? node17124 : node17119;
													assign node17119 = (inp[12]) ? node17121 : 4'b0011;
														assign node17121 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node17124 = (inp[11]) ? node17130 : node17125;
														assign node17125 = (inp[12]) ? 4'b0110 : node17126;
															assign node17126 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node17130 = (inp[12]) ? node17132 : 4'b0110;
															assign node17132 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node17135 = (inp[7]) ? node17143 : node17136;
													assign node17136 = (inp[1]) ? node17140 : node17137;
														assign node17137 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node17140 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node17143 = (inp[11]) ? 4'b0111 : 4'b0011;
										assign node17146 = (inp[12]) ? node17164 : node17147;
											assign node17147 = (inp[1]) ? node17157 : node17148;
												assign node17148 = (inp[13]) ? node17150 : 4'b0010;
													assign node17150 = (inp[11]) ? node17152 : 4'b0010;
														assign node17152 = (inp[15]) ? node17154 : 4'b0010;
															assign node17154 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node17157 = (inp[15]) ? node17159 : 4'b0110;
													assign node17159 = (inp[7]) ? node17161 : 4'b0110;
														assign node17161 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node17164 = (inp[1]) ? node17186 : node17165;
												assign node17165 = (inp[15]) ? node17171 : node17166;
													assign node17166 = (inp[7]) ? node17168 : 4'b0110;
														assign node17168 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node17171 = (inp[9]) ? node17179 : node17172;
														assign node17172 = (inp[13]) ? node17176 : node17173;
															assign node17173 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node17176 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node17179 = (inp[7]) ? node17183 : node17180;
															assign node17180 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node17183 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node17186 = (inp[15]) ? node17192 : node17187;
													assign node17187 = (inp[11]) ? node17189 : 4'b0010;
														assign node17189 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node17192 = (inp[7]) ? node17196 : node17193;
														assign node17193 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node17196 = (inp[13]) ? 4'b0010 : 4'b0011;
								assign node17199 = (inp[2]) ? node17325 : node17200;
									assign node17200 = (inp[0]) ? node17250 : node17201;
										assign node17201 = (inp[12]) ? node17239 : node17202;
											assign node17202 = (inp[1]) ? node17220 : node17203;
												assign node17203 = (inp[11]) ? node17213 : node17204;
													assign node17204 = (inp[7]) ? node17208 : node17205;
														assign node17205 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node17208 = (inp[13]) ? node17210 : 4'b0011;
															assign node17210 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node17213 = (inp[15]) ? 4'b0010 : node17214;
														assign node17214 = (inp[7]) ? node17216 : 4'b0010;
															assign node17216 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node17220 = (inp[15]) ? node17234 : node17221;
													assign node17221 = (inp[11]) ? node17229 : node17222;
														assign node17222 = (inp[13]) ? node17226 : node17223;
															assign node17223 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node17226 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node17229 = (inp[13]) ? 4'b0111 : node17230;
															assign node17230 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node17234 = (inp[7]) ? 4'b0110 : node17235;
														assign node17235 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node17239 = (inp[1]) ? 4'b0010 : node17240;
												assign node17240 = (inp[11]) ? 4'b0110 : node17241;
													assign node17241 = (inp[13]) ? node17243 : 4'b0110;
														assign node17243 = (inp[7]) ? 4'b0110 : node17244;
															assign node17244 = (inp[15]) ? 4'b0110 : 4'b0111;
										assign node17250 = (inp[15]) ? node17302 : node17251;
											assign node17251 = (inp[13]) ? node17281 : node17252;
												assign node17252 = (inp[7]) ? node17276 : node17253;
													assign node17253 = (inp[11]) ? node17263 : node17254;
														assign node17254 = (inp[9]) ? 4'b0111 : node17255;
															assign node17255 = (inp[1]) ? node17259 : node17256;
																assign node17256 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node17259 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node17263 = (inp[9]) ? node17271 : node17264;
															assign node17264 = (inp[1]) ? node17268 : node17265;
																assign node17265 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node17268 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node17271 = (inp[12]) ? 4'b0011 : node17272;
																assign node17272 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node17276 = (inp[12]) ? node17278 : 4'b0110;
														assign node17278 = (inp[1]) ? 4'b0010 : 4'b0111;
												assign node17281 = (inp[7]) ? node17293 : node17282;
													assign node17282 = (inp[11]) ? node17288 : node17283;
														assign node17283 = (inp[1]) ? 4'b0110 : node17284;
															assign node17284 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node17288 = (inp[1]) ? 4'b0011 : node17289;
															assign node17289 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node17293 = (inp[9]) ? node17295 : 4'b0011;
														assign node17295 = (inp[11]) ? 4'b0111 : node17296;
															assign node17296 = (inp[1]) ? 4'b0011 : node17297;
																assign node17297 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node17302 = (inp[9]) ? node17318 : node17303;
												assign node17303 = (inp[1]) ? node17311 : node17304;
													assign node17304 = (inp[12]) ? 4'b0111 : node17305;
														assign node17305 = (inp[7]) ? node17307 : 4'b0011;
															assign node17307 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node17311 = (inp[12]) ? 4'b0011 : node17312;
														assign node17312 = (inp[13]) ? 4'b0111 : node17313;
															assign node17313 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node17318 = (inp[1]) ? node17322 : node17319;
													assign node17319 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node17322 = (inp[12]) ? 4'b0011 : 4'b0111;
									assign node17325 = (inp[0]) ? node17389 : node17326;
										assign node17326 = (inp[15]) ? node17374 : node17327;
											assign node17327 = (inp[9]) ? node17353 : node17328;
												assign node17328 = (inp[1]) ? node17340 : node17329;
													assign node17329 = (inp[12]) ? node17335 : node17330;
														assign node17330 = (inp[13]) ? node17332 : 4'b0011;
															assign node17332 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17335 = (inp[13]) ? node17337 : 4'b0111;
															assign node17337 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node17340 = (inp[12]) ? node17348 : node17341;
														assign node17341 = (inp[11]) ? 4'b0111 : node17342;
															assign node17342 = (inp[13]) ? node17344 : 4'b0110;
																assign node17344 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17348 = (inp[13]) ? 4'b0011 : node17349;
															assign node17349 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node17353 = (inp[11]) ? node17365 : node17354;
													assign node17354 = (inp[12]) ? node17362 : node17355;
														assign node17355 = (inp[1]) ? node17357 : 4'b0010;
															assign node17357 = (inp[13]) ? node17359 : 4'b0110;
																assign node17359 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17362 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node17365 = (inp[1]) ? node17371 : node17366;
														assign node17366 = (inp[13]) ? node17368 : 4'b0111;
															assign node17368 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17371 = (inp[12]) ? 4'b0010 : 4'b0111;
											assign node17374 = (inp[12]) ? node17386 : node17375;
												assign node17375 = (inp[1]) ? node17381 : node17376;
													assign node17376 = (inp[7]) ? node17378 : 4'b0011;
														assign node17378 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node17381 = (inp[13]) ? 4'b0111 : node17382;
														assign node17382 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node17386 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node17389 = (inp[15]) ? node17423 : node17390;
											assign node17390 = (inp[12]) ? node17412 : node17391;
												assign node17391 = (inp[1]) ? node17405 : node17392;
													assign node17392 = (inp[9]) ? node17398 : node17393;
														assign node17393 = (inp[7]) ? 4'b0011 : node17394;
															assign node17394 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node17398 = (inp[13]) ? node17402 : node17399;
															assign node17399 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17402 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17405 = (inp[7]) ? node17409 : node17406;
														assign node17406 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node17409 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node17412 = (inp[1]) ? node17418 : node17413;
													assign node17413 = (inp[13]) ? node17415 : 4'b0110;
														assign node17415 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node17418 = (inp[7]) ? node17420 : 4'b0010;
														assign node17420 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node17423 = (inp[12]) ? node17435 : node17424;
												assign node17424 = (inp[1]) ? node17430 : node17425;
													assign node17425 = (inp[13]) ? node17427 : 4'b0010;
														assign node17427 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node17430 = (inp[13]) ? 4'b0110 : node17431;
														assign node17431 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node17435 = (inp[1]) ? 4'b0010 : 4'b0110;
							assign node17438 = (inp[1]) ? node17700 : node17439;
								assign node17439 = (inp[12]) ? node17589 : node17440;
									assign node17440 = (inp[13]) ? node17496 : node17441;
										assign node17441 = (inp[7]) ? node17463 : node17442;
											assign node17442 = (inp[5]) ? node17450 : node17443;
												assign node17443 = (inp[0]) ? node17447 : node17444;
													assign node17444 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17447 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node17450 = (inp[9]) ? node17458 : node17451;
													assign node17451 = (inp[0]) ? node17455 : node17452;
														assign node17452 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node17455 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node17458 = (inp[0]) ? 4'b0011 : node17459;
														assign node17459 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node17463 = (inp[15]) ? node17473 : node17464;
												assign node17464 = (inp[0]) ? 4'b0011 : node17465;
													assign node17465 = (inp[2]) ? node17469 : node17466;
														assign node17466 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node17469 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node17473 = (inp[11]) ? node17489 : node17474;
													assign node17474 = (inp[9]) ? node17482 : node17475;
														assign node17475 = (inp[2]) ? node17479 : node17476;
															assign node17476 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node17479 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node17482 = (inp[5]) ? node17484 : 4'b0010;
															assign node17484 = (inp[2]) ? 4'b0011 : node17485;
																assign node17485 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node17489 = (inp[2]) ? node17493 : node17490;
														assign node17490 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node17493 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node17496 = (inp[5]) ? node17546 : node17497;
											assign node17497 = (inp[9]) ? node17515 : node17498;
												assign node17498 = (inp[0]) ? node17506 : node17499;
													assign node17499 = (inp[2]) ? node17501 : 4'b0010;
														assign node17501 = (inp[15]) ? node17503 : 4'b0011;
															assign node17503 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node17506 = (inp[7]) ? node17512 : node17507;
														assign node17507 = (inp[2]) ? 4'b0011 : node17508;
															assign node17508 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node17512 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node17515 = (inp[11]) ? node17531 : node17516;
													assign node17516 = (inp[0]) ? node17526 : node17517;
														assign node17517 = (inp[15]) ? node17521 : node17518;
															assign node17518 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node17521 = (inp[7]) ? 4'b0010 : node17522;
																assign node17522 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node17526 = (inp[2]) ? 4'b0010 : node17527;
															assign node17527 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node17531 = (inp[15]) ? node17539 : node17532;
														assign node17532 = (inp[7]) ? node17534 : 4'b0011;
															assign node17534 = (inp[0]) ? node17536 : 4'b0010;
																assign node17536 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node17539 = (inp[2]) ? node17541 : 4'b0011;
															assign node17541 = (inp[7]) ? 4'b0011 : node17542;
																assign node17542 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node17546 = (inp[11]) ? node17574 : node17547;
												assign node17547 = (inp[9]) ? node17563 : node17548;
													assign node17548 = (inp[7]) ? node17554 : node17549;
														assign node17549 = (inp[15]) ? 4'b0010 : node17550;
															assign node17550 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node17554 = (inp[0]) ? 4'b0011 : node17555;
															assign node17555 = (inp[15]) ? node17559 : node17556;
																assign node17556 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node17559 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node17563 = (inp[2]) ? node17567 : node17564;
														assign node17564 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17567 = (inp[7]) ? node17569 : 4'b0010;
															assign node17569 = (inp[15]) ? 4'b0010 : node17570;
																assign node17570 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node17574 = (inp[15]) ? 4'b0010 : node17575;
													assign node17575 = (inp[2]) ? node17583 : node17576;
														assign node17576 = (inp[0]) ? node17580 : node17577;
															assign node17577 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node17580 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17583 = (inp[7]) ? 4'b0010 : node17584;
															assign node17584 = (inp[0]) ? 4'b0011 : 4'b0010;
									assign node17589 = (inp[7]) ? node17633 : node17590;
										assign node17590 = (inp[2]) ? node17614 : node17591;
											assign node17591 = (inp[0]) ? node17603 : node17592;
												assign node17592 = (inp[13]) ? node17594 : 4'b0110;
													assign node17594 = (inp[9]) ? node17600 : node17595;
														assign node17595 = (inp[15]) ? node17597 : 4'b0111;
															assign node17597 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node17600 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node17603 = (inp[13]) ? node17605 : 4'b0111;
													assign node17605 = (inp[11]) ? node17611 : node17606;
														assign node17606 = (inp[15]) ? 4'b0111 : node17607;
															assign node17607 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node17611 = (inp[15]) ? 4'b0110 : 4'b0111;
											assign node17614 = (inp[0]) ? node17626 : node17615;
												assign node17615 = (inp[13]) ? node17617 : 4'b0111;
													assign node17617 = (inp[11]) ? node17623 : node17618;
														assign node17618 = (inp[15]) ? 4'b0110 : node17619;
															assign node17619 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node17623 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node17626 = (inp[13]) ? node17628 : 4'b0110;
													assign node17628 = (inp[5]) ? 4'b0111 : node17629;
														assign node17629 = (inp[15]) ? 4'b0111 : 4'b0110;
										assign node17633 = (inp[9]) ? node17671 : node17634;
											assign node17634 = (inp[15]) ? node17652 : node17635;
												assign node17635 = (inp[0]) ? node17647 : node17636;
													assign node17636 = (inp[2]) ? node17642 : node17637;
														assign node17637 = (inp[5]) ? 4'b0110 : node17638;
															assign node17638 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node17642 = (inp[5]) ? 4'b0111 : node17643;
															assign node17643 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node17647 = (inp[2]) ? 4'b0110 : node17648;
														assign node17648 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node17652 = (inp[0]) ? node17660 : node17653;
													assign node17653 = (inp[2]) ? node17655 : 4'b0110;
														assign node17655 = (inp[11]) ? node17657 : 4'b0111;
															assign node17657 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node17660 = (inp[2]) ? node17666 : node17661;
														assign node17661 = (inp[5]) ? 4'b0111 : node17662;
															assign node17662 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node17666 = (inp[13]) ? 4'b0110 : node17667;
															assign node17667 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node17671 = (inp[0]) ? node17685 : node17672;
												assign node17672 = (inp[2]) ? node17680 : node17673;
													assign node17673 = (inp[15]) ? node17675 : 4'b0110;
														assign node17675 = (inp[5]) ? 4'b0110 : node17676;
															assign node17676 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node17680 = (inp[5]) ? 4'b0111 : node17681;
														assign node17681 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node17685 = (inp[2]) ? node17693 : node17686;
													assign node17686 = (inp[13]) ? 4'b0111 : node17687;
														assign node17687 = (inp[15]) ? node17689 : 4'b0111;
															assign node17689 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node17693 = (inp[5]) ? 4'b0110 : node17694;
														assign node17694 = (inp[13]) ? node17696 : 4'b0110;
															assign node17696 = (inp[15]) ? 4'b0110 : 4'b0111;
								assign node17700 = (inp[12]) ? node17826 : node17701;
									assign node17701 = (inp[5]) ? node17731 : node17702;
										assign node17702 = (inp[7]) ? node17718 : node17703;
											assign node17703 = (inp[11]) ? node17711 : node17704;
												assign node17704 = (inp[0]) ? node17708 : node17705;
													assign node17705 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node17708 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node17711 = (inp[0]) ? node17715 : node17712;
													assign node17712 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node17715 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node17718 = (inp[2]) ? node17724 : node17719;
												assign node17719 = (inp[0]) ? 4'b0111 : node17720;
													assign node17720 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node17724 = (inp[0]) ? node17726 : 4'b0111;
													assign node17726 = (inp[15]) ? node17728 : 4'b0110;
														assign node17728 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node17731 = (inp[15]) ? node17771 : node17732;
											assign node17732 = (inp[9]) ? node17754 : node17733;
												assign node17733 = (inp[13]) ? node17743 : node17734;
													assign node17734 = (inp[0]) ? 4'b0111 : node17735;
														assign node17735 = (inp[7]) ? node17739 : node17736;
															assign node17736 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node17739 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node17743 = (inp[7]) ? node17751 : node17744;
														assign node17744 = (inp[2]) ? node17748 : node17745;
															assign node17745 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node17748 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node17751 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node17754 = (inp[7]) ? node17756 : 4'b0110;
													assign node17756 = (inp[2]) ? node17766 : node17757;
														assign node17757 = (inp[11]) ? 4'b0111 : node17758;
															assign node17758 = (inp[13]) ? node17762 : node17759;
																assign node17759 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node17762 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node17766 = (inp[0]) ? node17768 : 4'b0110;
															assign node17768 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node17771 = (inp[13]) ? node17803 : node17772;
												assign node17772 = (inp[9]) ? node17786 : node17773;
													assign node17773 = (inp[7]) ? node17775 : 4'b0110;
														assign node17775 = (inp[11]) ? node17781 : node17776;
															assign node17776 = (inp[0]) ? node17778 : 4'b0110;
																assign node17778 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node17781 = (inp[2]) ? node17783 : 4'b0110;
																assign node17783 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node17786 = (inp[7]) ? node17798 : node17787;
														assign node17787 = (inp[11]) ? node17793 : node17788;
															assign node17788 = (inp[2]) ? node17790 : 4'b0111;
																assign node17790 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node17793 = (inp[0]) ? node17795 : 4'b0111;
																assign node17795 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node17798 = (inp[0]) ? 4'b0110 : node17799;
															assign node17799 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node17803 = (inp[11]) ? node17809 : node17804;
													assign node17804 = (inp[2]) ? node17806 : 4'b0111;
														assign node17806 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node17809 = (inp[7]) ? node17819 : node17810;
														assign node17810 = (inp[9]) ? 4'b0111 : node17811;
															assign node17811 = (inp[0]) ? node17815 : node17812;
																assign node17812 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node17815 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node17819 = (inp[0]) ? node17823 : node17820;
															assign node17820 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node17823 = (inp[2]) ? 4'b0110 : 4'b0111;
									assign node17826 = (inp[15]) ? node17866 : node17827;
										assign node17827 = (inp[2]) ? node17841 : node17828;
											assign node17828 = (inp[0]) ? 4'b0011 : node17829;
												assign node17829 = (inp[13]) ? 4'b0010 : node17830;
													assign node17830 = (inp[11]) ? node17832 : 4'b0011;
														assign node17832 = (inp[7]) ? node17836 : node17833;
															assign node17833 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node17836 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node17841 = (inp[0]) ? node17851 : node17842;
												assign node17842 = (inp[13]) ? 4'b0011 : node17843;
													assign node17843 = (inp[7]) ? node17847 : node17844;
														assign node17844 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node17847 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node17851 = (inp[13]) ? 4'b0010 : node17852;
													assign node17852 = (inp[11]) ? node17860 : node17853;
														assign node17853 = (inp[5]) ? node17857 : node17854;
															assign node17854 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node17857 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17860 = (inp[9]) ? 4'b0011 : node17861;
															assign node17861 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node17866 = (inp[9]) ? node17902 : node17867;
											assign node17867 = (inp[0]) ? node17885 : node17868;
												assign node17868 = (inp[2]) ? node17880 : node17869;
													assign node17869 = (inp[5]) ? 4'b0010 : node17870;
														assign node17870 = (inp[11]) ? 4'b0011 : node17871;
															assign node17871 = (inp[13]) ? node17875 : node17872;
																assign node17872 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node17875 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17880 = (inp[13]) ? 4'b0011 : node17881;
														assign node17881 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node17885 = (inp[2]) ? node17893 : node17886;
													assign node17886 = (inp[5]) ? 4'b0011 : node17887;
														assign node17887 = (inp[13]) ? 4'b0010 : node17888;
															assign node17888 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17893 = (inp[5]) ? 4'b0010 : node17894;
														assign node17894 = (inp[7]) ? node17898 : node17895;
															assign node17895 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node17898 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node17902 = (inp[2]) ? node17918 : node17903;
												assign node17903 = (inp[0]) ? node17911 : node17904;
													assign node17904 = (inp[5]) ? 4'b0010 : node17905;
														assign node17905 = (inp[13]) ? node17907 : 4'b0010;
															assign node17907 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17911 = (inp[5]) ? 4'b0011 : node17912;
														assign node17912 = (inp[13]) ? node17914 : 4'b0010;
															assign node17914 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node17918 = (inp[0]) ? node17920 : 4'b0011;
													assign node17920 = (inp[13]) ? node17922 : 4'b0010;
														assign node17922 = (inp[7]) ? 4'b0010 : 4'b0011;
					assign node17925 = (inp[14]) ? node19181 : node17926;
						assign node17926 = (inp[15]) ? node18572 : node17927;
							assign node17927 = (inp[10]) ? node18239 : node17928;
								assign node17928 = (inp[5]) ? node18074 : node17929;
									assign node17929 = (inp[1]) ? node18009 : node17930;
										assign node17930 = (inp[7]) ? node17974 : node17931;
											assign node17931 = (inp[12]) ? node17955 : node17932;
												assign node17932 = (inp[9]) ? node17944 : node17933;
													assign node17933 = (inp[2]) ? node17939 : node17934;
														assign node17934 = (inp[11]) ? node17936 : 4'b0011;
															assign node17936 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node17939 = (inp[13]) ? node17941 : 4'b0010;
															assign node17941 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node17944 = (inp[11]) ? node17946 : 4'b0010;
														assign node17946 = (inp[13]) ? node17952 : node17947;
															assign node17947 = (inp[0]) ? node17949 : 4'b0010;
																assign node17949 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node17952 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node17955 = (inp[0]) ? node17965 : node17956;
													assign node17956 = (inp[13]) ? node17962 : node17957;
														assign node17957 = (inp[2]) ? node17959 : 4'b0110;
															assign node17959 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node17962 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node17965 = (inp[2]) ? node17967 : 4'b0110;
														assign node17967 = (inp[9]) ? node17969 : 4'b0110;
															assign node17969 = (inp[13]) ? 4'b0111 : node17970;
																assign node17970 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node17974 = (inp[12]) ? node17994 : node17975;
												assign node17975 = (inp[0]) ? node17985 : node17976;
													assign node17976 = (inp[11]) ? node17980 : node17977;
														assign node17977 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node17980 = (inp[13]) ? 4'b0011 : node17981;
															assign node17981 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node17985 = (inp[13]) ? 4'b0010 : node17986;
														assign node17986 = (inp[11]) ? node17990 : node17987;
															assign node17987 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node17990 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node17994 = (inp[13]) ? node18002 : node17995;
													assign node17995 = (inp[11]) ? 4'b0010 : node17996;
														assign node17996 = (inp[0]) ? node17998 : 4'b0010;
															assign node17998 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node18002 = (inp[0]) ? node18006 : node18003;
														assign node18003 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18006 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node18009 = (inp[7]) ? node18049 : node18010;
											assign node18010 = (inp[12]) ? node18030 : node18011;
												assign node18011 = (inp[11]) ? node18021 : node18012;
													assign node18012 = (inp[13]) ? node18018 : node18013;
														assign node18013 = (inp[0]) ? node18015 : 4'b0111;
															assign node18015 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node18018 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node18021 = (inp[0]) ? node18025 : node18022;
														assign node18022 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node18025 = (inp[13]) ? 4'b0110 : node18026;
															assign node18026 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node18030 = (inp[13]) ? node18040 : node18031;
													assign node18031 = (inp[9]) ? node18033 : 4'b0010;
														assign node18033 = (inp[11]) ? node18037 : node18034;
															assign node18034 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node18037 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node18040 = (inp[0]) ? 4'b0011 : node18041;
														assign node18041 = (inp[11]) ? node18045 : node18042;
															assign node18042 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node18045 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node18049 = (inp[13]) ? node18067 : node18050;
												assign node18050 = (inp[0]) ? node18058 : node18051;
													assign node18051 = (inp[2]) ? node18055 : node18052;
														assign node18052 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node18055 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node18058 = (inp[9]) ? 4'b0111 : node18059;
														assign node18059 = (inp[11]) ? node18063 : node18060;
															assign node18060 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node18063 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node18067 = (inp[0]) ? node18071 : node18068;
													assign node18068 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node18071 = (inp[11]) ? 4'b0110 : 4'b0111;
									assign node18074 = (inp[1]) ? node18180 : node18075;
										assign node18075 = (inp[7]) ? node18127 : node18076;
											assign node18076 = (inp[12]) ? node18100 : node18077;
												assign node18077 = (inp[2]) ? node18089 : node18078;
													assign node18078 = (inp[13]) ? node18084 : node18079;
														assign node18079 = (inp[9]) ? 4'b0111 : node18080;
															assign node18080 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node18084 = (inp[0]) ? node18086 : 4'b0110;
															assign node18086 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node18089 = (inp[13]) ? node18091 : 4'b0110;
														assign node18091 = (inp[9]) ? node18093 : 4'b0110;
															assign node18093 = (inp[0]) ? node18097 : node18094;
																assign node18094 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node18097 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node18100 = (inp[9]) ? node18120 : node18101;
													assign node18101 = (inp[0]) ? node18111 : node18102;
														assign node18102 = (inp[2]) ? node18104 : 4'b0010;
															assign node18104 = (inp[13]) ? node18108 : node18105;
																assign node18105 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node18108 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18111 = (inp[2]) ? node18113 : 4'b0011;
															assign node18113 = (inp[11]) ? node18117 : node18114;
																assign node18114 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node18117 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node18120 = (inp[13]) ? node18122 : 4'b0010;
														assign node18122 = (inp[11]) ? node18124 : 4'b0010;
															assign node18124 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node18127 = (inp[9]) ? node18161 : node18128;
												assign node18128 = (inp[0]) ? node18138 : node18129;
													assign node18129 = (inp[11]) ? 4'b0111 : node18130;
														assign node18130 = (inp[12]) ? node18134 : node18131;
															assign node18131 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node18134 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node18138 = (inp[13]) ? node18148 : node18139;
														assign node18139 = (inp[2]) ? 4'b0110 : node18140;
															assign node18140 = (inp[11]) ? node18144 : node18141;
																assign node18141 = (inp[12]) ? 4'b0111 : 4'b0110;
																assign node18144 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node18148 = (inp[12]) ? node18154 : node18149;
															assign node18149 = (inp[11]) ? node18151 : 4'b0111;
																assign node18151 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node18154 = (inp[11]) ? node18158 : node18155;
																assign node18155 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node18158 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node18161 = (inp[0]) ? node18169 : node18162;
													assign node18162 = (inp[12]) ? 4'b0110 : node18163;
														assign node18163 = (inp[11]) ? 4'b0110 : node18164;
															assign node18164 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node18169 = (inp[11]) ? node18177 : node18170;
														assign node18170 = (inp[12]) ? 4'b0111 : node18171;
															assign node18171 = (inp[13]) ? node18173 : 4'b0110;
																assign node18173 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node18177 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node18180 = (inp[7]) ? node18210 : node18181;
											assign node18181 = (inp[12]) ? node18197 : node18182;
												assign node18182 = (inp[0]) ? node18194 : node18183;
													assign node18183 = (inp[9]) ? node18187 : node18184;
														assign node18184 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node18187 = (inp[13]) ? 4'b0011 : node18188;
															assign node18188 = (inp[11]) ? node18190 : 4'b0010;
																assign node18190 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node18194 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node18197 = (inp[0]) ? node18205 : node18198;
													assign node18198 = (inp[9]) ? node18200 : 4'b0111;
														assign node18200 = (inp[13]) ? 4'b0110 : node18201;
															assign node18201 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node18205 = (inp[2]) ? 4'b0110 : node18206;
														assign node18206 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node18210 = (inp[9]) ? node18228 : node18211;
												assign node18211 = (inp[0]) ? node18221 : node18212;
													assign node18212 = (inp[2]) ? node18214 : 4'b0011;
														assign node18214 = (inp[12]) ? 4'b0011 : node18215;
															assign node18215 = (inp[11]) ? 4'b0010 : node18216;
																assign node18216 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node18221 = (inp[11]) ? node18223 : 4'b0011;
														assign node18223 = (inp[2]) ? node18225 : 4'b0010;
															assign node18225 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node18228 = (inp[0]) ? node18230 : 4'b0010;
													assign node18230 = (inp[2]) ? node18234 : node18231;
														assign node18231 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18234 = (inp[11]) ? node18236 : 4'b0010;
															assign node18236 = (inp[13]) ? 4'b0010 : 4'b0011;
								assign node18239 = (inp[7]) ? node18409 : node18240;
									assign node18240 = (inp[0]) ? node18326 : node18241;
										assign node18241 = (inp[11]) ? node18291 : node18242;
											assign node18242 = (inp[13]) ? node18274 : node18243;
												assign node18243 = (inp[5]) ? node18257 : node18244;
													assign node18244 = (inp[2]) ? node18248 : node18245;
														assign node18245 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node18248 = (inp[9]) ? node18250 : 4'b0011;
															assign node18250 = (inp[1]) ? node18254 : node18251;
																assign node18251 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node18254 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node18257 = (inp[2]) ? node18267 : node18258;
														assign node18258 = (inp[9]) ? node18260 : 4'b0011;
															assign node18260 = (inp[12]) ? node18264 : node18261;
																assign node18261 = (inp[1]) ? 4'b0011 : 4'b0110;
																assign node18264 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node18267 = (inp[9]) ? 4'b0010 : node18268;
															assign node18268 = (inp[12]) ? 4'b0111 : node18269;
																assign node18269 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node18274 = (inp[5]) ? node18284 : node18275;
													assign node18275 = (inp[1]) ? node18279 : node18276;
														assign node18276 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node18279 = (inp[12]) ? node18281 : 4'b0110;
															assign node18281 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node18284 = (inp[1]) ? node18288 : node18285;
														assign node18285 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node18288 = (inp[2]) ? 4'b0011 : 4'b0110;
											assign node18291 = (inp[1]) ? node18305 : node18292;
												assign node18292 = (inp[12]) ? node18300 : node18293;
													assign node18293 = (inp[5]) ? 4'b0111 : node18294;
														assign node18294 = (inp[13]) ? 4'b0011 : node18295;
															assign node18295 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node18300 = (inp[5]) ? node18302 : 4'b0111;
														assign node18302 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node18305 = (inp[2]) ? node18313 : node18306;
													assign node18306 = (inp[12]) ? node18310 : node18307;
														assign node18307 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node18310 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node18313 = (inp[13]) ? node18319 : node18314;
														assign node18314 = (inp[5]) ? 4'b0110 : node18315;
															assign node18315 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node18319 = (inp[12]) ? node18323 : node18320;
															assign node18320 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node18323 = (inp[5]) ? 4'b0111 : 4'b0010;
										assign node18326 = (inp[12]) ? node18362 : node18327;
											assign node18327 = (inp[11]) ? node18345 : node18328;
												assign node18328 = (inp[1]) ? node18340 : node18329;
													assign node18329 = (inp[5]) ? node18335 : node18330;
														assign node18330 = (inp[2]) ? node18332 : 4'b0011;
															assign node18332 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node18335 = (inp[13]) ? node18337 : 4'b0111;
															assign node18337 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node18340 = (inp[5]) ? 4'b0010 : node18341;
														assign node18341 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node18345 = (inp[2]) ? node18355 : node18346;
													assign node18346 = (inp[5]) ? node18350 : node18347;
														assign node18347 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node18350 = (inp[1]) ? 4'b0011 : node18351;
															assign node18351 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node18355 = (inp[5]) ? node18359 : node18356;
														assign node18356 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node18359 = (inp[1]) ? 4'b0010 : 4'b0110;
											assign node18362 = (inp[11]) ? node18382 : node18363;
												assign node18363 = (inp[2]) ? node18371 : node18364;
													assign node18364 = (inp[5]) ? node18368 : node18365;
														assign node18365 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node18368 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node18371 = (inp[13]) ? node18373 : 4'b0110;
														assign node18373 = (inp[9]) ? 4'b0010 : node18374;
															assign node18374 = (inp[1]) ? node18378 : node18375;
																assign node18375 = (inp[5]) ? 4'b0010 : 4'b0111;
																assign node18378 = (inp[5]) ? 4'b0111 : 4'b0010;
												assign node18382 = (inp[2]) ? node18398 : node18383;
													assign node18383 = (inp[13]) ? node18391 : node18384;
														assign node18384 = (inp[9]) ? node18386 : 4'b0011;
															assign node18386 = (inp[5]) ? 4'b0110 : node18387;
																assign node18387 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node18391 = (inp[1]) ? node18395 : node18392;
															assign node18392 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node18395 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node18398 = (inp[1]) ? node18406 : node18399;
														assign node18399 = (inp[5]) ? node18403 : node18400;
															assign node18400 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node18403 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node18406 = (inp[5]) ? 4'b0111 : 4'b0011;
									assign node18409 = (inp[13]) ? node18501 : node18410;
										assign node18410 = (inp[2]) ? node18462 : node18411;
											assign node18411 = (inp[12]) ? node18439 : node18412;
												assign node18412 = (inp[11]) ? node18428 : node18413;
													assign node18413 = (inp[0]) ? node18421 : node18414;
														assign node18414 = (inp[1]) ? node18418 : node18415;
															assign node18415 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node18418 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node18421 = (inp[1]) ? node18425 : node18422;
															assign node18422 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node18425 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node18428 = (inp[1]) ? node18436 : node18429;
														assign node18429 = (inp[5]) ? node18433 : node18430;
															assign node18430 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node18433 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node18436 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node18439 = (inp[0]) ? node18447 : node18440;
													assign node18440 = (inp[5]) ? node18444 : node18441;
														assign node18441 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node18444 = (inp[9]) ? 4'b0110 : 4'b0011;
													assign node18447 = (inp[11]) ? node18455 : node18448;
														assign node18448 = (inp[9]) ? node18450 : 4'b0111;
															assign node18450 = (inp[1]) ? 4'b0111 : node18451;
																assign node18451 = (inp[5]) ? 4'b0111 : 4'b0010;
														assign node18455 = (inp[1]) ? node18459 : node18456;
															assign node18456 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node18459 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node18462 = (inp[5]) ? node18486 : node18463;
												assign node18463 = (inp[1]) ? node18481 : node18464;
													assign node18464 = (inp[0]) ? node18470 : node18465;
														assign node18465 = (inp[11]) ? 4'b0010 : node18466;
															assign node18466 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node18470 = (inp[9]) ? node18476 : node18471;
															assign node18471 = (inp[11]) ? node18473 : 4'b0010;
																assign node18473 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node18476 = (inp[11]) ? node18478 : 4'b0011;
																assign node18478 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node18481 = (inp[11]) ? node18483 : 4'b0110;
														assign node18483 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node18486 = (inp[1]) ? node18492 : node18487;
													assign node18487 = (inp[12]) ? node18489 : 4'b0111;
														assign node18489 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node18492 = (inp[12]) ? node18494 : 4'b0011;
														assign node18494 = (inp[0]) ? node18498 : node18495;
															assign node18495 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node18498 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node18501 = (inp[5]) ? node18531 : node18502;
											assign node18502 = (inp[1]) ? node18518 : node18503;
												assign node18503 = (inp[0]) ? node18509 : node18504;
													assign node18504 = (inp[9]) ? 4'b0010 : node18505;
														assign node18505 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node18509 = (inp[9]) ? node18511 : 4'b0011;
														assign node18511 = (inp[2]) ? 4'b0010 : node18512;
															assign node18512 = (inp[11]) ? node18514 : 4'b0011;
																assign node18514 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node18518 = (inp[9]) ? node18524 : node18519;
													assign node18519 = (inp[11]) ? node18521 : 4'b0110;
														assign node18521 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node18524 = (inp[0]) ? node18528 : node18525;
														assign node18525 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node18528 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node18531 = (inp[1]) ? node18563 : node18532;
												assign node18532 = (inp[12]) ? node18546 : node18533;
													assign node18533 = (inp[11]) ? 4'b0110 : node18534;
														assign node18534 = (inp[9]) ? node18540 : node18535;
															assign node18535 = (inp[2]) ? node18537 : 4'b0110;
																assign node18537 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node18540 = (inp[2]) ? node18542 : 4'b0111;
																assign node18542 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node18546 = (inp[2]) ? node18556 : node18547;
														assign node18547 = (inp[9]) ? node18551 : node18548;
															assign node18548 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node18551 = (inp[0]) ? node18553 : 4'b0111;
																assign node18553 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node18556 = (inp[0]) ? node18560 : node18557;
															assign node18557 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node18560 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node18563 = (inp[2]) ? node18567 : node18564;
													assign node18564 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node18567 = (inp[12]) ? 4'b0011 : node18568;
														assign node18568 = (inp[9]) ? 4'b0010 : 4'b0011;
							assign node18572 = (inp[10]) ? node18864 : node18573;
								assign node18573 = (inp[5]) ? node18701 : node18574;
									assign node18574 = (inp[1]) ? node18636 : node18575;
										assign node18575 = (inp[12]) ? node18607 : node18576;
											assign node18576 = (inp[7]) ? node18594 : node18577;
												assign node18577 = (inp[0]) ? node18583 : node18578;
													assign node18578 = (inp[11]) ? 4'b0100 : node18579;
														assign node18579 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node18583 = (inp[11]) ? node18589 : node18584;
														assign node18584 = (inp[13]) ? 4'b0100 : node18585;
															assign node18585 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18589 = (inp[13]) ? 4'b0101 : node18590;
															assign node18590 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node18594 = (inp[11]) ? node18598 : node18595;
													assign node18595 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node18598 = (inp[0]) ? node18604 : node18599;
														assign node18599 = (inp[13]) ? node18601 : 4'b0001;
															assign node18601 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node18604 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node18607 = (inp[9]) ? node18623 : node18608;
												assign node18608 = (inp[2]) ? node18618 : node18609;
													assign node18609 = (inp[13]) ? node18611 : 4'b0001;
														assign node18611 = (inp[11]) ? node18613 : 4'b0000;
															assign node18613 = (inp[0]) ? 4'b0000 : node18614;
																assign node18614 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18618 = (inp[13]) ? 4'b0001 : node18619;
														assign node18619 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node18623 = (inp[13]) ? 4'b0000 : node18624;
													assign node18624 = (inp[11]) ? node18630 : node18625;
														assign node18625 = (inp[7]) ? node18627 : 4'b0000;
															assign node18627 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node18630 = (inp[0]) ? 4'b0001 : node18631;
															assign node18631 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node18636 = (inp[12]) ? node18662 : node18637;
											assign node18637 = (inp[7]) ? node18657 : node18638;
												assign node18638 = (inp[9]) ? node18646 : node18639;
													assign node18639 = (inp[11]) ? 4'b0000 : node18640;
														assign node18640 = (inp[0]) ? node18642 : 4'b0000;
															assign node18642 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node18646 = (inp[13]) ? node18654 : node18647;
														assign node18647 = (inp[2]) ? 4'b0000 : node18648;
															assign node18648 = (inp[0]) ? node18650 : 4'b0001;
																assign node18650 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node18654 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node18657 = (inp[0]) ? node18659 : 4'b0100;
													assign node18659 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node18662 = (inp[7]) ? node18680 : node18663;
												assign node18663 = (inp[0]) ? node18675 : node18664;
													assign node18664 = (inp[11]) ? node18670 : node18665;
														assign node18665 = (inp[13]) ? 4'b0101 : node18666;
															assign node18666 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node18670 = (inp[13]) ? 4'b0100 : node18671;
															assign node18671 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node18675 = (inp[2]) ? node18677 : 4'b0101;
														assign node18677 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node18680 = (inp[11]) ? node18692 : node18681;
													assign node18681 = (inp[0]) ? node18687 : node18682;
														assign node18682 = (inp[13]) ? 4'b0100 : node18683;
															assign node18683 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18687 = (inp[2]) ? 4'b0101 : node18688;
															assign node18688 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node18692 = (inp[0]) ? node18696 : node18693;
														assign node18693 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node18696 = (inp[13]) ? 4'b0100 : node18697;
															assign node18697 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node18701 = (inp[1]) ? node18781 : node18702;
										assign node18702 = (inp[12]) ? node18746 : node18703;
											assign node18703 = (inp[7]) ? node18717 : node18704;
												assign node18704 = (inp[0]) ? node18710 : node18705;
													assign node18705 = (inp[11]) ? 4'b0001 : node18706;
														assign node18706 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node18710 = (inp[11]) ? 4'b0000 : node18711;
														assign node18711 = (inp[2]) ? 4'b0001 : node18712;
															assign node18712 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node18717 = (inp[9]) ? node18733 : node18718;
													assign node18718 = (inp[13]) ? node18722 : node18719;
														assign node18719 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18722 = (inp[2]) ? node18728 : node18723;
															assign node18723 = (inp[11]) ? node18725 : 4'b0100;
																assign node18725 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node18728 = (inp[11]) ? 4'b0101 : node18729;
																assign node18729 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node18733 = (inp[0]) ? node18741 : node18734;
														assign node18734 = (inp[11]) ? 4'b0100 : node18735;
															assign node18735 = (inp[2]) ? 4'b0101 : node18736;
																assign node18736 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node18741 = (inp[11]) ? node18743 : 4'b0100;
															assign node18743 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node18746 = (inp[7]) ? node18768 : node18747;
												assign node18747 = (inp[0]) ? node18757 : node18748;
													assign node18748 = (inp[11]) ? node18752 : node18749;
														assign node18749 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18752 = (inp[2]) ? 4'b0101 : node18753;
															assign node18753 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node18757 = (inp[11]) ? node18763 : node18758;
														assign node18758 = (inp[2]) ? 4'b0101 : node18759;
															assign node18759 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node18763 = (inp[2]) ? 4'b0100 : node18764;
															assign node18764 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node18768 = (inp[11]) ? node18776 : node18769;
													assign node18769 = (inp[13]) ? 4'b0101 : node18770;
														assign node18770 = (inp[2]) ? 4'b0100 : node18771;
															assign node18771 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node18776 = (inp[9]) ? 4'b0101 : node18777;
														assign node18777 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node18781 = (inp[7]) ? node18825 : node18782;
											assign node18782 = (inp[12]) ? node18814 : node18783;
												assign node18783 = (inp[0]) ? node18795 : node18784;
													assign node18784 = (inp[11]) ? node18790 : node18785;
														assign node18785 = (inp[13]) ? node18787 : 4'b0101;
															assign node18787 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node18790 = (inp[13]) ? node18792 : 4'b0100;
															assign node18792 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node18795 = (inp[9]) ? node18805 : node18796;
														assign node18796 = (inp[11]) ? node18802 : node18797;
															assign node18797 = (inp[13]) ? node18799 : 4'b0100;
																assign node18799 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node18802 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18805 = (inp[2]) ? node18809 : node18806;
															assign node18806 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node18809 = (inp[11]) ? node18811 : 4'b0101;
																assign node18811 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node18814 = (inp[2]) ? node18820 : node18815;
													assign node18815 = (inp[9]) ? node18817 : 4'b0000;
														assign node18817 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node18820 = (inp[11]) ? node18822 : 4'b0001;
														assign node18822 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node18825 = (inp[13]) ? node18851 : node18826;
												assign node18826 = (inp[12]) ? node18836 : node18827;
													assign node18827 = (inp[2]) ? node18829 : 4'b0001;
														assign node18829 = (inp[0]) ? node18833 : node18830;
															assign node18830 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node18833 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node18836 = (inp[11]) ? node18844 : node18837;
														assign node18837 = (inp[2]) ? node18841 : node18838;
															assign node18838 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node18841 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node18844 = (inp[9]) ? node18846 : 4'b0001;
															assign node18846 = (inp[0]) ? node18848 : 4'b0000;
																assign node18848 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node18851 = (inp[2]) ? node18857 : node18852;
													assign node18852 = (inp[11]) ? 4'b0000 : node18853;
														assign node18853 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node18857 = (inp[0]) ? node18861 : node18858;
														assign node18858 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node18861 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node18864 = (inp[5]) ? node19020 : node18865;
									assign node18865 = (inp[1]) ? node18945 : node18866;
										assign node18866 = (inp[7]) ? node18904 : node18867;
											assign node18867 = (inp[12]) ? node18877 : node18868;
												assign node18868 = (inp[2]) ? 4'b0100 : node18869;
													assign node18869 = (inp[13]) ? node18873 : node18870;
														assign node18870 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node18873 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node18877 = (inp[9]) ? node18891 : node18878;
													assign node18878 = (inp[13]) ? 4'b0001 : node18879;
														assign node18879 = (inp[2]) ? node18885 : node18880;
															assign node18880 = (inp[0]) ? node18882 : 4'b0001;
																assign node18882 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node18885 = (inp[11]) ? node18887 : 4'b0000;
																assign node18887 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node18891 = (inp[13]) ? node18899 : node18892;
														assign node18892 = (inp[2]) ? node18894 : 4'b0000;
															assign node18894 = (inp[0]) ? 4'b0001 : node18895;
																assign node18895 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node18899 = (inp[11]) ? 4'b0000 : node18900;
															assign node18900 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node18904 = (inp[0]) ? node18928 : node18905;
												assign node18905 = (inp[12]) ? node18917 : node18906;
													assign node18906 = (inp[9]) ? 4'b0000 : node18907;
														assign node18907 = (inp[11]) ? node18913 : node18908;
															assign node18908 = (inp[2]) ? node18910 : 4'b0000;
																assign node18910 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node18913 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node18917 = (inp[11]) ? node18923 : node18918;
														assign node18918 = (inp[9]) ? 4'b0001 : node18919;
															assign node18919 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node18923 = (inp[2]) ? node18925 : 4'b0000;
															assign node18925 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node18928 = (inp[11]) ? node18934 : node18929;
													assign node18929 = (inp[12]) ? node18931 : 4'b0001;
														assign node18931 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node18934 = (inp[12]) ? node18940 : node18935;
														assign node18935 = (inp[2]) ? node18937 : 4'b0000;
															assign node18937 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node18940 = (inp[2]) ? node18942 : 4'b0001;
															assign node18942 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node18945 = (inp[7]) ? node18991 : node18946;
											assign node18946 = (inp[12]) ? node18982 : node18947;
												assign node18947 = (inp[9]) ? node18967 : node18948;
													assign node18948 = (inp[2]) ? node18962 : node18949;
														assign node18949 = (inp[13]) ? node18955 : node18950;
															assign node18950 = (inp[11]) ? node18952 : 4'b0001;
																assign node18952 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node18955 = (inp[11]) ? node18959 : node18956;
																assign node18956 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node18959 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node18962 = (inp[11]) ? 4'b0001 : node18963;
															assign node18963 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node18967 = (inp[11]) ? node18977 : node18968;
														assign node18968 = (inp[2]) ? 4'b0001 : node18969;
															assign node18969 = (inp[13]) ? node18973 : node18970;
																assign node18970 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node18973 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node18977 = (inp[0]) ? 4'b0000 : node18978;
															assign node18978 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node18982 = (inp[0]) ? node18986 : node18983;
													assign node18983 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node18986 = (inp[9]) ? node18988 : 4'b0100;
														assign node18988 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node18991 = (inp[0]) ? node19003 : node18992;
												assign node18992 = (inp[11]) ? node18998 : node18993;
													assign node18993 = (inp[13]) ? 4'b0100 : node18994;
														assign node18994 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node18998 = (inp[13]) ? 4'b0101 : node18999;
														assign node18999 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node19003 = (inp[12]) ? node19013 : node19004;
													assign node19004 = (inp[2]) ? 4'b0100 : node19005;
														assign node19005 = (inp[9]) ? node19007 : 4'b0101;
															assign node19007 = (inp[13]) ? 4'b0100 : node19008;
																assign node19008 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node19013 = (inp[13]) ? 4'b0101 : node19014;
														assign node19014 = (inp[2]) ? 4'b0101 : node19015;
															assign node19015 = (inp[11]) ? 4'b0101 : 4'b0100;
									assign node19020 = (inp[1]) ? node19108 : node19021;
										assign node19021 = (inp[12]) ? node19069 : node19022;
											assign node19022 = (inp[7]) ? node19046 : node19023;
												assign node19023 = (inp[9]) ? node19029 : node19024;
													assign node19024 = (inp[0]) ? node19026 : 4'b0000;
														assign node19026 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node19029 = (inp[13]) ? node19041 : node19030;
														assign node19030 = (inp[0]) ? node19036 : node19031;
															assign node19031 = (inp[2]) ? 4'b0001 : node19032;
																assign node19032 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node19036 = (inp[2]) ? 4'b0000 : node19037;
																assign node19037 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node19041 = (inp[11]) ? 4'b0000 : node19042;
															assign node19042 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node19046 = (inp[9]) ? node19054 : node19047;
													assign node19047 = (inp[0]) ? 4'b0101 : node19048;
														assign node19048 = (inp[2]) ? node19050 : 4'b0101;
															assign node19050 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19054 = (inp[0]) ? node19060 : node19055;
														assign node19055 = (inp[11]) ? node19057 : 4'b0101;
															assign node19057 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node19060 = (inp[13]) ? 4'b0100 : node19061;
															assign node19061 = (inp[11]) ? node19065 : node19062;
																assign node19062 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node19065 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node19069 = (inp[7]) ? node19091 : node19070;
												assign node19070 = (inp[0]) ? node19080 : node19071;
													assign node19071 = (inp[13]) ? 4'b0101 : node19072;
														assign node19072 = (inp[2]) ? node19076 : node19073;
															assign node19073 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node19076 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node19080 = (inp[11]) ? node19086 : node19081;
														assign node19081 = (inp[13]) ? 4'b0101 : node19082;
															assign node19082 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node19086 = (inp[13]) ? 4'b0100 : node19087;
															assign node19087 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node19091 = (inp[9]) ? node19093 : 4'b0100;
													assign node19093 = (inp[13]) ? node19103 : node19094;
														assign node19094 = (inp[2]) ? 4'b0100 : node19095;
															assign node19095 = (inp[0]) ? node19099 : node19096;
																assign node19096 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node19099 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node19103 = (inp[2]) ? 4'b0101 : node19104;
															assign node19104 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node19108 = (inp[7]) ? node19150 : node19109;
											assign node19109 = (inp[12]) ? node19135 : node19110;
												assign node19110 = (inp[0]) ? node19122 : node19111;
													assign node19111 = (inp[11]) ? node19117 : node19112;
														assign node19112 = (inp[2]) ? node19114 : 4'b0101;
															assign node19114 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node19117 = (inp[13]) ? node19119 : 4'b0100;
															assign node19119 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node19122 = (inp[2]) ? node19124 : 4'b0100;
														assign node19124 = (inp[9]) ? node19130 : node19125;
															assign node19125 = (inp[11]) ? node19127 : 4'b0100;
																assign node19127 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node19130 = (inp[13]) ? 4'b0101 : node19131;
																assign node19131 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node19135 = (inp[13]) ? node19143 : node19136;
													assign node19136 = (inp[11]) ? 4'b0000 : node19137;
														assign node19137 = (inp[9]) ? node19139 : 4'b0000;
															assign node19139 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node19143 = (inp[2]) ? node19147 : node19144;
														assign node19144 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node19147 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node19150 = (inp[9]) ? node19166 : node19151;
												assign node19151 = (inp[11]) ? node19159 : node19152;
													assign node19152 = (inp[0]) ? 4'b0001 : node19153;
														assign node19153 = (inp[2]) ? 4'b0000 : node19154;
															assign node19154 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node19159 = (inp[0]) ? 4'b0000 : node19160;
														assign node19160 = (inp[12]) ? 4'b0001 : node19161;
															assign node19161 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node19166 = (inp[11]) ? node19174 : node19167;
													assign node19167 = (inp[0]) ? node19171 : node19168;
														assign node19168 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node19171 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19174 = (inp[2]) ? 4'b0001 : node19175;
														assign node19175 = (inp[12]) ? 4'b0000 : node19176;
															assign node19176 = (inp[13]) ? 4'b0000 : 4'b0001;
						assign node19181 = (inp[1]) ? node19611 : node19182;
							assign node19182 = (inp[15]) ? node19334 : node19183;
								assign node19183 = (inp[7]) ? node19327 : node19184;
									assign node19184 = (inp[10]) ? node19274 : node19185;
										assign node19185 = (inp[11]) ? node19229 : node19186;
											assign node19186 = (inp[9]) ? node19220 : node19187;
												assign node19187 = (inp[13]) ? node19201 : node19188;
													assign node19188 = (inp[2]) ? node19196 : node19189;
														assign node19189 = (inp[0]) ? node19193 : node19190;
															assign node19190 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node19193 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node19196 = (inp[12]) ? 4'b0000 : node19197;
															assign node19197 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node19201 = (inp[2]) ? node19215 : node19202;
														assign node19202 = (inp[5]) ? node19208 : node19203;
															assign node19203 = (inp[12]) ? 4'b0001 : node19204;
																assign node19204 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node19208 = (inp[12]) ? node19212 : node19209;
																assign node19209 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node19212 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19215 = (inp[12]) ? node19217 : 4'b0001;
															assign node19217 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node19220 = (inp[13]) ? 4'b0000 : node19221;
													assign node19221 = (inp[12]) ? node19223 : 4'b0001;
														assign node19223 = (inp[0]) ? node19225 : 4'b0000;
															assign node19225 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node19229 = (inp[13]) ? node19239 : node19230;
												assign node19230 = (inp[9]) ? 4'b0001 : node19231;
													assign node19231 = (inp[5]) ? node19235 : node19232;
														assign node19232 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19235 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node19239 = (inp[2]) ? node19255 : node19240;
													assign node19240 = (inp[9]) ? node19248 : node19241;
														assign node19241 = (inp[0]) ? node19243 : 4'b0001;
															assign node19243 = (inp[12]) ? node19245 : 4'b0000;
																assign node19245 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node19248 = (inp[5]) ? 4'b0000 : node19249;
															assign node19249 = (inp[12]) ? 4'b0000 : node19250;
																assign node19250 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node19255 = (inp[12]) ? node19261 : node19256;
														assign node19256 = (inp[9]) ? 4'b0001 : node19257;
															assign node19257 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node19261 = (inp[9]) ? node19267 : node19262;
															assign node19262 = (inp[0]) ? 4'b0001 : node19263;
																assign node19263 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node19267 = (inp[5]) ? node19271 : node19268;
																assign node19268 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node19271 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node19274 = (inp[11]) ? node19298 : node19275;
											assign node19275 = (inp[5]) ? node19287 : node19276;
												assign node19276 = (inp[0]) ? node19282 : node19277;
													assign node19277 = (inp[12]) ? node19279 : 4'b0000;
														assign node19279 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19282 = (inp[13]) ? node19284 : 4'b0001;
														assign node19284 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node19287 = (inp[0]) ? node19293 : node19288;
													assign node19288 = (inp[12]) ? node19290 : 4'b0001;
														assign node19290 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node19293 = (inp[12]) ? node19295 : 4'b0000;
														assign node19295 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node19298 = (inp[13]) ? node19306 : node19299;
												assign node19299 = (inp[0]) ? node19303 : node19300;
													assign node19300 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node19303 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node19306 = (inp[5]) ? node19320 : node19307;
													assign node19307 = (inp[9]) ? node19313 : node19308;
														assign node19308 = (inp[12]) ? 4'b0000 : node19309;
															assign node19309 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19313 = (inp[0]) ? node19317 : node19314;
															assign node19314 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node19317 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node19320 = (inp[12]) ? node19324 : node19321;
														assign node19321 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node19324 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node19327 = (inp[0]) ? node19331 : node19328;
										assign node19328 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node19331 = (inp[12]) ? 4'b0100 : 4'b0101;
								assign node19334 = (inp[2]) ? node19458 : node19335;
									assign node19335 = (inp[10]) ? node19399 : node19336;
										assign node19336 = (inp[13]) ? node19360 : node19337;
											assign node19337 = (inp[0]) ? node19349 : node19338;
												assign node19338 = (inp[5]) ? node19344 : node19339;
													assign node19339 = (inp[12]) ? node19341 : 4'b0100;
														assign node19341 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node19344 = (inp[7]) ? node19346 : 4'b0101;
														assign node19346 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node19349 = (inp[5]) ? node19355 : node19350;
													assign node19350 = (inp[7]) ? node19352 : 4'b0101;
														assign node19352 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node19355 = (inp[12]) ? 4'b0100 : node19356;
														assign node19356 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node19360 = (inp[11]) ? node19386 : node19361;
												assign node19361 = (inp[7]) ? node19375 : node19362;
													assign node19362 = (inp[12]) ? node19370 : node19363;
														assign node19363 = (inp[9]) ? node19365 : 4'b0100;
															assign node19365 = (inp[5]) ? node19367 : 4'b0100;
																assign node19367 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19370 = (inp[9]) ? 4'b0101 : node19371;
															assign node19371 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node19375 = (inp[9]) ? node19381 : node19376;
														assign node19376 = (inp[0]) ? 4'b0101 : node19377;
															assign node19377 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node19381 = (inp[0]) ? node19383 : 4'b0101;
															assign node19383 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node19386 = (inp[5]) ? node19394 : node19387;
													assign node19387 = (inp[12]) ? node19389 : 4'b0100;
														assign node19389 = (inp[0]) ? 4'b0101 : node19390;
															assign node19390 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node19394 = (inp[12]) ? 4'b0100 : node19395;
														assign node19395 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node19399 = (inp[9]) ? node19423 : node19400;
											assign node19400 = (inp[0]) ? node19410 : node19401;
												assign node19401 = (inp[12]) ? node19405 : node19402;
													assign node19402 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node19405 = (inp[5]) ? 4'b0101 : node19406;
														assign node19406 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node19410 = (inp[12]) ? node19418 : node19411;
													assign node19411 = (inp[7]) ? 4'b0101 : node19412;
														assign node19412 = (inp[5]) ? 4'b0101 : node19413;
															assign node19413 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node19418 = (inp[5]) ? 4'b0100 : node19419;
														assign node19419 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node19423 = (inp[7]) ? node19441 : node19424;
												assign node19424 = (inp[12]) ? node19436 : node19425;
													assign node19425 = (inp[13]) ? node19431 : node19426;
														assign node19426 = (inp[5]) ? 4'b0100 : node19427;
															assign node19427 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19431 = (inp[0]) ? node19433 : 4'b0101;
															assign node19433 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node19436 = (inp[5]) ? node19438 : 4'b0100;
														assign node19438 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node19441 = (inp[5]) ? node19447 : node19442;
													assign node19442 = (inp[12]) ? 4'b0101 : node19443;
														assign node19443 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node19447 = (inp[11]) ? node19453 : node19448;
														assign node19448 = (inp[12]) ? node19450 : 4'b0101;
															assign node19450 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node19453 = (inp[12]) ? node19455 : 4'b0100;
															assign node19455 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node19458 = (inp[13]) ? node19520 : node19459;
										assign node19459 = (inp[10]) ? node19487 : node19460;
											assign node19460 = (inp[11]) ? node19472 : node19461;
												assign node19461 = (inp[9]) ? 4'b0100 : node19462;
													assign node19462 = (inp[7]) ? node19464 : 4'b0100;
														assign node19464 = (inp[12]) ? node19468 : node19465;
															assign node19465 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node19468 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node19472 = (inp[12]) ? node19478 : node19473;
													assign node19473 = (inp[0]) ? node19475 : 4'b0100;
														assign node19475 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node19478 = (inp[0]) ? node19484 : node19479;
														assign node19479 = (inp[7]) ? 4'b0101 : node19480;
															assign node19480 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node19484 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node19487 = (inp[11]) ? node19505 : node19488;
												assign node19488 = (inp[5]) ? node19494 : node19489;
													assign node19489 = (inp[0]) ? node19491 : 4'b0100;
														assign node19491 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node19494 = (inp[0]) ? node19500 : node19495;
														assign node19495 = (inp[7]) ? node19497 : 4'b0101;
															assign node19497 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node19500 = (inp[7]) ? node19502 : 4'b0100;
															assign node19502 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node19505 = (inp[0]) ? node19511 : node19506;
													assign node19506 = (inp[5]) ? node19508 : 4'b0100;
														assign node19508 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node19511 = (inp[5]) ? node19517 : node19512;
														assign node19512 = (inp[12]) ? node19514 : 4'b0101;
															assign node19514 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node19517 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node19520 = (inp[7]) ? node19572 : node19521;
											assign node19521 = (inp[9]) ? node19543 : node19522;
												assign node19522 = (inp[11]) ? node19534 : node19523;
													assign node19523 = (inp[10]) ? 4'b0100 : node19524;
														assign node19524 = (inp[5]) ? 4'b0101 : node19525;
															assign node19525 = (inp[12]) ? node19529 : node19526;
																assign node19526 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node19529 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node19534 = (inp[5]) ? node19536 : 4'b0101;
														assign node19536 = (inp[12]) ? node19540 : node19537;
															assign node19537 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node19540 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node19543 = (inp[0]) ? node19559 : node19544;
													assign node19544 = (inp[10]) ? node19552 : node19545;
														assign node19545 = (inp[5]) ? node19549 : node19546;
															assign node19546 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node19549 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node19552 = (inp[12]) ? node19556 : node19553;
															assign node19553 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node19556 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node19559 = (inp[11]) ? node19561 : 4'b0101;
														assign node19561 = (inp[10]) ? node19567 : node19562;
															assign node19562 = (inp[5]) ? 4'b0101 : node19563;
																assign node19563 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node19567 = (inp[5]) ? node19569 : 4'b0101;
																assign node19569 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node19572 = (inp[9]) ? node19594 : node19573;
												assign node19573 = (inp[5]) ? node19581 : node19574;
													assign node19574 = (inp[12]) ? node19578 : node19575;
														assign node19575 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19578 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node19581 = (inp[11]) ? node19589 : node19582;
														assign node19582 = (inp[10]) ? node19584 : 4'b0100;
															assign node19584 = (inp[0]) ? node19586 : 4'b0101;
																assign node19586 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node19589 = (inp[10]) ? 4'b0100 : node19590;
															assign node19590 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node19594 = (inp[10]) ? node19604 : node19595;
													assign node19595 = (inp[5]) ? node19597 : 4'b0100;
														assign node19597 = (inp[0]) ? node19601 : node19598;
															assign node19598 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node19601 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node19604 = (inp[12]) ? node19608 : node19605;
														assign node19605 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19608 = (inp[0]) ? 4'b0100 : 4'b0101;
							assign node19611 = (inp[15]) ? node19809 : node19612;
								assign node19612 = (inp[7]) ? node19734 : node19613;
									assign node19613 = (inp[12]) ? node19643 : node19614;
										assign node19614 = (inp[11]) ? node19636 : node19615;
											assign node19615 = (inp[9]) ? node19629 : node19616;
												assign node19616 = (inp[10]) ? node19624 : node19617;
													assign node19617 = (inp[5]) ? node19621 : node19618;
														assign node19618 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19621 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node19624 = (inp[0]) ? node19626 : 4'b0100;
														assign node19626 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node19629 = (inp[5]) ? node19633 : node19630;
													assign node19630 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node19633 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node19636 = (inp[0]) ? node19640 : node19637;
												assign node19637 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node19640 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node19643 = (inp[9]) ? node19691 : node19644;
											assign node19644 = (inp[5]) ? node19674 : node19645;
												assign node19645 = (inp[2]) ? node19659 : node19646;
													assign node19646 = (inp[11]) ? node19654 : node19647;
														assign node19647 = (inp[0]) ? node19651 : node19648;
															assign node19648 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node19651 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node19654 = (inp[13]) ? 4'b0101 : node19655;
															assign node19655 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node19659 = (inp[11]) ? node19667 : node19660;
														assign node19660 = (inp[10]) ? node19662 : 4'b0100;
															assign node19662 = (inp[0]) ? node19664 : 4'b0100;
																assign node19664 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node19667 = (inp[0]) ? node19671 : node19668;
															assign node19668 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node19671 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node19674 = (inp[10]) ? node19684 : node19675;
													assign node19675 = (inp[2]) ? node19677 : 4'b0101;
														assign node19677 = (inp[13]) ? node19681 : node19678;
															assign node19678 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node19681 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node19684 = (inp[13]) ? node19688 : node19685;
														assign node19685 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node19688 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node19691 = (inp[5]) ? node19717 : node19692;
												assign node19692 = (inp[2]) ? node19712 : node19693;
													assign node19693 = (inp[11]) ? node19705 : node19694;
														assign node19694 = (inp[10]) ? node19700 : node19695;
															assign node19695 = (inp[13]) ? 4'b0101 : node19696;
																assign node19696 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node19700 = (inp[0]) ? node19702 : 4'b0100;
																assign node19702 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node19705 = (inp[13]) ? node19709 : node19706;
															assign node19706 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node19709 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node19712 = (inp[13]) ? node19714 : 4'b0101;
														assign node19714 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node19717 = (inp[10]) ? node19719 : 4'b0100;
													assign node19719 = (inp[11]) ? node19727 : node19720;
														assign node19720 = (inp[0]) ? node19724 : node19721;
															assign node19721 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node19724 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node19727 = (inp[0]) ? node19731 : node19728;
															assign node19728 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node19731 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node19734 = (inp[10]) ? node19774 : node19735;
										assign node19735 = (inp[11]) ? node19767 : node19736;
											assign node19736 = (inp[12]) ? node19758 : node19737;
												assign node19737 = (inp[5]) ? node19747 : node19738;
													assign node19738 = (inp[9]) ? 4'b0000 : node19739;
														assign node19739 = (inp[13]) ? node19743 : node19740;
															assign node19740 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node19743 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node19747 = (inp[9]) ? node19753 : node19748;
														assign node19748 = (inp[13]) ? node19750 : 4'b0000;
															assign node19750 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node19753 = (inp[0]) ? 4'b0001 : node19754;
															assign node19754 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node19758 = (inp[2]) ? node19764 : node19759;
													assign node19759 = (inp[0]) ? node19761 : 4'b0001;
														assign node19761 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node19764 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node19767 = (inp[13]) ? node19771 : node19768;
												assign node19768 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node19771 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node19774 = (inp[9]) ? node19788 : node19775;
											assign node19775 = (inp[5]) ? node19781 : node19776;
												assign node19776 = (inp[0]) ? node19778 : 4'b0001;
													assign node19778 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node19781 = (inp[13]) ? node19785 : node19782;
													assign node19782 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node19785 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node19788 = (inp[12]) ? node19802 : node19789;
												assign node19789 = (inp[2]) ? node19795 : node19790;
													assign node19790 = (inp[0]) ? 4'b0001 : node19791;
														assign node19791 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19795 = (inp[13]) ? node19799 : node19796;
														assign node19796 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19799 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node19802 = (inp[0]) ? node19806 : node19803;
													assign node19803 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19806 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node19809 = (inp[0]) ? node19835 : node19810;
									assign node19810 = (inp[7]) ? 4'b0001 : node19811;
										assign node19811 = (inp[11]) ? node19823 : node19812;
											assign node19812 = (inp[5]) ? node19818 : node19813;
												assign node19813 = (inp[13]) ? 4'b0000 : node19814;
													assign node19814 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node19818 = (inp[12]) ? 4'b0001 : node19819;
													assign node19819 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node19823 = (inp[5]) ? node19829 : node19824;
												assign node19824 = (inp[12]) ? 4'b0000 : node19825;
													assign node19825 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node19829 = (inp[13]) ? 4'b0001 : node19830;
													assign node19830 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node19835 = (inp[7]) ? 4'b0000 : node19836;
										assign node19836 = (inp[5]) ? node19842 : node19837;
											assign node19837 = (inp[12]) ? 4'b0001 : node19838;
												assign node19838 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node19842 = (inp[12]) ? 4'b0000 : node19843;
												assign node19843 = (inp[13]) ? 4'b0000 : 4'b0001;
		assign node19848 = (inp[8]) ? node30032 : node19849;
			assign node19849 = (inp[14]) ? node25325 : node19850;
				assign node19850 = (inp[2]) ? node22758 : node19851;
					assign node19851 = (inp[13]) ? node21327 : node19852;
						assign node19852 = (inp[5]) ? node20576 : node19853;
							assign node19853 = (inp[6]) ? node20231 : node19854;
								assign node19854 = (inp[1]) ? node20052 : node19855;
									assign node19855 = (inp[15]) ? node19957 : node19856;
										assign node19856 = (inp[12]) ? node19918 : node19857;
											assign node19857 = (inp[7]) ? node19891 : node19858;
												assign node19858 = (inp[4]) ? node19870 : node19859;
													assign node19859 = (inp[11]) ? node19865 : node19860;
														assign node19860 = (inp[0]) ? 4'b1000 : node19861;
															assign node19861 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node19865 = (inp[10]) ? node19867 : 4'b1001;
															assign node19867 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node19870 = (inp[0]) ? node19876 : node19871;
														assign node19871 = (inp[11]) ? 4'b1010 : node19872;
															assign node19872 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node19876 = (inp[10]) ? node19884 : node19877;
															assign node19877 = (inp[11]) ? node19881 : node19878;
																assign node19878 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node19881 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node19884 = (inp[11]) ? node19888 : node19885;
																assign node19885 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node19888 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node19891 = (inp[4]) ? node19903 : node19892;
													assign node19892 = (inp[10]) ? node19894 : 4'b1011;
														assign node19894 = (inp[11]) ? node19900 : node19895;
															assign node19895 = (inp[9]) ? node19897 : 4'b1010;
																assign node19897 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node19900 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node19903 = (inp[0]) ? node19911 : node19904;
														assign node19904 = (inp[9]) ? node19908 : node19905;
															assign node19905 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node19908 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node19911 = (inp[11]) ? 4'b1101 : node19912;
															assign node19912 = (inp[9]) ? node19914 : 4'b1101;
																assign node19914 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node19918 = (inp[9]) ? node19940 : node19919;
												assign node19919 = (inp[10]) ? node19927 : node19920;
													assign node19920 = (inp[4]) ? node19922 : 4'b1100;
														assign node19922 = (inp[7]) ? node19924 : 4'b1100;
															assign node19924 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node19927 = (inp[0]) ? node19929 : 4'b1101;
														assign node19929 = (inp[7]) ? node19937 : node19930;
															assign node19930 = (inp[4]) ? node19934 : node19931;
																assign node19931 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node19934 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node19937 = (inp[4]) ? 4'b1011 : 4'b1101;
												assign node19940 = (inp[4]) ? node19948 : node19941;
													assign node19941 = (inp[7]) ? 4'b1100 : node19942;
														assign node19942 = (inp[10]) ? 4'b1010 : node19943;
															assign node19943 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19948 = (inp[7]) ? node19954 : node19949;
														assign node19949 = (inp[11]) ? node19951 : 4'b1101;
															assign node19951 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node19954 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node19957 = (inp[12]) ? node20003 : node19958;
											assign node19958 = (inp[7]) ? node19976 : node19959;
												assign node19959 = (inp[4]) ? node19969 : node19960;
													assign node19960 = (inp[11]) ? node19962 : 4'b1001;
														assign node19962 = (inp[0]) ? node19964 : 4'b1001;
															assign node19964 = (inp[10]) ? node19966 : 4'b1000;
																assign node19966 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node19969 = (inp[0]) ? 4'b1100 : node19970;
														assign node19970 = (inp[10]) ? 4'b1101 : node19971;
															assign node19971 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node19976 = (inp[4]) ? node19986 : node19977;
													assign node19977 = (inp[11]) ? node19979 : 4'b1111;
														assign node19979 = (inp[0]) ? node19981 : 4'b1111;
															assign node19981 = (inp[10]) ? node19983 : 4'b1110;
																assign node19983 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node19986 = (inp[11]) ? node19994 : node19987;
														assign node19987 = (inp[9]) ? node19991 : node19988;
															assign node19988 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node19991 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node19994 = (inp[10]) ? 4'b1011 : node19995;
															assign node19995 = (inp[0]) ? node19999 : node19996;
																assign node19996 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node19999 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node20003 = (inp[7]) ? node20027 : node20004;
												assign node20004 = (inp[9]) ? node20016 : node20005;
													assign node20005 = (inp[0]) ? node20007 : 4'b1010;
														assign node20007 = (inp[4]) ? 4'b1010 : node20008;
															assign node20008 = (inp[10]) ? node20012 : node20009;
																assign node20009 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node20012 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node20016 = (inp[10]) ? node20018 : 4'b1011;
														assign node20018 = (inp[4]) ? node20024 : node20019;
															assign node20019 = (inp[11]) ? 4'b1010 : node20020;
																assign node20020 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node20024 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node20027 = (inp[0]) ? node20041 : node20028;
													assign node20028 = (inp[4]) ? node20030 : 4'b1001;
														assign node20030 = (inp[9]) ? node20036 : node20031;
															assign node20031 = (inp[10]) ? node20033 : 4'b1001;
																assign node20033 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node20036 = (inp[11]) ? 4'b1000 : node20037;
																assign node20037 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node20041 = (inp[10]) ? node20047 : node20042;
														assign node20042 = (inp[9]) ? 4'b1000 : node20043;
															assign node20043 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20047 = (inp[9]) ? node20049 : 4'b1000;
															assign node20049 = (inp[4]) ? 4'b1001 : 4'b1000;
									assign node20052 = (inp[12]) ? node20154 : node20053;
										assign node20053 = (inp[7]) ? node20101 : node20054;
											assign node20054 = (inp[15]) ? node20076 : node20055;
												assign node20055 = (inp[4]) ? node20067 : node20056;
													assign node20056 = (inp[9]) ? node20060 : node20057;
														assign node20057 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node20060 = (inp[10]) ? 4'b1100 : node20061;
															assign node20061 = (inp[11]) ? 4'b1101 : node20062;
																assign node20062 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node20067 = (inp[10]) ? node20071 : node20068;
														assign node20068 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node20071 = (inp[9]) ? node20073 : 4'b1111;
															assign node20073 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node20076 = (inp[4]) ? node20086 : node20077;
													assign node20077 = (inp[0]) ? node20079 : 4'b1100;
														assign node20079 = (inp[10]) ? node20083 : node20080;
															assign node20080 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node20083 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node20086 = (inp[0]) ? node20094 : node20087;
														assign node20087 = (inp[10]) ? node20091 : node20088;
															assign node20088 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node20091 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node20094 = (inp[9]) ? 4'b1001 : node20095;
															assign node20095 = (inp[10]) ? 4'b1001 : node20096;
																assign node20096 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20101 = (inp[4]) ? node20129 : node20102;
												assign node20102 = (inp[15]) ? node20118 : node20103;
													assign node20103 = (inp[11]) ? node20105 : 4'b1011;
														assign node20105 = (inp[10]) ? node20111 : node20106;
															assign node20106 = (inp[9]) ? 4'b1010 : node20107;
																assign node20107 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node20111 = (inp[0]) ? node20115 : node20112;
																assign node20112 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node20115 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node20118 = (inp[9]) ? node20126 : node20119;
														assign node20119 = (inp[11]) ? 4'b1111 : node20120;
															assign node20120 = (inp[10]) ? node20122 : 4'b1110;
																assign node20122 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node20126 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node20129 = (inp[15]) ? node20141 : node20130;
													assign node20130 = (inp[11]) ? node20136 : node20131;
														assign node20131 = (inp[9]) ? node20133 : 4'b1000;
															assign node20133 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node20136 = (inp[0]) ? node20138 : 4'b1001;
															assign node20138 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node20141 = (inp[9]) ? node20143 : 4'b1010;
														assign node20143 = (inp[10]) ? node20149 : node20144;
															assign node20144 = (inp[11]) ? node20146 : 4'b1010;
																assign node20146 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node20149 = (inp[0]) ? 4'b1011 : node20150;
																assign node20150 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node20154 = (inp[7]) ? node20196 : node20155;
											assign node20155 = (inp[15]) ? node20175 : node20156;
												assign node20156 = (inp[4]) ? node20164 : node20157;
													assign node20157 = (inp[10]) ? 4'b1111 : node20158;
														assign node20158 = (inp[9]) ? node20160 : 4'b1111;
															assign node20160 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node20164 = (inp[10]) ? node20170 : node20165;
														assign node20165 = (inp[11]) ? 4'b1100 : node20166;
															assign node20166 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node20170 = (inp[9]) ? 4'b1101 : node20171;
															assign node20171 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node20175 = (inp[10]) ? node20187 : node20176;
													assign node20176 = (inp[4]) ? node20182 : node20177;
														assign node20177 = (inp[11]) ? 4'b1111 : node20178;
															assign node20178 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node20182 = (inp[11]) ? 4'b1110 : node20183;
															assign node20183 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node20187 = (inp[11]) ? node20189 : 4'b1111;
														assign node20189 = (inp[9]) ? 4'b1110 : node20190;
															assign node20190 = (inp[0]) ? node20192 : 4'b1111;
																assign node20192 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node20196 = (inp[15]) ? node20212 : node20197;
												assign node20197 = (inp[4]) ? node20205 : node20198;
													assign node20198 = (inp[9]) ? node20200 : 4'b1000;
														assign node20200 = (inp[10]) ? node20202 : 4'b1001;
															assign node20202 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node20205 = (inp[10]) ? 4'b1110 : node20206;
														assign node20206 = (inp[0]) ? 4'b1111 : node20207;
															assign node20207 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node20212 = (inp[9]) ? node20224 : node20213;
													assign node20213 = (inp[4]) ? node20219 : node20214;
														assign node20214 = (inp[10]) ? 4'b1101 : node20215;
															assign node20215 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node20219 = (inp[10]) ? 4'b1100 : node20220;
															assign node20220 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node20224 = (inp[11]) ? node20226 : 4'b1100;
														assign node20226 = (inp[10]) ? node20228 : 4'b1100;
															assign node20228 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node20231 = (inp[12]) ? node20431 : node20232;
									assign node20232 = (inp[15]) ? node20336 : node20233;
										assign node20233 = (inp[7]) ? node20283 : node20234;
											assign node20234 = (inp[1]) ? node20256 : node20235;
												assign node20235 = (inp[0]) ? node20243 : node20236;
													assign node20236 = (inp[4]) ? node20238 : 4'b1001;
														assign node20238 = (inp[9]) ? node20240 : 4'b1000;
															assign node20240 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node20243 = (inp[4]) ? node20251 : node20244;
														assign node20244 = (inp[9]) ? node20248 : node20245;
															assign node20245 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node20248 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20251 = (inp[9]) ? node20253 : 4'b1000;
															assign node20253 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node20256 = (inp[4]) ? node20272 : node20257;
													assign node20257 = (inp[11]) ? node20263 : node20258;
														assign node20258 = (inp[10]) ? node20260 : 4'b1101;
															assign node20260 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node20263 = (inp[10]) ? node20267 : node20264;
															assign node20264 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node20267 = (inp[9]) ? node20269 : 4'b1100;
																assign node20269 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node20272 = (inp[10]) ? node20278 : node20273;
														assign node20273 = (inp[11]) ? node20275 : 4'b1000;
															assign node20275 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node20278 = (inp[9]) ? 4'b1001 : node20279;
															assign node20279 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20283 = (inp[1]) ? node20307 : node20284;
												assign node20284 = (inp[4]) ? node20294 : node20285;
													assign node20285 = (inp[11]) ? 4'b1011 : node20286;
														assign node20286 = (inp[10]) ? 4'b1011 : node20287;
															assign node20287 = (inp[9]) ? node20289 : 4'b1010;
																assign node20289 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node20294 = (inp[0]) ? node20302 : node20295;
														assign node20295 = (inp[9]) ? node20299 : node20296;
															assign node20296 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node20299 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node20302 = (inp[11]) ? 4'b1111 : node20303;
															assign node20303 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node20307 = (inp[0]) ? node20323 : node20308;
													assign node20308 = (inp[4]) ? node20318 : node20309;
														assign node20309 = (inp[10]) ? node20311 : 4'b1010;
															assign node20311 = (inp[9]) ? node20315 : node20312;
																assign node20312 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node20315 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20318 = (inp[10]) ? node20320 : 4'b1011;
															assign node20320 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node20323 = (inp[10]) ? node20331 : node20324;
														assign node20324 = (inp[9]) ? node20328 : node20325;
															assign node20325 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node20328 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20331 = (inp[11]) ? 4'b1011 : node20332;
															assign node20332 = (inp[9]) ? 4'b1011 : 4'b1010;
										assign node20336 = (inp[7]) ? node20384 : node20337;
											assign node20337 = (inp[4]) ? node20363 : node20338;
												assign node20338 = (inp[1]) ? node20354 : node20339;
													assign node20339 = (inp[9]) ? node20345 : node20340;
														assign node20340 = (inp[10]) ? node20342 : 4'b1011;
															assign node20342 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node20345 = (inp[10]) ? 4'b1010 : node20346;
															assign node20346 = (inp[11]) ? node20350 : node20347;
																assign node20347 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node20350 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node20354 = (inp[0]) ? 4'b1111 : node20355;
														assign node20355 = (inp[11]) ? node20359 : node20356;
															assign node20356 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node20359 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node20363 = (inp[1]) ? node20373 : node20364;
													assign node20364 = (inp[11]) ? node20366 : 4'b1110;
														assign node20366 = (inp[9]) ? node20370 : node20367;
															assign node20367 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node20370 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node20373 = (inp[9]) ? node20375 : 4'b1010;
														assign node20375 = (inp[10]) ? node20377 : 4'b1010;
															assign node20377 = (inp[11]) ? node20381 : node20378;
																assign node20378 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node20381 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node20384 = (inp[9]) ? node20412 : node20385;
												assign node20385 = (inp[10]) ? node20399 : node20386;
													assign node20386 = (inp[4]) ? node20396 : node20387;
														assign node20387 = (inp[1]) ? node20389 : 4'b1001;
															assign node20389 = (inp[11]) ? node20393 : node20390;
																assign node20390 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node20393 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node20396 = (inp[11]) ? 4'b1000 : 4'b1100;
													assign node20399 = (inp[11]) ? node20405 : node20400;
														assign node20400 = (inp[1]) ? node20402 : 4'b1000;
															assign node20402 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node20405 = (inp[1]) ? node20407 : 4'b1101;
															assign node20407 = (inp[4]) ? 4'b1000 : node20408;
																assign node20408 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node20412 = (inp[1]) ? node20420 : node20413;
													assign node20413 = (inp[11]) ? node20417 : node20414;
														assign node20414 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node20417 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20420 = (inp[4]) ? node20428 : node20421;
														assign node20421 = (inp[0]) ? node20425 : node20422;
															assign node20422 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node20425 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node20428 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node20431 = (inp[15]) ? node20511 : node20432;
										assign node20432 = (inp[7]) ? node20480 : node20433;
											assign node20433 = (inp[4]) ? node20459 : node20434;
												assign node20434 = (inp[10]) ? node20450 : node20435;
													assign node20435 = (inp[0]) ? node20443 : node20436;
														assign node20436 = (inp[9]) ? 4'b1001 : node20437;
															assign node20437 = (inp[1]) ? node20439 : 4'b1001;
																assign node20439 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node20443 = (inp[9]) ? node20447 : node20444;
															assign node20444 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node20447 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node20450 = (inp[1]) ? 4'b1000 : node20451;
														assign node20451 = (inp[0]) ? 4'b1000 : node20452;
															assign node20452 = (inp[9]) ? node20454 : 4'b1001;
																assign node20454 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node20459 = (inp[1]) ? node20469 : node20460;
													assign node20460 = (inp[10]) ? 4'b1000 : node20461;
														assign node20461 = (inp[11]) ? node20465 : node20462;
															assign node20462 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node20465 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node20469 = (inp[10]) ? node20475 : node20470;
														assign node20470 = (inp[9]) ? 4'b1100 : node20471;
															assign node20471 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20475 = (inp[11]) ? 4'b1101 : node20476;
															assign node20476 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node20480 = (inp[4]) ? node20496 : node20481;
												assign node20481 = (inp[1]) ? node20489 : node20482;
													assign node20482 = (inp[9]) ? node20486 : node20483;
														assign node20483 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node20486 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node20489 = (inp[9]) ? node20491 : 4'b1011;
														assign node20491 = (inp[11]) ? node20493 : 4'b1010;
															assign node20493 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node20496 = (inp[9]) ? node20502 : node20497;
													assign node20497 = (inp[11]) ? node20499 : 4'b1010;
														assign node20499 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node20502 = (inp[1]) ? 4'b1011 : node20503;
														assign node20503 = (inp[10]) ? node20505 : 4'b1011;
															assign node20505 = (inp[11]) ? 4'b1010 : node20506;
																assign node20506 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node20511 = (inp[7]) ? node20535 : node20512;
											assign node20512 = (inp[11]) ? node20524 : node20513;
												assign node20513 = (inp[9]) ? node20519 : node20514;
													assign node20514 = (inp[0]) ? node20516 : 4'b1010;
														assign node20516 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node20519 = (inp[4]) ? 4'b1011 : node20520;
														assign node20520 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node20524 = (inp[9]) ? node20530 : node20525;
													assign node20525 = (inp[4]) ? 4'b1011 : node20526;
														assign node20526 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node20530 = (inp[4]) ? 4'b1010 : node20531;
														assign node20531 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node20535 = (inp[4]) ? node20561 : node20536;
												assign node20536 = (inp[0]) ? node20542 : node20537;
													assign node20537 = (inp[11]) ? 4'b1001 : node20538;
														assign node20538 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node20542 = (inp[1]) ? node20552 : node20543;
														assign node20543 = (inp[10]) ? 4'b1001 : node20544;
															assign node20544 = (inp[11]) ? node20548 : node20545;
																assign node20545 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node20548 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node20552 = (inp[10]) ? node20554 : 4'b1001;
															assign node20554 = (inp[11]) ? node20558 : node20555;
																assign node20555 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node20558 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node20561 = (inp[1]) ? node20569 : node20562;
													assign node20562 = (inp[11]) ? node20566 : node20563;
														assign node20563 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node20566 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node20569 = (inp[0]) ? 4'b1001 : node20570;
														assign node20570 = (inp[11]) ? 4'b1000 : node20571;
															assign node20571 = (inp[9]) ? 4'b1000 : 4'b1001;
							assign node20576 = (inp[6]) ? node20976 : node20577;
								assign node20577 = (inp[7]) ? node20771 : node20578;
									assign node20578 = (inp[12]) ? node20680 : node20579;
										assign node20579 = (inp[15]) ? node20627 : node20580;
											assign node20580 = (inp[4]) ? node20596 : node20581;
												assign node20581 = (inp[11]) ? node20587 : node20582;
													assign node20582 = (inp[10]) ? 4'b1001 : node20583;
														assign node20583 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node20587 = (inp[1]) ? 4'b1001 : node20588;
														assign node20588 = (inp[0]) ? 4'b1000 : node20589;
															assign node20589 = (inp[9]) ? 4'b1001 : node20590;
																assign node20590 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node20596 = (inp[1]) ? node20616 : node20597;
													assign node20597 = (inp[11]) ? node20603 : node20598;
														assign node20598 = (inp[9]) ? node20600 : 4'b1011;
															assign node20600 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node20603 = (inp[0]) ? node20611 : node20604;
															assign node20604 = (inp[10]) ? node20608 : node20605;
																assign node20605 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node20608 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node20611 = (inp[10]) ? 4'b1011 : node20612;
																assign node20612 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node20616 = (inp[9]) ? node20620 : node20617;
														assign node20617 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node20620 = (inp[10]) ? node20624 : node20621;
															assign node20621 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node20624 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node20627 = (inp[4]) ? node20657 : node20628;
												assign node20628 = (inp[9]) ? node20642 : node20629;
													assign node20629 = (inp[1]) ? node20635 : node20630;
														assign node20630 = (inp[11]) ? 4'b1001 : node20631;
															assign node20631 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node20635 = (inp[0]) ? node20637 : 4'b1000;
															assign node20637 = (inp[11]) ? 4'b1000 : node20638;
																assign node20638 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node20642 = (inp[0]) ? node20648 : node20643;
														assign node20643 = (inp[1]) ? 4'b1001 : node20644;
															assign node20644 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node20648 = (inp[1]) ? node20650 : 4'b1000;
															assign node20650 = (inp[10]) ? node20654 : node20651;
																assign node20651 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node20654 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node20657 = (inp[0]) ? node20667 : node20658;
													assign node20658 = (inp[11]) ? node20660 : 4'b1101;
														assign node20660 = (inp[10]) ? node20664 : node20661;
															assign node20661 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node20664 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node20667 = (inp[11]) ? node20669 : 4'b1100;
														assign node20669 = (inp[9]) ? node20675 : node20670;
															assign node20670 = (inp[10]) ? node20672 : 4'b1100;
																assign node20672 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node20675 = (inp[1]) ? 4'b1101 : node20676;
																assign node20676 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node20680 = (inp[15]) ? node20720 : node20681;
											assign node20681 = (inp[4]) ? node20703 : node20682;
												assign node20682 = (inp[1]) ? node20692 : node20683;
													assign node20683 = (inp[9]) ? node20687 : node20684;
														assign node20684 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node20687 = (inp[11]) ? node20689 : 4'b1011;
															assign node20689 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node20692 = (inp[10]) ? node20698 : node20693;
														assign node20693 = (inp[9]) ? 4'b1010 : node20694;
															assign node20694 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20698 = (inp[9]) ? node20700 : 4'b1010;
															assign node20700 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node20703 = (inp[1]) ? node20711 : node20704;
													assign node20704 = (inp[0]) ? 4'b1001 : node20705;
														assign node20705 = (inp[11]) ? node20707 : 4'b1000;
															assign node20707 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node20711 = (inp[9]) ? 4'b1100 : node20712;
														assign node20712 = (inp[0]) ? node20716 : node20713;
															assign node20713 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node20716 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node20720 = (inp[0]) ? node20748 : node20721;
												assign node20721 = (inp[1]) ? node20735 : node20722;
													assign node20722 = (inp[9]) ? node20730 : node20723;
														assign node20723 = (inp[4]) ? node20727 : node20724;
															assign node20724 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node20727 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node20730 = (inp[10]) ? 4'b1010 : node20731;
															assign node20731 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node20735 = (inp[9]) ? 4'b1011 : node20736;
														assign node20736 = (inp[11]) ? node20742 : node20737;
															assign node20737 = (inp[4]) ? node20739 : 4'b1011;
																assign node20739 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node20742 = (inp[10]) ? node20744 : 4'b1010;
																assign node20744 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node20748 = (inp[4]) ? node20758 : node20749;
													assign node20749 = (inp[1]) ? 4'b1010 : node20750;
														assign node20750 = (inp[9]) ? 4'b1010 : node20751;
															assign node20751 = (inp[10]) ? 4'b1011 : node20752;
																assign node20752 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20758 = (inp[1]) ? node20764 : node20759;
														assign node20759 = (inp[11]) ? 4'b1010 : node20760;
															assign node20760 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node20764 = (inp[11]) ? 4'b1011 : node20765;
															assign node20765 = (inp[10]) ? 4'b1010 : node20766;
																assign node20766 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node20771 = (inp[12]) ? node20879 : node20772;
										assign node20772 = (inp[15]) ? node20824 : node20773;
											assign node20773 = (inp[4]) ? node20801 : node20774;
												assign node20774 = (inp[1]) ? node20788 : node20775;
													assign node20775 = (inp[10]) ? node20781 : node20776;
														assign node20776 = (inp[11]) ? 4'b1110 : node20777;
															assign node20777 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node20781 = (inp[9]) ? node20785 : node20782;
															assign node20782 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node20785 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node20788 = (inp[11]) ? node20798 : node20789;
														assign node20789 = (inp[0]) ? 4'b1011 : node20790;
															assign node20790 = (inp[9]) ? node20794 : node20791;
																assign node20791 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node20794 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node20798 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node20801 = (inp[1]) ? node20809 : node20802;
													assign node20802 = (inp[10]) ? node20804 : 4'b1101;
														assign node20804 = (inp[9]) ? node20806 : 4'b1100;
															assign node20806 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node20809 = (inp[0]) ? node20815 : node20810;
														assign node20810 = (inp[9]) ? node20812 : 4'b1100;
															assign node20812 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node20815 = (inp[9]) ? 4'b1101 : node20816;
															assign node20816 = (inp[10]) ? node20820 : node20817;
																assign node20817 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node20820 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node20824 = (inp[0]) ? node20844 : node20825;
												assign node20825 = (inp[4]) ? node20833 : node20826;
													assign node20826 = (inp[1]) ? 4'b1110 : node20827;
														assign node20827 = (inp[10]) ? 4'b1010 : node20828;
															assign node20828 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20833 = (inp[1]) ? node20837 : node20834;
														assign node20834 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node20837 = (inp[11]) ? node20839 : 4'b1011;
															assign node20839 = (inp[10]) ? 4'b1010 : node20840;
																assign node20840 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node20844 = (inp[9]) ? node20862 : node20845;
													assign node20845 = (inp[10]) ? node20855 : node20846;
														assign node20846 = (inp[11]) ? 4'b1011 : node20847;
															assign node20847 = (inp[1]) ? node20851 : node20848;
																assign node20848 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node20851 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node20855 = (inp[1]) ? node20859 : node20856;
															assign node20856 = (inp[11]) ? 4'b1010 : 4'b1110;
															assign node20859 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node20862 = (inp[10]) ? node20872 : node20863;
														assign node20863 = (inp[1]) ? node20867 : node20864;
															assign node20864 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node20867 = (inp[4]) ? node20869 : 4'b1111;
																assign node20869 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20872 = (inp[1]) ? node20876 : node20873;
															assign node20873 = (inp[11]) ? 4'b1011 : 4'b1111;
															assign node20876 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node20879 = (inp[4]) ? node20925 : node20880;
											assign node20880 = (inp[15]) ? node20902 : node20881;
												assign node20881 = (inp[11]) ? node20889 : node20882;
													assign node20882 = (inp[10]) ? 4'b1100 : node20883;
														assign node20883 = (inp[9]) ? 4'b1100 : node20884;
															assign node20884 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node20889 = (inp[0]) ? node20897 : node20890;
														assign node20890 = (inp[9]) ? 4'b1100 : node20891;
															assign node20891 = (inp[10]) ? 4'b1101 : node20892;
																assign node20892 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node20897 = (inp[9]) ? 4'b1101 : node20898;
															assign node20898 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node20902 = (inp[0]) ? node20916 : node20903;
													assign node20903 = (inp[1]) ? node20905 : 4'b1001;
														assign node20905 = (inp[11]) ? node20911 : node20906;
															assign node20906 = (inp[10]) ? 4'b1000 : node20907;
																assign node20907 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node20911 = (inp[10]) ? node20913 : 4'b1001;
																assign node20913 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node20916 = (inp[10]) ? node20918 : 4'b1000;
														assign node20918 = (inp[11]) ? node20922 : node20919;
															assign node20919 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node20922 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node20925 = (inp[15]) ? node20951 : node20926;
												assign node20926 = (inp[9]) ? node20934 : node20927;
													assign node20927 = (inp[10]) ? 4'b1011 : node20928;
														assign node20928 = (inp[11]) ? 4'b1011 : node20929;
															assign node20929 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node20934 = (inp[10]) ? node20940 : node20935;
														assign node20935 = (inp[1]) ? node20937 : 4'b1011;
															assign node20937 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node20940 = (inp[11]) ? node20946 : node20941;
															assign node20941 = (inp[1]) ? node20943 : 4'b1010;
																assign node20943 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node20946 = (inp[1]) ? 4'b1010 : node20947;
																assign node20947 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node20951 = (inp[1]) ? node20961 : node20952;
													assign node20952 = (inp[9]) ? 4'b1001 : node20953;
														assign node20953 = (inp[10]) ? 4'b1000 : node20954;
															assign node20954 = (inp[11]) ? 4'b1001 : node20955;
																assign node20955 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node20961 = (inp[10]) ? node20967 : node20962;
														assign node20962 = (inp[9]) ? 4'b1000 : node20963;
															assign node20963 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node20967 = (inp[9]) ? node20973 : node20968;
															assign node20968 = (inp[11]) ? 4'b1000 : node20969;
																assign node20969 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node20973 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node20976 = (inp[12]) ? node21170 : node20977;
									assign node20977 = (inp[15]) ? node21069 : node20978;
										assign node20978 = (inp[7]) ? node21024 : node20979;
											assign node20979 = (inp[4]) ? node20999 : node20980;
												assign node20980 = (inp[1]) ? node20994 : node20981;
													assign node20981 = (inp[10]) ? node20987 : node20982;
														assign node20982 = (inp[0]) ? 4'b1100 : node20983;
															assign node20983 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node20987 = (inp[11]) ? node20989 : 4'b1101;
															assign node20989 = (inp[9]) ? node20991 : 4'b1100;
																assign node20991 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node20994 = (inp[0]) ? 4'b1000 : node20995;
														assign node20995 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node20999 = (inp[10]) ? node21009 : node21000;
													assign node21000 = (inp[11]) ? node21006 : node21001;
														assign node21001 = (inp[9]) ? 4'b1101 : node21002;
															assign node21002 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node21006 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node21009 = (inp[0]) ? node21019 : node21010;
														assign node21010 = (inp[11]) ? node21012 : 4'b1100;
															assign node21012 = (inp[1]) ? node21016 : node21013;
																assign node21013 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node21016 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node21019 = (inp[11]) ? 4'b1100 : node21020;
															assign node21020 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node21024 = (inp[1]) ? node21042 : node21025;
												assign node21025 = (inp[4]) ? node21035 : node21026;
													assign node21026 = (inp[0]) ? node21028 : 4'b1111;
														assign node21028 = (inp[9]) ? node21032 : node21029;
															assign node21029 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node21032 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node21035 = (inp[11]) ? 4'b1011 : node21036;
														assign node21036 = (inp[0]) ? node21038 : 4'b1011;
															assign node21038 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node21042 = (inp[10]) ? node21052 : node21043;
													assign node21043 = (inp[0]) ? node21045 : 4'b1110;
														assign node21045 = (inp[11]) ? node21049 : node21046;
															assign node21046 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node21049 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node21052 = (inp[4]) ? node21058 : node21053;
														assign node21053 = (inp[9]) ? node21055 : 4'b1111;
															assign node21055 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node21058 = (inp[9]) ? node21064 : node21059;
															assign node21059 = (inp[0]) ? node21061 : 4'b1111;
																assign node21061 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node21064 = (inp[11]) ? node21066 : 4'b1110;
																assign node21066 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node21069 = (inp[7]) ? node21119 : node21070;
											assign node21070 = (inp[4]) ? node21100 : node21071;
												assign node21071 = (inp[1]) ? node21083 : node21072;
													assign node21072 = (inp[10]) ? 4'b1111 : node21073;
														assign node21073 = (inp[0]) ? 4'b1111 : node21074;
															assign node21074 = (inp[9]) ? node21078 : node21075;
																assign node21075 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node21078 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node21083 = (inp[11]) ? node21089 : node21084;
														assign node21084 = (inp[0]) ? 4'b1010 : node21085;
															assign node21085 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node21089 = (inp[10]) ? node21095 : node21090;
															assign node21090 = (inp[0]) ? 4'b1011 : node21091;
																assign node21091 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node21095 = (inp[0]) ? node21097 : 4'b1011;
																assign node21097 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node21100 = (inp[1]) ? node21112 : node21101;
													assign node21101 = (inp[11]) ? node21107 : node21102;
														assign node21102 = (inp[0]) ? 4'b1011 : node21103;
															assign node21103 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node21107 = (inp[9]) ? node21109 : 4'b1010;
															assign node21109 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node21112 = (inp[9]) ? node21116 : node21113;
														assign node21113 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node21116 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node21119 = (inp[10]) ? node21141 : node21120;
												assign node21120 = (inp[4]) ? node21128 : node21121;
													assign node21121 = (inp[1]) ? node21123 : 4'b1101;
														assign node21123 = (inp[9]) ? 4'b1001 : node21124;
															assign node21124 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node21128 = (inp[1]) ? node21134 : node21129;
														assign node21129 = (inp[9]) ? node21131 : 4'b1001;
															assign node21131 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node21134 = (inp[9]) ? node21136 : 4'b1101;
															assign node21136 = (inp[11]) ? node21138 : 4'b1100;
																assign node21138 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node21141 = (inp[0]) ? node21159 : node21142;
													assign node21142 = (inp[1]) ? node21150 : node21143;
														assign node21143 = (inp[4]) ? 4'b1001 : node21144;
															assign node21144 = (inp[9]) ? 4'b1101 : node21145;
																assign node21145 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node21150 = (inp[4]) ? 4'b1100 : node21151;
															assign node21151 = (inp[9]) ? node21155 : node21152;
																assign node21152 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node21155 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node21159 = (inp[4]) ? node21163 : node21160;
														assign node21160 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node21163 = (inp[1]) ? node21165 : 4'b1000;
															assign node21165 = (inp[11]) ? 4'b1101 : node21166;
																assign node21166 = (inp[9]) ? 4'b1101 : 4'b1100;
									assign node21170 = (inp[15]) ? node21266 : node21171;
										assign node21171 = (inp[7]) ? node21221 : node21172;
											assign node21172 = (inp[1]) ? node21202 : node21173;
												assign node21173 = (inp[10]) ? node21185 : node21174;
													assign node21174 = (inp[9]) ? 4'b1101 : node21175;
														assign node21175 = (inp[11]) ? node21177 : 4'b1101;
															assign node21177 = (inp[4]) ? node21181 : node21178;
																assign node21178 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node21181 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node21185 = (inp[11]) ? node21199 : node21186;
														assign node21186 = (inp[9]) ? node21192 : node21187;
															assign node21187 = (inp[4]) ? node21189 : 4'b1101;
																assign node21189 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node21192 = (inp[0]) ? node21196 : node21193;
																assign node21193 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node21196 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node21199 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node21202 = (inp[4]) ? node21214 : node21203;
													assign node21203 = (inp[0]) ? node21209 : node21204;
														assign node21204 = (inp[9]) ? node21206 : 4'b1100;
															assign node21206 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node21209 = (inp[11]) ? 4'b1101 : node21210;
															assign node21210 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node21214 = (inp[9]) ? node21218 : node21215;
														assign node21215 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node21218 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node21221 = (inp[4]) ? node21245 : node21222;
												assign node21222 = (inp[1]) ? node21238 : node21223;
													assign node21223 = (inp[11]) ? node21231 : node21224;
														assign node21224 = (inp[9]) ? node21228 : node21225;
															assign node21225 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node21228 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node21231 = (inp[0]) ? node21235 : node21232;
															assign node21232 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node21235 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node21238 = (inp[0]) ? 4'b1110 : node21239;
														assign node21239 = (inp[11]) ? node21241 : 4'b1111;
															assign node21241 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node21245 = (inp[10]) ? node21253 : node21246;
													assign node21246 = (inp[9]) ? node21248 : 4'b1111;
														assign node21248 = (inp[11]) ? node21250 : 4'b1111;
															assign node21250 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node21253 = (inp[0]) ? node21259 : node21254;
														assign node21254 = (inp[9]) ? 4'b1111 : node21255;
															assign node21255 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node21259 = (inp[1]) ? 4'b1110 : node21260;
															assign node21260 = (inp[9]) ? node21262 : 4'b1111;
																assign node21262 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node21266 = (inp[7]) ? node21290 : node21267;
											assign node21267 = (inp[4]) ? node21281 : node21268;
												assign node21268 = (inp[11]) ? node21274 : node21269;
													assign node21269 = (inp[0]) ? 4'b1111 : node21270;
														assign node21270 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node21274 = (inp[0]) ? node21278 : node21275;
														assign node21275 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node21278 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node21281 = (inp[9]) ? 4'b1110 : node21282;
													assign node21282 = (inp[11]) ? node21286 : node21283;
														assign node21283 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node21286 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node21290 = (inp[1]) ? node21304 : node21291;
												assign node21291 = (inp[0]) ? node21299 : node21292;
													assign node21292 = (inp[4]) ? 4'b1101 : node21293;
														assign node21293 = (inp[11]) ? node21295 : 4'b1100;
															assign node21295 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node21299 = (inp[9]) ? node21301 : 4'b1100;
														assign node21301 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node21304 = (inp[9]) ? node21316 : node21305;
													assign node21305 = (inp[11]) ? node21307 : 4'b1101;
														assign node21307 = (inp[10]) ? node21313 : node21308;
															assign node21308 = (inp[0]) ? node21310 : 4'b1101;
																assign node21310 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node21313 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node21316 = (inp[11]) ? node21322 : node21317;
														assign node21317 = (inp[0]) ? 4'b1100 : node21318;
															assign node21318 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node21322 = (inp[4]) ? 4'b1101 : node21323;
															assign node21323 = (inp[0]) ? 4'b1101 : 4'b1100;
						assign node21327 = (inp[5]) ? node22051 : node21328;
							assign node21328 = (inp[6]) ? node21680 : node21329;
								assign node21329 = (inp[1]) ? node21481 : node21330;
									assign node21330 = (inp[12]) ? node21408 : node21331;
										assign node21331 = (inp[7]) ? node21373 : node21332;
											assign node21332 = (inp[4]) ? node21350 : node21333;
												assign node21333 = (inp[9]) ? node21339 : node21334;
													assign node21334 = (inp[0]) ? node21336 : 4'b1101;
														assign node21336 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node21339 = (inp[11]) ? node21341 : 4'b1100;
														assign node21341 = (inp[0]) ? node21343 : 4'b1100;
															assign node21343 = (inp[10]) ? node21347 : node21344;
																assign node21344 = (inp[15]) ? 4'b1100 : 4'b1101;
																assign node21347 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node21350 = (inp[15]) ? node21364 : node21351;
													assign node21351 = (inp[0]) ? node21359 : node21352;
														assign node21352 = (inp[11]) ? 4'b1111 : node21353;
															assign node21353 = (inp[9]) ? 4'b1110 : node21354;
																assign node21354 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node21359 = (inp[9]) ? node21361 : 4'b1111;
															assign node21361 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node21364 = (inp[0]) ? node21366 : 4'b1001;
														assign node21366 = (inp[11]) ? 4'b1000 : node21367;
															assign node21367 = (inp[10]) ? node21369 : 4'b1001;
																assign node21369 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node21373 = (inp[4]) ? node21395 : node21374;
												assign node21374 = (inp[15]) ? node21382 : node21375;
													assign node21375 = (inp[11]) ? node21377 : 4'b1111;
														assign node21377 = (inp[10]) ? node21379 : 4'b1111;
															assign node21379 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node21382 = (inp[0]) ? node21388 : node21383;
														assign node21383 = (inp[11]) ? 4'b1011 : node21384;
															assign node21384 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node21388 = (inp[9]) ? node21390 : 4'b1010;
															assign node21390 = (inp[11]) ? node21392 : 4'b1011;
																assign node21392 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node21395 = (inp[15]) ? node21399 : node21396;
													assign node21396 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node21399 = (inp[11]) ? 4'b1110 : node21400;
														assign node21400 = (inp[9]) ? node21402 : 4'b1111;
															assign node21402 = (inp[0]) ? node21404 : 4'b1110;
																assign node21404 = (inp[10]) ? 4'b1111 : 4'b1110;
										assign node21408 = (inp[7]) ? node21442 : node21409;
											assign node21409 = (inp[4]) ? node21429 : node21410;
												assign node21410 = (inp[0]) ? node21420 : node21411;
													assign node21411 = (inp[10]) ? 4'b1110 : node21412;
														assign node21412 = (inp[9]) ? node21416 : node21413;
															assign node21413 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node21416 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node21420 = (inp[15]) ? node21426 : node21421;
														assign node21421 = (inp[10]) ? 4'b1111 : node21422;
															assign node21422 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node21426 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node21429 = (inp[15]) ? node21437 : node21430;
													assign node21430 = (inp[10]) ? node21432 : 4'b1000;
														assign node21432 = (inp[9]) ? 4'b1001 : node21433;
															assign node21433 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node21437 = (inp[10]) ? node21439 : 4'b1111;
														assign node21439 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node21442 = (inp[15]) ? node21462 : node21443;
												assign node21443 = (inp[4]) ? node21453 : node21444;
													assign node21444 = (inp[9]) ? node21448 : node21445;
														assign node21445 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node21448 = (inp[10]) ? 4'b1001 : node21449;
															assign node21449 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node21453 = (inp[11]) ? node21455 : 4'b1110;
														assign node21455 = (inp[9]) ? 4'b1111 : node21456;
															assign node21456 = (inp[10]) ? 4'b1110 : node21457;
																assign node21457 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node21462 = (inp[11]) ? node21476 : node21463;
													assign node21463 = (inp[0]) ? node21469 : node21464;
														assign node21464 = (inp[9]) ? 4'b1101 : node21465;
															assign node21465 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node21469 = (inp[9]) ? node21473 : node21470;
															assign node21470 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node21473 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node21476 = (inp[9]) ? node21478 : 4'b1100;
														assign node21478 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node21481 = (inp[12]) ? node21583 : node21482;
										assign node21482 = (inp[7]) ? node21540 : node21483;
											assign node21483 = (inp[4]) ? node21515 : node21484;
												assign node21484 = (inp[11]) ? node21502 : node21485;
													assign node21485 = (inp[15]) ? node21497 : node21486;
														assign node21486 = (inp[0]) ? node21492 : node21487;
															assign node21487 = (inp[9]) ? 4'b1001 : node21488;
																assign node21488 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node21492 = (inp[9]) ? 4'b1000 : node21493;
																assign node21493 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node21497 = (inp[10]) ? 4'b1001 : node21498;
															assign node21498 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node21502 = (inp[15]) ? node21508 : node21503;
														assign node21503 = (inp[10]) ? 4'b1000 : node21504;
															assign node21504 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node21508 = (inp[10]) ? 4'b1001 : node21509;
															assign node21509 = (inp[9]) ? 4'b1000 : node21510;
																assign node21510 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node21515 = (inp[15]) ? node21527 : node21516;
													assign node21516 = (inp[0]) ? node21518 : 4'b1011;
														assign node21518 = (inp[10]) ? 4'b1010 : node21519;
															assign node21519 = (inp[9]) ? node21523 : node21520;
																assign node21520 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node21523 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node21527 = (inp[11]) ? node21533 : node21528;
														assign node21528 = (inp[9]) ? node21530 : 4'b1100;
															assign node21530 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node21533 = (inp[9]) ? node21535 : 4'b1101;
															assign node21535 = (inp[10]) ? node21537 : 4'b1101;
																assign node21537 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node21540 = (inp[15]) ? node21564 : node21541;
												assign node21541 = (inp[4]) ? node21549 : node21542;
													assign node21542 = (inp[10]) ? node21544 : 4'b1110;
														assign node21544 = (inp[9]) ? 4'b1111 : node21545;
															assign node21545 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node21549 = (inp[11]) ? node21557 : node21550;
														assign node21550 = (inp[0]) ? node21552 : 4'b1101;
															assign node21552 = (inp[10]) ? 4'b1101 : node21553;
																assign node21553 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node21557 = (inp[0]) ? node21559 : 4'b1100;
															assign node21559 = (inp[9]) ? 4'b1101 : node21560;
																assign node21560 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node21564 = (inp[4]) ? node21580 : node21565;
													assign node21565 = (inp[11]) ? node21575 : node21566;
														assign node21566 = (inp[9]) ? 4'b1011 : node21567;
															assign node21567 = (inp[0]) ? node21571 : node21568;
																assign node21568 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node21571 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node21575 = (inp[9]) ? 4'b1010 : node21576;
															assign node21576 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node21580 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node21583 = (inp[7]) ? node21623 : node21584;
											assign node21584 = (inp[15]) ? node21602 : node21585;
												assign node21585 = (inp[4]) ? node21593 : node21586;
													assign node21586 = (inp[10]) ? 4'b1011 : node21587;
														assign node21587 = (inp[9]) ? node21589 : 4'b1010;
															assign node21589 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node21593 = (inp[9]) ? 4'b1000 : node21594;
														assign node21594 = (inp[10]) ? node21596 : 4'b1001;
															assign node21596 = (inp[11]) ? node21598 : 4'b1001;
																assign node21598 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node21602 = (inp[9]) ? node21620 : node21603;
													assign node21603 = (inp[0]) ? node21613 : node21604;
														assign node21604 = (inp[10]) ? node21608 : node21605;
															assign node21605 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node21608 = (inp[4]) ? 4'b1011 : node21609;
																assign node21609 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node21613 = (inp[11]) ? node21615 : 4'b1010;
															assign node21615 = (inp[10]) ? node21617 : 4'b1010;
																assign node21617 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node21620 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node21623 = (inp[15]) ? node21651 : node21624;
												assign node21624 = (inp[4]) ? node21636 : node21625;
													assign node21625 = (inp[0]) ? node21627 : 4'b1101;
														assign node21627 = (inp[11]) ? node21633 : node21628;
															assign node21628 = (inp[9]) ? node21630 : 4'b1101;
																assign node21630 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node21633 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node21636 = (inp[11]) ? node21646 : node21637;
														assign node21637 = (inp[10]) ? node21639 : 4'b1010;
															assign node21639 = (inp[9]) ? node21643 : node21640;
																assign node21640 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node21643 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node21646 = (inp[9]) ? 4'b1010 : node21647;
															assign node21647 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node21651 = (inp[4]) ? node21667 : node21652;
													assign node21652 = (inp[11]) ? node21654 : 4'b1000;
														assign node21654 = (inp[10]) ? node21662 : node21655;
															assign node21655 = (inp[0]) ? node21659 : node21656;
																assign node21656 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node21659 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node21662 = (inp[9]) ? 4'b1000 : node21663;
																assign node21663 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node21667 = (inp[11]) ? node21673 : node21668;
														assign node21668 = (inp[0]) ? 4'b1001 : node21669;
															assign node21669 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node21673 = (inp[10]) ? node21677 : node21674;
															assign node21674 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node21677 = (inp[9]) ? 4'b1001 : 4'b1000;
								assign node21680 = (inp[12]) ? node21862 : node21681;
									assign node21681 = (inp[15]) ? node21777 : node21682;
										assign node21682 = (inp[7]) ? node21734 : node21683;
											assign node21683 = (inp[1]) ? node21711 : node21684;
												assign node21684 = (inp[4]) ? node21704 : node21685;
													assign node21685 = (inp[10]) ? node21697 : node21686;
														assign node21686 = (inp[0]) ? node21692 : node21687;
															assign node21687 = (inp[11]) ? node21689 : 4'b1100;
																assign node21689 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node21692 = (inp[9]) ? node21694 : 4'b1100;
																assign node21694 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node21697 = (inp[11]) ? node21701 : node21698;
															assign node21698 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node21701 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node21704 = (inp[9]) ? node21708 : node21705;
														assign node21705 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node21708 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node21711 = (inp[4]) ? node21719 : node21712;
													assign node21712 = (inp[9]) ? 4'b1001 : node21713;
														assign node21713 = (inp[0]) ? node21715 : 4'b1000;
															assign node21715 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node21719 = (inp[0]) ? node21725 : node21720;
														assign node21720 = (inp[11]) ? node21722 : 4'b1100;
															assign node21722 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node21725 = (inp[10]) ? node21727 : 4'b1101;
															assign node21727 = (inp[9]) ? node21731 : node21728;
																assign node21728 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node21731 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node21734 = (inp[1]) ? node21754 : node21735;
												assign node21735 = (inp[4]) ? node21739 : node21736;
													assign node21736 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node21739 = (inp[10]) ? 4'b1010 : node21740;
														assign node21740 = (inp[0]) ? node21748 : node21741;
															assign node21741 = (inp[11]) ? node21745 : node21742;
																assign node21742 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node21745 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node21748 = (inp[9]) ? node21750 : 4'b1011;
																assign node21750 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node21754 = (inp[11]) ? node21766 : node21755;
													assign node21755 = (inp[10]) ? node21761 : node21756;
														assign node21756 = (inp[9]) ? 4'b1110 : node21757;
															assign node21757 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node21761 = (inp[9]) ? node21763 : 4'b1110;
															assign node21763 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node21766 = (inp[4]) ? node21768 : 4'b1111;
														assign node21768 = (inp[10]) ? node21774 : node21769;
															assign node21769 = (inp[0]) ? 4'b1111 : node21770;
																assign node21770 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node21774 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node21777 = (inp[7]) ? node21819 : node21778;
											assign node21778 = (inp[0]) ? node21800 : node21779;
												assign node21779 = (inp[1]) ? node21791 : node21780;
													assign node21780 = (inp[4]) ? node21786 : node21781;
														assign node21781 = (inp[11]) ? node21783 : 4'b1110;
															assign node21783 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node21786 = (inp[11]) ? node21788 : 4'b1010;
															assign node21788 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node21791 = (inp[4]) ? 4'b1111 : node21792;
														assign node21792 = (inp[11]) ? node21796 : node21793;
															assign node21793 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node21796 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node21800 = (inp[1]) ? node21808 : node21801;
													assign node21801 = (inp[4]) ? node21803 : 4'b1111;
														assign node21803 = (inp[11]) ? node21805 : 4'b1011;
															assign node21805 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node21808 = (inp[4]) ? 4'b1110 : node21809;
														assign node21809 = (inp[10]) ? 4'b1011 : node21810;
															assign node21810 = (inp[11]) ? node21814 : node21811;
																assign node21811 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node21814 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node21819 = (inp[4]) ? node21853 : node21820;
												assign node21820 = (inp[1]) ? node21836 : node21821;
													assign node21821 = (inp[0]) ? node21829 : node21822;
														assign node21822 = (inp[9]) ? node21826 : node21823;
															assign node21823 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node21826 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node21829 = (inp[10]) ? node21831 : 4'b1101;
															assign node21831 = (inp[9]) ? 4'b1101 : node21832;
																assign node21832 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node21836 = (inp[0]) ? 4'b1000 : node21837;
														assign node21837 = (inp[10]) ? node21845 : node21838;
															assign node21838 = (inp[11]) ? node21842 : node21839;
																assign node21839 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node21842 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node21845 = (inp[11]) ? node21849 : node21846;
																assign node21846 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node21849 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node21853 = (inp[1]) ? node21855 : 4'b1000;
													assign node21855 = (inp[11]) ? 4'b1100 : node21856;
														assign node21856 = (inp[0]) ? node21858 : 4'b1100;
															assign node21858 = (inp[9]) ? 4'b1101 : 4'b1100;
									assign node21862 = (inp[15]) ? node21964 : node21863;
										assign node21863 = (inp[7]) ? node21909 : node21864;
											assign node21864 = (inp[4]) ? node21892 : node21865;
												assign node21865 = (inp[1]) ? node21873 : node21866;
													assign node21866 = (inp[0]) ? node21868 : 4'b1101;
														assign node21868 = (inp[9]) ? node21870 : 4'b1100;
															assign node21870 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node21873 = (inp[0]) ? node21879 : node21874;
														assign node21874 = (inp[9]) ? 4'b1100 : node21875;
															assign node21875 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node21879 = (inp[10]) ? node21887 : node21880;
															assign node21880 = (inp[11]) ? node21884 : node21881;
																assign node21881 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node21884 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node21887 = (inp[9]) ? 4'b1101 : node21888;
																assign node21888 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node21892 = (inp[1]) ? node21902 : node21893;
													assign node21893 = (inp[0]) ? node21895 : 4'b1100;
														assign node21895 = (inp[9]) ? node21899 : node21896;
															assign node21896 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node21899 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node21902 = (inp[10]) ? node21904 : 4'b1000;
														assign node21904 = (inp[11]) ? 4'b1001 : node21905;
															assign node21905 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node21909 = (inp[1]) ? node21931 : node21910;
												assign node21910 = (inp[4]) ? node21918 : node21911;
													assign node21911 = (inp[9]) ? node21915 : node21912;
														assign node21912 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node21915 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node21918 = (inp[10]) ? node21926 : node21919;
														assign node21919 = (inp[9]) ? node21923 : node21920;
															assign node21920 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node21923 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node21926 = (inp[0]) ? 4'b1111 : node21927;
															assign node21927 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node21931 = (inp[10]) ? node21943 : node21932;
													assign node21932 = (inp[0]) ? node21934 : 4'b1110;
														assign node21934 = (inp[4]) ? 4'b1111 : node21935;
															assign node21935 = (inp[9]) ? node21939 : node21936;
																assign node21936 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node21939 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node21943 = (inp[4]) ? node21949 : node21944;
														assign node21944 = (inp[11]) ? 4'b1111 : node21945;
															assign node21945 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node21949 = (inp[9]) ? node21957 : node21950;
															assign node21950 = (inp[11]) ? node21954 : node21951;
																assign node21951 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node21954 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node21957 = (inp[0]) ? node21961 : node21958;
																assign node21958 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node21961 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node21964 = (inp[7]) ? node22016 : node21965;
											assign node21965 = (inp[4]) ? node21993 : node21966;
												assign node21966 = (inp[10]) ? node21986 : node21967;
													assign node21967 = (inp[0]) ? node21981 : node21968;
														assign node21968 = (inp[1]) ? node21976 : node21969;
															assign node21969 = (inp[9]) ? node21973 : node21970;
																assign node21970 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node21973 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node21976 = (inp[11]) ? 4'b1110 : node21977;
																assign node21977 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node21981 = (inp[1]) ? node21983 : 4'b1111;
															assign node21983 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node21986 = (inp[11]) ? node21990 : node21987;
														assign node21987 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node21990 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node21993 = (inp[0]) ? node22001 : node21994;
													assign node21994 = (inp[11]) ? node21998 : node21995;
														assign node21995 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node21998 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node22001 = (inp[1]) ? node22009 : node22002;
														assign node22002 = (inp[9]) ? node22006 : node22003;
															assign node22003 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node22006 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node22009 = (inp[9]) ? node22013 : node22010;
															assign node22010 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node22013 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node22016 = (inp[4]) ? node22032 : node22017;
												assign node22017 = (inp[1]) ? node22019 : 4'b1100;
													assign node22019 = (inp[10]) ? node22027 : node22020;
														assign node22020 = (inp[11]) ? node22024 : node22021;
															assign node22021 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node22024 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node22027 = (inp[9]) ? 4'b1100 : node22028;
															assign node22028 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node22032 = (inp[1]) ? node22044 : node22033;
													assign node22033 = (inp[11]) ? 4'b1101 : node22034;
														assign node22034 = (inp[10]) ? 4'b1101 : node22035;
															assign node22035 = (inp[0]) ? node22039 : node22036;
																assign node22036 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node22039 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node22044 = (inp[11]) ? 4'b1100 : node22045;
														assign node22045 = (inp[0]) ? 4'b1100 : node22046;
															assign node22046 = (inp[9]) ? 4'b1100 : 4'b1101;
							assign node22051 = (inp[6]) ? node22419 : node22052;
								assign node22052 = (inp[12]) ? node22236 : node22053;
									assign node22053 = (inp[7]) ? node22143 : node22054;
										assign node22054 = (inp[4]) ? node22106 : node22055;
											assign node22055 = (inp[9]) ? node22073 : node22056;
												assign node22056 = (inp[10]) ? node22068 : node22057;
													assign node22057 = (inp[15]) ? node22059 : 4'b1100;
														assign node22059 = (inp[0]) ? 4'b1101 : node22060;
															assign node22060 = (inp[1]) ? node22064 : node22061;
																assign node22061 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node22064 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node22068 = (inp[0]) ? 4'b1101 : node22069;
														assign node22069 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node22073 = (inp[15]) ? node22087 : node22074;
													assign node22074 = (inp[0]) ? node22080 : node22075;
														assign node22075 = (inp[11]) ? node22077 : 4'b1101;
															assign node22077 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node22080 = (inp[10]) ? node22082 : 4'b1100;
															assign node22082 = (inp[1]) ? node22084 : 4'b1100;
																assign node22084 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node22087 = (inp[0]) ? node22101 : node22088;
														assign node22088 = (inp[10]) ? node22096 : node22089;
															assign node22089 = (inp[11]) ? node22093 : node22090;
																assign node22090 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node22093 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node22096 = (inp[1]) ? node22098 : 4'b1100;
																assign node22098 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node22101 = (inp[11]) ? 4'b1101 : node22102;
															assign node22102 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node22106 = (inp[15]) ? node22122 : node22107;
												assign node22107 = (inp[1]) ? node22117 : node22108;
													assign node22108 = (inp[0]) ? 4'b1110 : node22109;
														assign node22109 = (inp[10]) ? node22113 : node22110;
															assign node22110 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node22113 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22117 = (inp[11]) ? node22119 : 4'b1111;
														assign node22119 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node22122 = (inp[1]) ? node22130 : node22123;
													assign node22123 = (inp[11]) ? 4'b1001 : node22124;
														assign node22124 = (inp[0]) ? 4'b1000 : node22125;
															assign node22125 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node22130 = (inp[11]) ? node22136 : node22131;
														assign node22131 = (inp[0]) ? 4'b1001 : node22132;
															assign node22132 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node22136 = (inp[9]) ? node22138 : 4'b1000;
															assign node22138 = (inp[10]) ? node22140 : 4'b1000;
																assign node22140 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node22143 = (inp[15]) ? node22185 : node22144;
											assign node22144 = (inp[4]) ? node22170 : node22145;
												assign node22145 = (inp[1]) ? node22165 : node22146;
													assign node22146 = (inp[0]) ? node22156 : node22147;
														assign node22147 = (inp[11]) ? 4'b1010 : node22148;
															assign node22148 = (inp[10]) ? node22152 : node22149;
																assign node22149 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node22152 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node22156 = (inp[9]) ? 4'b1011 : node22157;
															assign node22157 = (inp[10]) ? node22161 : node22158;
																assign node22158 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node22161 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node22165 = (inp[10]) ? 4'b1111 : node22166;
														assign node22166 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node22170 = (inp[10]) ? node22180 : node22171;
													assign node22171 = (inp[9]) ? node22175 : node22172;
														assign node22172 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node22175 = (inp[0]) ? node22177 : 4'b1000;
															assign node22177 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node22180 = (inp[9]) ? node22182 : 4'b1000;
														assign node22182 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node22185 = (inp[9]) ? node22209 : node22186;
												assign node22186 = (inp[10]) ? node22200 : node22187;
													assign node22187 = (inp[11]) ? node22193 : node22188;
														assign node22188 = (inp[1]) ? 4'b1110 : node22189;
															assign node22189 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node22193 = (inp[1]) ? node22195 : 4'b1010;
															assign node22195 = (inp[4]) ? node22197 : 4'b1010;
																assign node22197 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node22200 = (inp[0]) ? node22202 : 4'b1011;
														assign node22202 = (inp[4]) ? node22206 : node22203;
															assign node22203 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node22206 = (inp[1]) ? 4'b1111 : 4'b1010;
												assign node22209 = (inp[1]) ? node22223 : node22210;
													assign node22210 = (inp[4]) ? 4'b1011 : node22211;
														assign node22211 = (inp[10]) ? node22217 : node22212;
															assign node22212 = (inp[0]) ? node22214 : 4'b1110;
																assign node22214 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node22217 = (inp[0]) ? node22219 : 4'b1111;
																assign node22219 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22223 = (inp[4]) ? node22231 : node22224;
														assign node22224 = (inp[11]) ? 4'b1010 : node22225;
															assign node22225 = (inp[10]) ? 4'b1011 : node22226;
																assign node22226 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node22231 = (inp[11]) ? 4'b1111 : node22232;
															assign node22232 = (inp[10]) ? 4'b1110 : 4'b1111;
									assign node22236 = (inp[7]) ? node22336 : node22237;
										assign node22237 = (inp[15]) ? node22281 : node22238;
											assign node22238 = (inp[4]) ? node22258 : node22239;
												assign node22239 = (inp[9]) ? node22247 : node22240;
													assign node22240 = (inp[0]) ? node22242 : 4'b1111;
														assign node22242 = (inp[10]) ? node22244 : 4'b1110;
															assign node22244 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22247 = (inp[11]) ? 4'b1110 : node22248;
														assign node22248 = (inp[10]) ? node22252 : node22249;
															assign node22249 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node22252 = (inp[1]) ? node22254 : 4'b1110;
																assign node22254 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node22258 = (inp[1]) ? node22276 : node22259;
													assign node22259 = (inp[0]) ? node22271 : node22260;
														assign node22260 = (inp[11]) ? node22266 : node22261;
															assign node22261 = (inp[10]) ? 4'b1101 : node22262;
																assign node22262 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node22266 = (inp[9]) ? node22268 : 4'b1100;
																assign node22268 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node22271 = (inp[9]) ? 4'b1101 : node22272;
															assign node22272 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node22276 = (inp[9]) ? node22278 : 4'b1001;
														assign node22278 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node22281 = (inp[1]) ? node22307 : node22282;
												assign node22282 = (inp[4]) ? node22296 : node22283;
													assign node22283 = (inp[9]) ? node22289 : node22284;
														assign node22284 = (inp[10]) ? node22286 : 4'b1111;
															assign node22286 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node22289 = (inp[11]) ? node22291 : 4'b1110;
															assign node22291 = (inp[10]) ? 4'b1110 : node22292;
																assign node22292 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node22296 = (inp[0]) ? node22300 : node22297;
														assign node22297 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node22300 = (inp[11]) ? 4'b1111 : node22301;
															assign node22301 = (inp[9]) ? node22303 : 4'b1110;
																assign node22303 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node22307 = (inp[10]) ? node22323 : node22308;
													assign node22308 = (inp[9]) ? node22316 : node22309;
														assign node22309 = (inp[4]) ? node22311 : 4'b1111;
															assign node22311 = (inp[0]) ? 4'b1110 : node22312;
																assign node22312 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node22316 = (inp[4]) ? 4'b1111 : node22317;
															assign node22317 = (inp[0]) ? 4'b1110 : node22318;
																assign node22318 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22323 = (inp[9]) ? node22329 : node22324;
														assign node22324 = (inp[4]) ? 4'b1111 : node22325;
															assign node22325 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node22329 = (inp[4]) ? 4'b1110 : node22330;
															assign node22330 = (inp[11]) ? node22332 : 4'b1111;
																assign node22332 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node22336 = (inp[15]) ? node22380 : node22337;
											assign node22337 = (inp[4]) ? node22357 : node22338;
												assign node22338 = (inp[11]) ? node22346 : node22339;
													assign node22339 = (inp[10]) ? 4'b1001 : node22340;
														assign node22340 = (inp[1]) ? 4'b1001 : node22341;
															assign node22341 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node22346 = (inp[0]) ? 4'b1000 : node22347;
														assign node22347 = (inp[10]) ? 4'b1001 : node22348;
															assign node22348 = (inp[9]) ? node22352 : node22349;
																assign node22349 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node22352 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node22357 = (inp[9]) ? node22371 : node22358;
													assign node22358 = (inp[11]) ? node22366 : node22359;
														assign node22359 = (inp[10]) ? node22361 : 4'b1110;
															assign node22361 = (inp[1]) ? 4'b1111 : node22362;
																assign node22362 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node22366 = (inp[10]) ? 4'b1110 : node22367;
															assign node22367 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node22371 = (inp[0]) ? node22373 : 4'b1111;
														assign node22373 = (inp[1]) ? 4'b1111 : node22374;
															assign node22374 = (inp[11]) ? node22376 : 4'b1110;
																assign node22376 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node22380 = (inp[9]) ? node22400 : node22381;
												assign node22381 = (inp[1]) ? node22389 : node22382;
													assign node22382 = (inp[10]) ? 4'b1101 : node22383;
														assign node22383 = (inp[11]) ? node22385 : 4'b1101;
															assign node22385 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node22389 = (inp[10]) ? node22393 : node22390;
														assign node22390 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node22393 = (inp[4]) ? node22395 : 4'b1100;
															assign node22395 = (inp[0]) ? 4'b1101 : node22396;
																assign node22396 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node22400 = (inp[11]) ? node22410 : node22401;
													assign node22401 = (inp[0]) ? 4'b1101 : node22402;
														assign node22402 = (inp[4]) ? node22406 : node22403;
															assign node22403 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node22406 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node22410 = (inp[10]) ? node22412 : 4'b1100;
														assign node22412 = (inp[1]) ? node22414 : 4'b1100;
															assign node22414 = (inp[0]) ? 4'b1101 : node22415;
																assign node22415 = (inp[4]) ? 4'b1101 : 4'b1100;
								assign node22419 = (inp[12]) ? node22617 : node22420;
									assign node22420 = (inp[15]) ? node22534 : node22421;
										assign node22421 = (inp[7]) ? node22483 : node22422;
											assign node22422 = (inp[4]) ? node22450 : node22423;
												assign node22423 = (inp[1]) ? node22437 : node22424;
													assign node22424 = (inp[11]) ? node22432 : node22425;
														assign node22425 = (inp[10]) ? node22429 : node22426;
															assign node22426 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node22429 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node22432 = (inp[10]) ? 4'b1001 : node22433;
															assign node22433 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node22437 = (inp[0]) ? node22443 : node22438;
														assign node22438 = (inp[11]) ? node22440 : 4'b1101;
															assign node22440 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node22443 = (inp[11]) ? node22447 : node22444;
															assign node22444 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node22447 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node22450 = (inp[1]) ? node22460 : node22451;
													assign node22451 = (inp[0]) ? node22457 : node22452;
														assign node22452 = (inp[11]) ? node22454 : 4'b1000;
															assign node22454 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node22457 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node22460 = (inp[10]) ? node22470 : node22461;
														assign node22461 = (inp[11]) ? 4'b1001 : node22462;
															assign node22462 = (inp[9]) ? node22466 : node22463;
																assign node22463 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node22466 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node22470 = (inp[11]) ? node22478 : node22471;
															assign node22471 = (inp[0]) ? node22475 : node22472;
																assign node22472 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node22475 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node22478 = (inp[0]) ? 4'b1000 : node22479;
																assign node22479 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node22483 = (inp[4]) ? node22507 : node22484;
												assign node22484 = (inp[10]) ? node22502 : node22485;
													assign node22485 = (inp[11]) ? node22493 : node22486;
														assign node22486 = (inp[1]) ? 4'b1010 : node22487;
															assign node22487 = (inp[0]) ? node22489 : 4'b1010;
																assign node22489 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node22493 = (inp[9]) ? node22497 : node22494;
															assign node22494 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node22497 = (inp[1]) ? 4'b1010 : node22498;
																assign node22498 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node22502 = (inp[11]) ? 4'b1010 : node22503;
														assign node22503 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node22507 = (inp[1]) ? node22521 : node22508;
													assign node22508 = (inp[10]) ? node22516 : node22509;
														assign node22509 = (inp[0]) ? node22511 : 4'b1111;
															assign node22511 = (inp[11]) ? 4'b1111 : node22512;
																assign node22512 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node22516 = (inp[0]) ? 4'b1110 : node22517;
															assign node22517 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22521 = (inp[11]) ? node22529 : node22522;
														assign node22522 = (inp[10]) ? 4'b1010 : node22523;
															assign node22523 = (inp[9]) ? 4'b1011 : node22524;
																assign node22524 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node22529 = (inp[0]) ? node22531 : 4'b1010;
															assign node22531 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node22534 = (inp[7]) ? node22578 : node22535;
											assign node22535 = (inp[11]) ? node22553 : node22536;
												assign node22536 = (inp[9]) ? node22546 : node22537;
													assign node22537 = (inp[0]) ? 4'b1110 : node22538;
														assign node22538 = (inp[10]) ? 4'b1110 : node22539;
															assign node22539 = (inp[4]) ? 4'b1011 : node22540;
																assign node22540 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node22546 = (inp[1]) ? 4'b1111 : node22547;
														assign node22547 = (inp[4]) ? 4'b1111 : node22548;
															assign node22548 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node22553 = (inp[9]) ? node22569 : node22554;
													assign node22554 = (inp[0]) ? node22562 : node22555;
														assign node22555 = (inp[10]) ? node22557 : 4'b1111;
															assign node22557 = (inp[4]) ? 4'b1010 : node22558;
																assign node22558 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node22562 = (inp[10]) ? 4'b1111 : node22563;
															assign node22563 = (inp[1]) ? node22565 : 4'b1010;
																assign node22565 = (inp[4]) ? 4'b1010 : 4'b1111;
													assign node22569 = (inp[4]) ? node22575 : node22570;
														assign node22570 = (inp[1]) ? 4'b1110 : node22571;
															assign node22571 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node22575 = (inp[1]) ? 4'b1011 : 4'b1110;
											assign node22578 = (inp[1]) ? node22596 : node22579;
												assign node22579 = (inp[4]) ? node22589 : node22580;
													assign node22580 = (inp[0]) ? node22586 : node22581;
														assign node22581 = (inp[9]) ? 4'b1001 : node22582;
															assign node22582 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node22586 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node22589 = (inp[10]) ? 4'b1101 : node22590;
														assign node22590 = (inp[9]) ? node22592 : 4'b1100;
															assign node22592 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node22596 = (inp[4]) ? node22606 : node22597;
													assign node22597 = (inp[9]) ? node22599 : 4'b1101;
														assign node22599 = (inp[10]) ? node22601 : 4'b1101;
															assign node22601 = (inp[0]) ? 4'b1100 : node22602;
																assign node22602 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node22606 = (inp[10]) ? node22608 : 4'b1000;
														assign node22608 = (inp[11]) ? 4'b1000 : node22609;
															assign node22609 = (inp[9]) ? node22613 : node22610;
																assign node22610 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node22613 = (inp[0]) ? 4'b1001 : 4'b1000;
									assign node22617 = (inp[15]) ? node22693 : node22618;
										assign node22618 = (inp[7]) ? node22648 : node22619;
											assign node22619 = (inp[4]) ? node22635 : node22620;
												assign node22620 = (inp[10]) ? node22626 : node22621;
													assign node22621 = (inp[9]) ? node22623 : 4'b1000;
														assign node22623 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node22626 = (inp[0]) ? 4'b1000 : node22627;
														assign node22627 = (inp[11]) ? 4'b1001 : node22628;
															assign node22628 = (inp[9]) ? node22630 : 4'b1000;
																assign node22630 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node22635 = (inp[1]) ? node22641 : node22636;
													assign node22636 = (inp[9]) ? node22638 : 4'b1001;
														assign node22638 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node22641 = (inp[11]) ? node22643 : 4'b1101;
														assign node22643 = (inp[9]) ? node22645 : 4'b1100;
															assign node22645 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node22648 = (inp[4]) ? node22664 : node22649;
												assign node22649 = (inp[1]) ? node22655 : node22650;
													assign node22650 = (inp[10]) ? 4'b1111 : node22651;
														assign node22651 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node22655 = (inp[0]) ? node22657 : 4'b1011;
														assign node22657 = (inp[11]) ? node22661 : node22658;
															assign node22658 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node22661 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node22664 = (inp[10]) ? node22678 : node22665;
													assign node22665 = (inp[1]) ? node22671 : node22666;
														assign node22666 = (inp[11]) ? node22668 : 4'b1011;
															assign node22668 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node22671 = (inp[9]) ? 4'b1010 : node22672;
															assign node22672 = (inp[0]) ? node22674 : 4'b1010;
																assign node22674 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node22678 = (inp[1]) ? node22688 : node22679;
														assign node22679 = (inp[0]) ? node22685 : node22680;
															assign node22680 = (inp[11]) ? node22682 : 4'b1010;
																assign node22682 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node22685 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node22688 = (inp[9]) ? 4'b1011 : node22689;
															assign node22689 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node22693 = (inp[7]) ? node22727 : node22694;
											assign node22694 = (inp[0]) ? node22714 : node22695;
												assign node22695 = (inp[1]) ? node22705 : node22696;
													assign node22696 = (inp[4]) ? 4'b1011 : node22697;
														assign node22697 = (inp[11]) ? node22701 : node22698;
															assign node22698 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node22701 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node22705 = (inp[4]) ? 4'b1010 : node22706;
														assign node22706 = (inp[11]) ? node22710 : node22707;
															assign node22707 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node22710 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node22714 = (inp[11]) ? node22720 : node22715;
													assign node22715 = (inp[4]) ? node22717 : 4'b1011;
														assign node22717 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node22720 = (inp[9]) ? node22724 : node22721;
														assign node22721 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node22724 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node22727 = (inp[4]) ? node22745 : node22728;
												assign node22728 = (inp[1]) ? node22740 : node22729;
													assign node22729 = (inp[9]) ? node22735 : node22730;
														assign node22730 = (inp[0]) ? 4'b1000 : node22731;
															assign node22731 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node22735 = (inp[10]) ? node22737 : 4'b1001;
															assign node22737 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node22740 = (inp[9]) ? node22742 : 4'b1001;
														assign node22742 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node22745 = (inp[0]) ? node22755 : node22746;
													assign node22746 = (inp[10]) ? 4'b1001 : node22747;
														assign node22747 = (inp[11]) ? node22751 : node22748;
															assign node22748 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node22751 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node22755 = (inp[1]) ? 4'b1000 : 4'b1001;
					assign node22758 = (inp[13]) ? node24046 : node22759;
						assign node22759 = (inp[5]) ? node23459 : node22760;
							assign node22760 = (inp[6]) ? node23152 : node22761;
								assign node22761 = (inp[1]) ? node22937 : node22762;
									assign node22762 = (inp[7]) ? node22836 : node22763;
										assign node22763 = (inp[12]) ? node22803 : node22764;
											assign node22764 = (inp[4]) ? node22782 : node22765;
												assign node22765 = (inp[11]) ? node22775 : node22766;
													assign node22766 = (inp[0]) ? 4'b1101 : node22767;
														assign node22767 = (inp[9]) ? node22771 : node22768;
															assign node22768 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node22771 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node22775 = (inp[10]) ? node22779 : node22776;
														assign node22776 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node22779 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node22782 = (inp[15]) ? node22794 : node22783;
													assign node22783 = (inp[0]) ? node22785 : 4'b1111;
														assign node22785 = (inp[9]) ? 4'b1110 : node22786;
															assign node22786 = (inp[10]) ? node22790 : node22787;
																assign node22787 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node22790 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node22794 = (inp[0]) ? node22796 : 4'b1001;
														assign node22796 = (inp[10]) ? node22800 : node22797;
															assign node22797 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node22800 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node22803 = (inp[4]) ? node22819 : node22804;
												assign node22804 = (inp[0]) ? node22810 : node22805;
													assign node22805 = (inp[10]) ? 4'b1111 : node22806;
														assign node22806 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node22810 = (inp[9]) ? node22812 : 4'b1110;
														assign node22812 = (inp[10]) ? node22816 : node22813;
															assign node22813 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node22816 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node22819 = (inp[15]) ? node22827 : node22820;
													assign node22820 = (inp[11]) ? 4'b1001 : node22821;
														assign node22821 = (inp[0]) ? node22823 : 4'b1000;
															assign node22823 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node22827 = (inp[10]) ? node22829 : 4'b1110;
														assign node22829 = (inp[11]) ? node22831 : 4'b1111;
															assign node22831 = (inp[9]) ? 4'b1110 : node22832;
																assign node22832 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node22836 = (inp[12]) ? node22886 : node22837;
											assign node22837 = (inp[15]) ? node22855 : node22838;
												assign node22838 = (inp[4]) ? node22852 : node22839;
													assign node22839 = (inp[11]) ? node22845 : node22840;
														assign node22840 = (inp[9]) ? 4'b1111 : node22841;
															assign node22841 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node22845 = (inp[10]) ? node22849 : node22846;
															assign node22846 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node22849 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node22852 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node22855 = (inp[4]) ? node22875 : node22856;
													assign node22856 = (inp[0]) ? node22870 : node22857;
														assign node22857 = (inp[9]) ? node22863 : node22858;
															assign node22858 = (inp[11]) ? 4'b1011 : node22859;
																assign node22859 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node22863 = (inp[11]) ? node22867 : node22864;
																assign node22864 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node22867 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node22870 = (inp[9]) ? node22872 : 4'b1010;
															assign node22872 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node22875 = (inp[10]) ? node22881 : node22876;
														assign node22876 = (inp[11]) ? 4'b1111 : node22877;
															assign node22877 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node22881 = (inp[0]) ? node22883 : 4'b1110;
															assign node22883 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node22886 = (inp[15]) ? node22906 : node22887;
												assign node22887 = (inp[4]) ? node22897 : node22888;
													assign node22888 = (inp[11]) ? node22890 : 4'b1000;
														assign node22890 = (inp[9]) ? node22894 : node22891;
															assign node22891 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node22894 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node22897 = (inp[10]) ? 4'b1110 : node22898;
														assign node22898 = (inp[11]) ? node22902 : node22899;
															assign node22899 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node22902 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node22906 = (inp[11]) ? node22922 : node22907;
													assign node22907 = (inp[0]) ? node22909 : 4'b1100;
														assign node22909 = (inp[4]) ? node22917 : node22910;
															assign node22910 = (inp[10]) ? node22914 : node22911;
																assign node22911 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node22914 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node22917 = (inp[9]) ? node22919 : 4'b1100;
																assign node22919 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node22922 = (inp[0]) ? node22930 : node22923;
														assign node22923 = (inp[10]) ? node22927 : node22924;
															assign node22924 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node22927 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node22930 = (inp[10]) ? node22932 : 4'b1101;
															assign node22932 = (inp[9]) ? 4'b1101 : node22933;
																assign node22933 = (inp[4]) ? 4'b1101 : 4'b1100;
									assign node22937 = (inp[7]) ? node23041 : node22938;
										assign node22938 = (inp[12]) ? node22996 : node22939;
											assign node22939 = (inp[4]) ? node22973 : node22940;
												assign node22940 = (inp[11]) ? node22954 : node22941;
													assign node22941 = (inp[15]) ? node22947 : node22942;
														assign node22942 = (inp[9]) ? node22944 : 4'b1000;
															assign node22944 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node22947 = (inp[10]) ? node22949 : 4'b1000;
															assign node22949 = (inp[0]) ? node22951 : 4'b1001;
																assign node22951 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node22954 = (inp[10]) ? node22964 : node22955;
														assign node22955 = (inp[15]) ? 4'b1001 : node22956;
															assign node22956 = (inp[9]) ? node22960 : node22957;
																assign node22957 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node22960 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node22964 = (inp[15]) ? node22970 : node22965;
															assign node22965 = (inp[9]) ? node22967 : 4'b1001;
																assign node22967 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node22970 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node22973 = (inp[15]) ? node22985 : node22974;
													assign node22974 = (inp[0]) ? node22980 : node22975;
														assign node22975 = (inp[9]) ? 4'b1010 : node22976;
															assign node22976 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node22980 = (inp[9]) ? 4'b1011 : node22981;
															assign node22981 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node22985 = (inp[9]) ? node22987 : 4'b1100;
														assign node22987 = (inp[11]) ? 4'b1100 : node22988;
															assign node22988 = (inp[10]) ? node22992 : node22989;
																assign node22989 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node22992 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node22996 = (inp[4]) ? node23022 : node22997;
												assign node22997 = (inp[9]) ? node23007 : node22998;
													assign node22998 = (inp[15]) ? node23002 : node22999;
														assign node22999 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node23002 = (inp[10]) ? node23004 : 4'b1010;
															assign node23004 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node23007 = (inp[11]) ? node23017 : node23008;
														assign node23008 = (inp[0]) ? 4'b1011 : node23009;
															assign node23009 = (inp[15]) ? node23013 : node23010;
																assign node23010 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node23013 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node23017 = (inp[15]) ? 4'b1011 : node23018;
															assign node23018 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node23022 = (inp[15]) ? node23034 : node23023;
													assign node23023 = (inp[9]) ? node23029 : node23024;
														assign node23024 = (inp[10]) ? 4'b1000 : node23025;
															assign node23025 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node23029 = (inp[10]) ? 4'b1001 : node23030;
															assign node23030 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node23034 = (inp[9]) ? 4'b1011 : node23035;
														assign node23035 = (inp[0]) ? 4'b1010 : node23036;
															assign node23036 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node23041 = (inp[12]) ? node23099 : node23042;
											assign node23042 = (inp[4]) ? node23076 : node23043;
												assign node23043 = (inp[15]) ? node23061 : node23044;
													assign node23044 = (inp[11]) ? node23050 : node23045;
														assign node23045 = (inp[9]) ? node23047 : 4'b1111;
															assign node23047 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node23050 = (inp[10]) ? node23056 : node23051;
															assign node23051 = (inp[0]) ? 4'b1110 : node23052;
																assign node23052 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node23056 = (inp[0]) ? 4'b1111 : node23057;
																assign node23057 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node23061 = (inp[0]) ? node23071 : node23062;
														assign node23062 = (inp[11]) ? 4'b1010 : node23063;
															assign node23063 = (inp[9]) ? node23067 : node23064;
																assign node23064 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node23067 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node23071 = (inp[11]) ? 4'b1011 : node23072;
															assign node23072 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node23076 = (inp[15]) ? node23088 : node23077;
													assign node23077 = (inp[11]) ? node23079 : 4'b1100;
														assign node23079 = (inp[0]) ? 4'b1101 : node23080;
															assign node23080 = (inp[9]) ? node23084 : node23081;
																assign node23081 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node23084 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node23088 = (inp[9]) ? node23090 : 4'b1110;
														assign node23090 = (inp[0]) ? node23096 : node23091;
															assign node23091 = (inp[11]) ? node23093 : 4'b1110;
																assign node23093 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node23096 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node23099 = (inp[4]) ? node23125 : node23100;
												assign node23100 = (inp[15]) ? node23116 : node23101;
													assign node23101 = (inp[10]) ? node23105 : node23102;
														assign node23102 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node23105 = (inp[9]) ? node23111 : node23106;
															assign node23106 = (inp[11]) ? 4'b1101 : node23107;
																assign node23107 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node23111 = (inp[0]) ? node23113 : 4'b1100;
																assign node23113 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23116 = (inp[0]) ? node23118 : 4'b1001;
														assign node23118 = (inp[9]) ? node23122 : node23119;
															assign node23119 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node23122 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node23125 = (inp[15]) ? node23141 : node23126;
													assign node23126 = (inp[10]) ? node23136 : node23127;
														assign node23127 = (inp[9]) ? node23131 : node23128;
															assign node23128 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node23131 = (inp[11]) ? node23133 : 4'b1010;
																assign node23133 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node23136 = (inp[0]) ? node23138 : 4'b1010;
															assign node23138 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node23141 = (inp[9]) ? node23149 : node23142;
														assign node23142 = (inp[10]) ? node23144 : 4'b1000;
															assign node23144 = (inp[11]) ? node23146 : 4'b1001;
																assign node23146 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node23149 = (inp[10]) ? 4'b1000 : 4'b1001;
								assign node23152 = (inp[12]) ? node23320 : node23153;
									assign node23153 = (inp[15]) ? node23229 : node23154;
										assign node23154 = (inp[7]) ? node23194 : node23155;
											assign node23155 = (inp[1]) ? node23169 : node23156;
												assign node23156 = (inp[11]) ? node23162 : node23157;
													assign node23157 = (inp[4]) ? node23159 : 4'b1001;
														assign node23159 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node23162 = (inp[4]) ? node23166 : node23163;
														assign node23163 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node23166 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node23169 = (inp[4]) ? node23181 : node23170;
													assign node23170 = (inp[10]) ? node23176 : node23171;
														assign node23171 = (inp[9]) ? 4'b1100 : node23172;
															assign node23172 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node23176 = (inp[0]) ? 4'b1101 : node23177;
															assign node23177 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node23181 = (inp[11]) ? node23189 : node23182;
														assign node23182 = (inp[9]) ? node23186 : node23183;
															assign node23183 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node23186 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node23189 = (inp[9]) ? node23191 : 4'b1000;
															assign node23191 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node23194 = (inp[1]) ? node23208 : node23195;
												assign node23195 = (inp[4]) ? node23203 : node23196;
													assign node23196 = (inp[10]) ? 4'b1011 : node23197;
														assign node23197 = (inp[11]) ? node23199 : 4'b1011;
															assign node23199 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node23203 = (inp[9]) ? node23205 : 4'b1110;
														assign node23205 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node23208 = (inp[0]) ? node23226 : node23209;
													assign node23209 = (inp[9]) ? node23219 : node23210;
														assign node23210 = (inp[10]) ? 4'b1011 : node23211;
															assign node23211 = (inp[11]) ? node23215 : node23212;
																assign node23212 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node23215 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node23219 = (inp[10]) ? node23221 : 4'b1011;
															assign node23221 = (inp[4]) ? node23223 : 4'b1010;
																assign node23223 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node23226 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node23229 = (inp[7]) ? node23279 : node23230;
											assign node23230 = (inp[9]) ? node23250 : node23231;
												assign node23231 = (inp[1]) ? node23239 : node23232;
													assign node23232 = (inp[4]) ? node23236 : node23233;
														assign node23233 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node23236 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node23239 = (inp[4]) ? 4'b1011 : node23240;
														assign node23240 = (inp[10]) ? node23244 : node23241;
															assign node23241 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node23244 = (inp[11]) ? node23246 : 4'b1111;
																assign node23246 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node23250 = (inp[11]) ? node23266 : node23251;
													assign node23251 = (inp[0]) ? node23263 : node23252;
														assign node23252 = (inp[10]) ? node23258 : node23253;
															assign node23253 = (inp[4]) ? 4'b1110 : node23254;
																assign node23254 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node23258 = (inp[4]) ? node23260 : 4'b1110;
																assign node23260 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node23263 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node23266 = (inp[10]) ? node23272 : node23267;
														assign node23267 = (inp[4]) ? 4'b1010 : node23268;
															assign node23268 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node23272 = (inp[1]) ? node23276 : node23273;
															assign node23273 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node23276 = (inp[4]) ? 4'b1010 : 4'b1111;
											assign node23279 = (inp[10]) ? node23299 : node23280;
												assign node23280 = (inp[1]) ? node23290 : node23281;
													assign node23281 = (inp[4]) ? node23283 : 4'b1001;
														assign node23283 = (inp[0]) ? node23285 : 4'b1101;
															assign node23285 = (inp[11]) ? node23287 : 4'b1100;
																assign node23287 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node23290 = (inp[4]) ? node23292 : 4'b1100;
														assign node23292 = (inp[9]) ? node23294 : 4'b1001;
															assign node23294 = (inp[11]) ? 4'b1001 : node23295;
																assign node23295 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node23299 = (inp[4]) ? node23313 : node23300;
													assign node23300 = (inp[1]) ? node23306 : node23301;
														assign node23301 = (inp[11]) ? node23303 : 4'b1001;
															assign node23303 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node23306 = (inp[9]) ? node23310 : node23307;
															assign node23307 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node23310 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node23313 = (inp[1]) ? 4'b1000 : node23314;
														assign node23314 = (inp[11]) ? node23316 : 4'b1100;
															assign node23316 = (inp[9]) ? 4'b1101 : 4'b1100;
									assign node23320 = (inp[15]) ? node23416 : node23321;
										assign node23321 = (inp[7]) ? node23367 : node23322;
											assign node23322 = (inp[1]) ? node23346 : node23323;
												assign node23323 = (inp[9]) ? node23335 : node23324;
													assign node23324 = (inp[10]) ? node23326 : 4'b1001;
														assign node23326 = (inp[4]) ? node23328 : 4'b1000;
															assign node23328 = (inp[11]) ? node23332 : node23329;
																assign node23329 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node23332 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node23335 = (inp[11]) ? node23341 : node23336;
														assign node23336 = (inp[0]) ? node23338 : 4'b1001;
															assign node23338 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node23341 = (inp[10]) ? node23343 : 4'b1000;
															assign node23343 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node23346 = (inp[4]) ? node23362 : node23347;
													assign node23347 = (inp[10]) ? node23353 : node23348;
														assign node23348 = (inp[9]) ? 4'b1000 : node23349;
															assign node23349 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node23353 = (inp[9]) ? 4'b1001 : node23354;
															assign node23354 = (inp[0]) ? node23358 : node23355;
																assign node23355 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node23358 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node23362 = (inp[9]) ? 4'b1101 : node23363;
														assign node23363 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node23367 = (inp[1]) ? node23387 : node23368;
												assign node23368 = (inp[4]) ? node23380 : node23369;
													assign node23369 = (inp[10]) ? 4'b1110 : node23370;
														assign node23370 = (inp[9]) ? 4'b1110 : node23371;
															assign node23371 = (inp[11]) ? node23375 : node23372;
																assign node23372 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node23375 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node23380 = (inp[0]) ? 4'b1011 : node23381;
														assign node23381 = (inp[11]) ? 4'b1011 : node23382;
															assign node23382 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node23387 = (inp[10]) ? node23399 : node23388;
													assign node23388 = (inp[4]) ? node23394 : node23389;
														assign node23389 = (inp[0]) ? node23391 : 4'b1010;
															assign node23391 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node23394 = (inp[0]) ? 4'b1010 : node23395;
															assign node23395 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node23399 = (inp[9]) ? node23411 : node23400;
														assign node23400 = (inp[11]) ? node23406 : node23401;
															assign node23401 = (inp[0]) ? node23403 : 4'b1010;
																assign node23403 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node23406 = (inp[4]) ? node23408 : 4'b1011;
																assign node23408 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node23411 = (inp[11]) ? node23413 : 4'b1011;
															assign node23413 = (inp[4]) ? 4'b1011 : 4'b1010;
										assign node23416 = (inp[7]) ? node23436 : node23417;
											assign node23417 = (inp[9]) ? node23431 : node23418;
												assign node23418 = (inp[0]) ? node23420 : 4'b1010;
													assign node23420 = (inp[10]) ? node23426 : node23421;
														assign node23421 = (inp[4]) ? node23423 : 4'b1011;
															assign node23423 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node23426 = (inp[4]) ? node23428 : 4'b1010;
															assign node23428 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node23431 = (inp[11]) ? node23433 : 4'b1011;
													assign node23433 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node23436 = (inp[11]) ? node23448 : node23437;
												assign node23437 = (inp[9]) ? node23443 : node23438;
													assign node23438 = (inp[0]) ? node23440 : 4'b1001;
														assign node23440 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node23443 = (inp[4]) ? node23445 : 4'b1000;
														assign node23445 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node23448 = (inp[9]) ? node23454 : node23449;
													assign node23449 = (inp[4]) ? node23451 : 4'b1000;
														assign node23451 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node23454 = (inp[4]) ? node23456 : 4'b1001;
														assign node23456 = (inp[1]) ? 4'b1001 : 4'b1000;
							assign node23459 = (inp[12]) ? node23811 : node23460;
								assign node23460 = (inp[7]) ? node23630 : node23461;
									assign node23461 = (inp[15]) ? node23555 : node23462;
										assign node23462 = (inp[6]) ? node23510 : node23463;
											assign node23463 = (inp[4]) ? node23491 : node23464;
												assign node23464 = (inp[0]) ? node23472 : node23465;
													assign node23465 = (inp[1]) ? node23469 : node23466;
														assign node23466 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node23469 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node23472 = (inp[1]) ? node23486 : node23473;
														assign node23473 = (inp[10]) ? node23479 : node23474;
															assign node23474 = (inp[9]) ? 4'b1101 : node23475;
																assign node23475 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node23479 = (inp[9]) ? node23483 : node23480;
																assign node23480 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node23483 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node23486 = (inp[9]) ? node23488 : 4'b1101;
															assign node23488 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node23491 = (inp[0]) ? node23501 : node23492;
													assign node23492 = (inp[10]) ? node23498 : node23493;
														assign node23493 = (inp[9]) ? node23495 : 4'b1110;
															assign node23495 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node23498 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node23501 = (inp[1]) ? 4'b1111 : node23502;
														assign node23502 = (inp[11]) ? node23504 : 4'b1110;
															assign node23504 = (inp[9]) ? node23506 : 4'b1111;
																assign node23506 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node23510 = (inp[4]) ? node23534 : node23511;
												assign node23511 = (inp[1]) ? node23521 : node23512;
													assign node23512 = (inp[10]) ? 4'b1100 : node23513;
														assign node23513 = (inp[9]) ? node23517 : node23514;
															assign node23514 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node23517 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23521 = (inp[10]) ? 4'b1001 : node23522;
														assign node23522 = (inp[0]) ? node23528 : node23523;
															assign node23523 = (inp[11]) ? 4'b1000 : node23524;
																assign node23524 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node23528 = (inp[9]) ? 4'b1001 : node23529;
																assign node23529 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node23534 = (inp[9]) ? node23546 : node23535;
													assign node23535 = (inp[11]) ? node23541 : node23536;
														assign node23536 = (inp[1]) ? 4'b1100 : node23537;
															assign node23537 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node23541 = (inp[1]) ? 4'b1101 : node23542;
															assign node23542 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node23546 = (inp[11]) ? node23550 : node23547;
														assign node23547 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node23550 = (inp[1]) ? 4'b1100 : node23551;
															assign node23551 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node23555 = (inp[6]) ? node23593 : node23556;
											assign node23556 = (inp[4]) ? node23574 : node23557;
												assign node23557 = (inp[11]) ? node23569 : node23558;
													assign node23558 = (inp[9]) ? node23564 : node23559;
														assign node23559 = (inp[10]) ? 4'b1101 : node23560;
															assign node23560 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node23564 = (inp[0]) ? 4'b1101 : node23565;
															assign node23565 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node23569 = (inp[10]) ? node23571 : 4'b1100;
														assign node23571 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node23574 = (inp[1]) ? node23582 : node23575;
													assign node23575 = (inp[10]) ? 4'b1000 : node23576;
														assign node23576 = (inp[9]) ? node23578 : 4'b1000;
															assign node23578 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node23582 = (inp[11]) ? 4'b1001 : node23583;
														assign node23583 = (inp[0]) ? 4'b1000 : node23584;
															assign node23584 = (inp[9]) ? node23588 : node23585;
																assign node23585 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node23588 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node23593 = (inp[10]) ? node23611 : node23594;
												assign node23594 = (inp[1]) ? node23608 : node23595;
													assign node23595 = (inp[4]) ? node23599 : node23596;
														assign node23596 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node23599 = (inp[0]) ? node23601 : 4'b1011;
															assign node23601 = (inp[11]) ? node23605 : node23602;
																assign node23602 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node23605 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node23608 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node23611 = (inp[1]) ? node23623 : node23612;
													assign node23612 = (inp[4]) ? node23616 : node23613;
														assign node23613 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node23616 = (inp[9]) ? node23620 : node23617;
															assign node23617 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node23620 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node23623 = (inp[4]) ? node23625 : 4'b1010;
														assign node23625 = (inp[0]) ? node23627 : 4'b1110;
															assign node23627 = (inp[9]) ? 4'b1111 : 4'b1110;
									assign node23630 = (inp[4]) ? node23720 : node23631;
										assign node23631 = (inp[15]) ? node23675 : node23632;
											assign node23632 = (inp[6]) ? node23652 : node23633;
												assign node23633 = (inp[1]) ? node23643 : node23634;
													assign node23634 = (inp[0]) ? 4'b1010 : node23635;
														assign node23635 = (inp[11]) ? 4'b1011 : node23636;
															assign node23636 = (inp[10]) ? node23638 : 4'b1011;
																assign node23638 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node23643 = (inp[9]) ? node23645 : 4'b1111;
														assign node23645 = (inp[11]) ? node23647 : 4'b1110;
															assign node23647 = (inp[10]) ? node23649 : 4'b1111;
																assign node23649 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node23652 = (inp[1]) ? node23662 : node23653;
													assign node23653 = (inp[10]) ? node23657 : node23654;
														assign node23654 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node23657 = (inp[11]) ? node23659 : 4'b1110;
															assign node23659 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node23662 = (inp[0]) ? node23668 : node23663;
														assign node23663 = (inp[9]) ? 4'b1110 : node23664;
															assign node23664 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node23668 = (inp[11]) ? node23672 : node23669;
															assign node23669 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node23672 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node23675 = (inp[6]) ? node23701 : node23676;
												assign node23676 = (inp[1]) ? node23690 : node23677;
													assign node23677 = (inp[11]) ? node23683 : node23678;
														assign node23678 = (inp[10]) ? 4'b1110 : node23679;
															assign node23679 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node23683 = (inp[9]) ? 4'b1111 : node23684;
															assign node23684 = (inp[0]) ? 4'b1110 : node23685;
																assign node23685 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node23690 = (inp[9]) ? node23692 : 4'b1011;
														assign node23692 = (inp[11]) ? node23694 : 4'b1010;
															assign node23694 = (inp[10]) ? node23698 : node23695;
																assign node23695 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node23698 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node23701 = (inp[1]) ? node23713 : node23702;
													assign node23702 = (inp[10]) ? node23708 : node23703;
														assign node23703 = (inp[11]) ? 4'b1101 : node23704;
															assign node23704 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node23708 = (inp[9]) ? 4'b1100 : node23709;
															assign node23709 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23713 = (inp[9]) ? 4'b1000 : node23714;
														assign node23714 = (inp[0]) ? 4'b1001 : node23715;
															assign node23715 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node23720 = (inp[1]) ? node23770 : node23721;
											assign node23721 = (inp[0]) ? node23743 : node23722;
												assign node23722 = (inp[9]) ? node23734 : node23723;
													assign node23723 = (inp[15]) ? node23727 : node23724;
														assign node23724 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node23727 = (inp[6]) ? 4'b1000 : node23728;
															assign node23728 = (inp[11]) ? node23730 : 4'b1010;
																assign node23730 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node23734 = (inp[11]) ? node23736 : 4'b1001;
														assign node23736 = (inp[15]) ? 4'b1000 : node23737;
															assign node23737 = (inp[6]) ? 4'b1011 : node23738;
																assign node23738 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node23743 = (inp[15]) ? node23755 : node23744;
													assign node23744 = (inp[6]) ? node23750 : node23745;
														assign node23745 = (inp[10]) ? node23747 : 4'b1001;
															assign node23747 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node23750 = (inp[11]) ? 4'b1010 : node23751;
															assign node23751 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node23755 = (inp[6]) ? node23761 : node23756;
														assign node23756 = (inp[9]) ? node23758 : 4'b1011;
															assign node23758 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node23761 = (inp[10]) ? node23763 : 4'b1001;
															assign node23763 = (inp[9]) ? node23767 : node23764;
																assign node23764 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node23767 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node23770 = (inp[15]) ? node23786 : node23771;
												assign node23771 = (inp[6]) ? node23779 : node23772;
													assign node23772 = (inp[9]) ? node23774 : 4'b1000;
														assign node23774 = (inp[11]) ? 4'b1001 : node23775;
															assign node23775 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node23779 = (inp[0]) ? node23781 : 4'b1110;
														assign node23781 = (inp[9]) ? 4'b1111 : node23782;
															assign node23782 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node23786 = (inp[6]) ? node23800 : node23787;
													assign node23787 = (inp[9]) ? node23795 : node23788;
														assign node23788 = (inp[11]) ? 4'b1110 : node23789;
															assign node23789 = (inp[10]) ? node23791 : 4'b1111;
																assign node23791 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node23795 = (inp[11]) ? 4'b1111 : node23796;
															assign node23796 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node23800 = (inp[10]) ? node23806 : node23801;
														assign node23801 = (inp[0]) ? 4'b1101 : node23802;
															assign node23802 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node23806 = (inp[9]) ? 4'b1100 : node23807;
															assign node23807 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node23811 = (inp[15]) ? node23969 : node23812;
									assign node23812 = (inp[7]) ? node23898 : node23813;
										assign node23813 = (inp[4]) ? node23859 : node23814;
											assign node23814 = (inp[6]) ? node23832 : node23815;
												assign node23815 = (inp[11]) ? node23823 : node23816;
													assign node23816 = (inp[9]) ? 4'b1110 : node23817;
														assign node23817 = (inp[0]) ? 4'b1111 : node23818;
															assign node23818 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node23823 = (inp[1]) ? 4'b1111 : node23824;
														assign node23824 = (inp[0]) ? node23826 : 4'b1110;
															assign node23826 = (inp[10]) ? node23828 : 4'b1111;
																assign node23828 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node23832 = (inp[1]) ? node23842 : node23833;
													assign node23833 = (inp[10]) ? node23835 : 4'b1101;
														assign node23835 = (inp[9]) ? node23839 : node23836;
															assign node23836 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node23839 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23842 = (inp[10]) ? node23850 : node23843;
														assign node23843 = (inp[11]) ? node23845 : 4'b1100;
															assign node23845 = (inp[9]) ? 4'b1100 : node23846;
																assign node23846 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node23850 = (inp[11]) ? 4'b1101 : node23851;
															assign node23851 = (inp[9]) ? node23855 : node23852;
																assign node23852 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node23855 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node23859 = (inp[1]) ? node23877 : node23860;
												assign node23860 = (inp[9]) ? node23868 : node23861;
													assign node23861 = (inp[0]) ? node23863 : 4'b1101;
														assign node23863 = (inp[6]) ? 4'b1101 : node23864;
															assign node23864 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23868 = (inp[0]) ? node23870 : 4'b1100;
														assign node23870 = (inp[11]) ? node23872 : 4'b1101;
															assign node23872 = (inp[10]) ? 4'b1100 : node23873;
																assign node23873 = (inp[6]) ? 4'b1100 : 4'b1101;
												assign node23877 = (inp[0]) ? node23887 : node23878;
													assign node23878 = (inp[9]) ? 4'b1000 : node23879;
														assign node23879 = (inp[6]) ? 4'b1001 : node23880;
															assign node23880 = (inp[11]) ? 4'b1000 : node23881;
																assign node23881 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node23887 = (inp[6]) ? node23893 : node23888;
														assign node23888 = (inp[10]) ? node23890 : 4'b1001;
															assign node23890 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node23893 = (inp[9]) ? node23895 : 4'b1000;
															assign node23895 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node23898 = (inp[4]) ? node23936 : node23899;
											assign node23899 = (inp[6]) ? node23923 : node23900;
												assign node23900 = (inp[0]) ? node23908 : node23901;
													assign node23901 = (inp[9]) ? node23903 : 4'b1001;
														assign node23903 = (inp[1]) ? 4'b1000 : node23904;
															assign node23904 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node23908 = (inp[10]) ? node23918 : node23909;
														assign node23909 = (inp[1]) ? node23915 : node23910;
															assign node23910 = (inp[9]) ? node23912 : 4'b1000;
																assign node23912 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node23915 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node23918 = (inp[9]) ? node23920 : 4'b1000;
															assign node23920 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node23923 = (inp[1]) ? node23929 : node23924;
													assign node23924 = (inp[11]) ? node23926 : 4'b1010;
														assign node23926 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node23929 = (inp[9]) ? node23933 : node23930;
														assign node23930 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node23933 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node23936 = (inp[10]) ? node23952 : node23937;
												assign node23937 = (inp[9]) ? node23943 : node23938;
													assign node23938 = (inp[6]) ? node23940 : 4'b1111;
														assign node23940 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node23943 = (inp[1]) ? node23945 : 4'b1110;
														assign node23945 = (inp[0]) ? node23949 : node23946;
															assign node23946 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node23949 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node23952 = (inp[6]) ? node23958 : node23953;
													assign node23953 = (inp[9]) ? node23955 : 4'b1110;
														assign node23955 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node23958 = (inp[11]) ? node23964 : node23959;
														assign node23959 = (inp[0]) ? 4'b1110 : node23960;
															assign node23960 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node23964 = (inp[0]) ? node23966 : 4'b1111;
															assign node23966 = (inp[9]) ? 4'b1111 : 4'b1110;
									assign node23969 = (inp[7]) ? node24007 : node23970;
										assign node23970 = (inp[11]) ? node23996 : node23971;
											assign node23971 = (inp[9]) ? node23983 : node23972;
												assign node23972 = (inp[6]) ? 4'b1110 : node23973;
													assign node23973 = (inp[4]) ? node23979 : node23974;
														assign node23974 = (inp[0]) ? 4'b1110 : node23975;
															assign node23975 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node23979 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node23983 = (inp[6]) ? 4'b1111 : node23984;
													assign node23984 = (inp[4]) ? 4'b1110 : node23985;
														assign node23985 = (inp[1]) ? 4'b1111 : node23986;
															assign node23986 = (inp[10]) ? node23990 : node23987;
																assign node23987 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node23990 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node23996 = (inp[9]) ? node24002 : node23997;
												assign node23997 = (inp[6]) ? 4'b1111 : node23998;
													assign node23998 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node24002 = (inp[10]) ? 4'b1110 : node24003;
													assign node24003 = (inp[6]) ? 4'b1110 : 4'b1111;
										assign node24007 = (inp[9]) ? node24023 : node24008;
											assign node24008 = (inp[11]) ? node24018 : node24009;
												assign node24009 = (inp[6]) ? 4'b1100 : node24010;
													assign node24010 = (inp[1]) ? 4'b1101 : node24011;
														assign node24011 = (inp[10]) ? 4'b1100 : node24012;
															assign node24012 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node24018 = (inp[10]) ? 4'b1101 : node24019;
													assign node24019 = (inp[6]) ? 4'b1101 : 4'b1100;
											assign node24023 = (inp[11]) ? node24041 : node24024;
												assign node24024 = (inp[6]) ? 4'b1101 : node24025;
													assign node24025 = (inp[1]) ? node24031 : node24026;
														assign node24026 = (inp[10]) ? 4'b1101 : node24027;
															assign node24027 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node24031 = (inp[4]) ? node24037 : node24032;
															assign node24032 = (inp[10]) ? node24034 : 4'b1100;
																assign node24034 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node24037 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node24041 = (inp[10]) ? 4'b1100 : node24042;
													assign node24042 = (inp[6]) ? 4'b1100 : 4'b1101;
						assign node24046 = (inp[5]) ? node24720 : node24047;
							assign node24047 = (inp[6]) ? node24431 : node24048;
								assign node24048 = (inp[1]) ? node24236 : node24049;
									assign node24049 = (inp[7]) ? node24147 : node24050;
										assign node24050 = (inp[12]) ? node24094 : node24051;
											assign node24051 = (inp[4]) ? node24073 : node24052;
												assign node24052 = (inp[9]) ? node24060 : node24053;
													assign node24053 = (inp[15]) ? 4'b1000 : node24054;
														assign node24054 = (inp[10]) ? 4'b1000 : node24055;
															assign node24055 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node24060 = (inp[15]) ? node24068 : node24061;
														assign node24061 = (inp[10]) ? 4'b1001 : node24062;
															assign node24062 = (inp[0]) ? node24064 : 4'b1000;
																assign node24064 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node24068 = (inp[0]) ? node24070 : 4'b1001;
															assign node24070 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node24073 = (inp[15]) ? node24083 : node24074;
													assign node24074 = (inp[11]) ? node24078 : node24075;
														assign node24075 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node24078 = (inp[10]) ? node24080 : 4'b1010;
															assign node24080 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node24083 = (inp[11]) ? 4'b1100 : node24084;
														assign node24084 = (inp[10]) ? 4'b1101 : node24085;
															assign node24085 = (inp[0]) ? node24089 : node24086;
																assign node24086 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node24089 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node24094 = (inp[15]) ? node24122 : node24095;
												assign node24095 = (inp[4]) ? node24113 : node24096;
													assign node24096 = (inp[0]) ? node24102 : node24097;
														assign node24097 = (inp[11]) ? node24099 : 4'b1010;
															assign node24099 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node24102 = (inp[9]) ? node24108 : node24103;
															assign node24103 = (inp[11]) ? node24105 : 4'b1011;
																assign node24105 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node24108 = (inp[10]) ? node24110 : 4'b1010;
																assign node24110 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node24113 = (inp[9]) ? 4'b1100 : node24114;
														assign node24114 = (inp[0]) ? node24118 : node24115;
															assign node24115 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node24118 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node24122 = (inp[11]) ? node24138 : node24123;
													assign node24123 = (inp[9]) ? node24129 : node24124;
														assign node24124 = (inp[10]) ? 4'b1010 : node24125;
															assign node24125 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node24129 = (inp[10]) ? node24135 : node24130;
															assign node24130 = (inp[0]) ? 4'b1010 : node24131;
																assign node24131 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node24135 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node24138 = (inp[0]) ? 4'b1011 : node24139;
														assign node24139 = (inp[9]) ? node24143 : node24140;
															assign node24140 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node24143 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node24147 = (inp[12]) ? node24195 : node24148;
											assign node24148 = (inp[4]) ? node24176 : node24149;
												assign node24149 = (inp[15]) ? node24165 : node24150;
													assign node24150 = (inp[11]) ? node24160 : node24151;
														assign node24151 = (inp[10]) ? 4'b1010 : node24152;
															assign node24152 = (inp[0]) ? node24156 : node24153;
																assign node24153 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node24156 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node24160 = (inp[10]) ? node24162 : 4'b1011;
															assign node24162 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node24165 = (inp[10]) ? node24173 : node24166;
														assign node24166 = (inp[11]) ? 4'b1110 : node24167;
															assign node24167 = (inp[0]) ? 4'b1111 : node24168;
																assign node24168 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node24173 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node24176 = (inp[15]) ? node24188 : node24177;
													assign node24177 = (inp[11]) ? 4'b1101 : node24178;
														assign node24178 = (inp[0]) ? 4'b1101 : node24179;
															assign node24179 = (inp[10]) ? node24183 : node24180;
																assign node24180 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node24183 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node24188 = (inp[11]) ? 4'b1010 : node24189;
														assign node24189 = (inp[0]) ? node24191 : 4'b1010;
															assign node24191 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node24195 = (inp[15]) ? node24213 : node24196;
												assign node24196 = (inp[4]) ? node24208 : node24197;
													assign node24197 = (inp[11]) ? node24201 : node24198;
														assign node24198 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node24201 = (inp[10]) ? 4'b1100 : node24202;
															assign node24202 = (inp[9]) ? 4'b1101 : node24203;
																assign node24203 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node24208 = (inp[9]) ? node24210 : 4'b1011;
														assign node24210 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node24213 = (inp[11]) ? node24231 : node24214;
													assign node24214 = (inp[0]) ? node24224 : node24215;
														assign node24215 = (inp[4]) ? node24217 : 4'b1000;
															assign node24217 = (inp[10]) ? node24221 : node24218;
																assign node24218 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node24221 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node24224 = (inp[4]) ? node24226 : 4'b1001;
															assign node24226 = (inp[9]) ? node24228 : 4'b1000;
																assign node24228 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node24231 = (inp[10]) ? node24233 : 4'b1001;
														assign node24233 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node24236 = (inp[7]) ? node24336 : node24237;
										assign node24237 = (inp[12]) ? node24281 : node24238;
											assign node24238 = (inp[15]) ? node24256 : node24239;
												assign node24239 = (inp[4]) ? node24247 : node24240;
													assign node24240 = (inp[0]) ? node24242 : 4'b1101;
														assign node24242 = (inp[11]) ? node24244 : 4'b1100;
															assign node24244 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node24247 = (inp[11]) ? node24249 : 4'b1111;
														assign node24249 = (inp[9]) ? node24253 : node24250;
															assign node24250 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node24253 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node24256 = (inp[4]) ? node24270 : node24257;
													assign node24257 = (inp[10]) ? node24259 : 4'b1101;
														assign node24259 = (inp[9]) ? node24265 : node24260;
															assign node24260 = (inp[11]) ? node24262 : 4'b1101;
																assign node24262 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node24265 = (inp[0]) ? 4'b1100 : node24266;
																assign node24266 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node24270 = (inp[9]) ? node24272 : 4'b1001;
														assign node24272 = (inp[0]) ? node24274 : 4'b1001;
															assign node24274 = (inp[11]) ? node24278 : node24275;
																assign node24275 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node24278 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node24281 = (inp[15]) ? node24303 : node24282;
												assign node24282 = (inp[4]) ? node24296 : node24283;
													assign node24283 = (inp[11]) ? node24289 : node24284;
														assign node24284 = (inp[10]) ? 4'b1110 : node24285;
															assign node24285 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node24289 = (inp[9]) ? node24293 : node24290;
															assign node24290 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node24293 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node24296 = (inp[11]) ? 4'b1100 : node24297;
														assign node24297 = (inp[10]) ? 4'b1101 : node24298;
															assign node24298 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node24303 = (inp[0]) ? node24317 : node24304;
													assign node24304 = (inp[9]) ? node24312 : node24305;
														assign node24305 = (inp[4]) ? 4'b1111 : node24306;
															assign node24306 = (inp[11]) ? 4'b1110 : node24307;
																assign node24307 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node24312 = (inp[10]) ? node24314 : 4'b1110;
															assign node24314 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node24317 = (inp[4]) ? node24323 : node24318;
														assign node24318 = (inp[10]) ? 4'b1111 : node24319;
															assign node24319 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node24323 = (inp[9]) ? node24331 : node24324;
															assign node24324 = (inp[11]) ? node24328 : node24325;
																assign node24325 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node24328 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node24331 = (inp[11]) ? 4'b1111 : node24332;
																assign node24332 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node24336 = (inp[12]) ? node24378 : node24337;
											assign node24337 = (inp[15]) ? node24355 : node24338;
												assign node24338 = (inp[4]) ? node24346 : node24339;
													assign node24339 = (inp[0]) ? 4'b1010 : node24340;
														assign node24340 = (inp[11]) ? node24342 : 4'b1011;
															assign node24342 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node24346 = (inp[9]) ? node24350 : node24347;
														assign node24347 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node24350 = (inp[10]) ? 4'b1000 : node24351;
															assign node24351 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node24355 = (inp[4]) ? node24365 : node24356;
													assign node24356 = (inp[10]) ? 4'b1111 : node24357;
														assign node24357 = (inp[9]) ? node24359 : 4'b1111;
															assign node24359 = (inp[11]) ? 4'b1110 : node24360;
																assign node24360 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node24365 = (inp[0]) ? node24373 : node24366;
														assign node24366 = (inp[10]) ? 4'b1010 : node24367;
															assign node24367 = (inp[11]) ? node24369 : 4'b1010;
																assign node24369 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node24373 = (inp[10]) ? node24375 : 4'b1011;
															assign node24375 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node24378 = (inp[4]) ? node24406 : node24379;
												assign node24379 = (inp[15]) ? node24401 : node24380;
													assign node24380 = (inp[0]) ? node24394 : node24381;
														assign node24381 = (inp[11]) ? node24389 : node24382;
															assign node24382 = (inp[10]) ? node24386 : node24383;
																assign node24383 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node24386 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node24389 = (inp[10]) ? 4'b1000 : node24390;
																assign node24390 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node24394 = (inp[10]) ? 4'b1001 : node24395;
															assign node24395 = (inp[11]) ? node24397 : 4'b1001;
																assign node24397 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node24401 = (inp[10]) ? node24403 : 4'b1100;
														assign node24403 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node24406 = (inp[15]) ? node24420 : node24407;
													assign node24407 = (inp[9]) ? node24411 : node24408;
														assign node24408 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node24411 = (inp[0]) ? node24415 : node24412;
															assign node24412 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node24415 = (inp[10]) ? node24417 : 4'b1110;
																assign node24417 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node24420 = (inp[0]) ? 4'b1101 : node24421;
														assign node24421 = (inp[11]) ? 4'b1101 : node24422;
															assign node24422 = (inp[10]) ? node24426 : node24423;
																assign node24423 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node24426 = (inp[9]) ? 4'b1100 : 4'b1101;
								assign node24431 = (inp[12]) ? node24565 : node24432;
									assign node24432 = (inp[15]) ? node24486 : node24433;
										assign node24433 = (inp[7]) ? node24463 : node24434;
											assign node24434 = (inp[1]) ? node24450 : node24435;
												assign node24435 = (inp[0]) ? node24437 : 4'b1101;
													assign node24437 = (inp[11]) ? node24445 : node24438;
														assign node24438 = (inp[10]) ? node24440 : 4'b1101;
															assign node24440 = (inp[9]) ? node24442 : 4'b1100;
																assign node24442 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node24445 = (inp[4]) ? 4'b1101 : node24446;
															assign node24446 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node24450 = (inp[4]) ? node24458 : node24451;
													assign node24451 = (inp[0]) ? 4'b1001 : node24452;
														assign node24452 = (inp[11]) ? 4'b1000 : node24453;
															assign node24453 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node24458 = (inp[9]) ? node24460 : 4'b1101;
														assign node24460 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node24463 = (inp[1]) ? node24475 : node24464;
												assign node24464 = (inp[4]) ? node24470 : node24465;
													assign node24465 = (inp[11]) ? node24467 : 4'b1111;
														assign node24467 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node24470 = (inp[9]) ? node24472 : 4'b1010;
														assign node24472 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node24475 = (inp[11]) ? node24481 : node24476;
													assign node24476 = (inp[4]) ? node24478 : 4'b1110;
														assign node24478 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node24481 = (inp[9]) ? node24483 : 4'b1111;
														assign node24483 = (inp[4]) ? 4'b1110 : 4'b1111;
										assign node24486 = (inp[7]) ? node24530 : node24487;
											assign node24487 = (inp[4]) ? node24515 : node24488;
												assign node24488 = (inp[1]) ? node24506 : node24489;
													assign node24489 = (inp[11]) ? node24501 : node24490;
														assign node24490 = (inp[10]) ? node24496 : node24491;
															assign node24491 = (inp[0]) ? node24493 : 4'b1111;
																assign node24493 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node24496 = (inp[9]) ? node24498 : 4'b1110;
																assign node24498 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node24501 = (inp[9]) ? 4'b1111 : node24502;
															assign node24502 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node24506 = (inp[0]) ? node24508 : 4'b1011;
														assign node24508 = (inp[10]) ? node24510 : 4'b1010;
															assign node24510 = (inp[11]) ? node24512 : 4'b1011;
																assign node24512 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node24515 = (inp[1]) ? node24521 : node24516;
													assign node24516 = (inp[11]) ? node24518 : 4'b1011;
														assign node24518 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node24521 = (inp[10]) ? node24523 : 4'b1111;
														assign node24523 = (inp[11]) ? node24525 : 4'b1111;
															assign node24525 = (inp[0]) ? node24527 : 4'b1111;
																assign node24527 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node24530 = (inp[4]) ? node24548 : node24531;
												assign node24531 = (inp[1]) ? node24541 : node24532;
													assign node24532 = (inp[10]) ? 4'b1101 : node24533;
														assign node24533 = (inp[0]) ? 4'b1100 : node24534;
															assign node24534 = (inp[9]) ? node24536 : 4'b1101;
																assign node24536 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node24541 = (inp[11]) ? node24545 : node24542;
														assign node24542 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node24545 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node24548 = (inp[1]) ? node24558 : node24549;
													assign node24549 = (inp[0]) ? 4'b1000 : node24550;
														assign node24550 = (inp[10]) ? node24552 : 4'b1000;
															assign node24552 = (inp[11]) ? 4'b1001 : node24553;
																assign node24553 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node24558 = (inp[11]) ? node24562 : node24559;
														assign node24559 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node24562 = (inp[9]) ? 4'b1100 : 4'b1101;
									assign node24565 = (inp[15]) ? node24641 : node24566;
										assign node24566 = (inp[7]) ? node24600 : node24567;
											assign node24567 = (inp[4]) ? node24581 : node24568;
												assign node24568 = (inp[9]) ? node24574 : node24569;
													assign node24569 = (inp[11]) ? 4'b1101 : node24570;
														assign node24570 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node24574 = (inp[11]) ? node24576 : 4'b1101;
														assign node24576 = (inp[0]) ? 4'b1100 : node24577;
															assign node24577 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node24581 = (inp[1]) ? node24589 : node24582;
													assign node24582 = (inp[9]) ? node24586 : node24583;
														assign node24583 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node24586 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node24589 = (inp[11]) ? node24595 : node24590;
														assign node24590 = (inp[9]) ? 4'b1000 : node24591;
															assign node24591 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node24595 = (inp[9]) ? 4'b1001 : node24596;
															assign node24596 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node24600 = (inp[4]) ? node24618 : node24601;
												assign node24601 = (inp[1]) ? node24609 : node24602;
													assign node24602 = (inp[9]) ? 4'b1010 : node24603;
														assign node24603 = (inp[0]) ? node24605 : 4'b1011;
															assign node24605 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node24609 = (inp[10]) ? 4'b1110 : node24610;
														assign node24610 = (inp[11]) ? 4'b1111 : node24611;
															assign node24611 = (inp[9]) ? node24613 : 4'b1111;
																assign node24613 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node24618 = (inp[0]) ? node24628 : node24619;
													assign node24619 = (inp[11]) ? node24621 : 4'b1110;
														assign node24621 = (inp[1]) ? node24625 : node24622;
															assign node24622 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node24625 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node24628 = (inp[1]) ? node24636 : node24629;
														assign node24629 = (inp[11]) ? node24633 : node24630;
															assign node24630 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node24633 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node24636 = (inp[9]) ? 4'b1111 : node24637;
															assign node24637 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node24641 = (inp[7]) ? node24695 : node24642;
											assign node24642 = (inp[1]) ? node24668 : node24643;
												assign node24643 = (inp[4]) ? node24653 : node24644;
													assign node24644 = (inp[10]) ? 4'b1111 : node24645;
														assign node24645 = (inp[11]) ? node24647 : 4'b1111;
															assign node24647 = (inp[0]) ? 4'b1110 : node24648;
																assign node24648 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node24653 = (inp[0]) ? node24661 : node24654;
														assign node24654 = (inp[11]) ? node24658 : node24655;
															assign node24655 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node24658 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node24661 = (inp[9]) ? node24665 : node24662;
															assign node24662 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node24665 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node24668 = (inp[10]) ? node24674 : node24669;
													assign node24669 = (inp[0]) ? 4'b1110 : node24670;
														assign node24670 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node24674 = (inp[4]) ? node24684 : node24675;
														assign node24675 = (inp[11]) ? 4'b1110 : node24676;
															assign node24676 = (inp[0]) ? node24680 : node24677;
																assign node24677 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node24680 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node24684 = (inp[0]) ? node24690 : node24685;
															assign node24685 = (inp[9]) ? node24687 : 4'b1110;
																assign node24687 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node24690 = (inp[9]) ? 4'b1111 : node24691;
																assign node24691 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node24695 = (inp[0]) ? node24713 : node24696;
												assign node24696 = (inp[10]) ? node24708 : node24697;
													assign node24697 = (inp[4]) ? node24703 : node24698;
														assign node24698 = (inp[1]) ? 4'b1100 : node24699;
															assign node24699 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node24703 = (inp[11]) ? 4'b1101 : node24704;
															assign node24704 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node24708 = (inp[9]) ? node24710 : 4'b1100;
														assign node24710 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node24713 = (inp[11]) ? node24717 : node24714;
													assign node24714 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node24717 = (inp[9]) ? 4'b1100 : 4'b1101;
							assign node24720 = (inp[12]) ? node25068 : node24721;
								assign node24721 = (inp[7]) ? node24899 : node24722;
									assign node24722 = (inp[15]) ? node24798 : node24723;
										assign node24723 = (inp[4]) ? node24757 : node24724;
											assign node24724 = (inp[1]) ? node24744 : node24725;
												assign node24725 = (inp[0]) ? node24735 : node24726;
													assign node24726 = (inp[9]) ? node24732 : node24727;
														assign node24727 = (inp[10]) ? node24729 : 4'b1001;
															assign node24729 = (inp[6]) ? 4'b1001 : 4'b1000;
														assign node24732 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node24735 = (inp[9]) ? node24739 : node24736;
														assign node24736 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node24739 = (inp[11]) ? 4'b1001 : node24740;
															assign node24740 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node24744 = (inp[6]) ? node24750 : node24745;
													assign node24745 = (inp[11]) ? node24747 : 4'b1000;
														assign node24747 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node24750 = (inp[11]) ? node24754 : node24751;
														assign node24751 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node24754 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node24757 = (inp[6]) ? node24781 : node24758;
												assign node24758 = (inp[11]) ? node24770 : node24759;
													assign node24759 = (inp[9]) ? node24767 : node24760;
														assign node24760 = (inp[10]) ? node24764 : node24761;
															assign node24761 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node24764 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node24767 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node24770 = (inp[10]) ? 4'b1011 : node24771;
														assign node24771 = (inp[1]) ? 4'b1010 : node24772;
															assign node24772 = (inp[9]) ? node24776 : node24773;
																assign node24773 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node24776 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node24781 = (inp[9]) ? node24789 : node24782;
													assign node24782 = (inp[0]) ? node24784 : 4'b1001;
														assign node24784 = (inp[10]) ? 4'b1000 : node24785;
															assign node24785 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node24789 = (inp[11]) ? node24795 : node24790;
														assign node24790 = (inp[1]) ? 4'b1000 : node24791;
															assign node24791 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node24795 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node24798 = (inp[6]) ? node24856 : node24799;
											assign node24799 = (inp[4]) ? node24835 : node24800;
												assign node24800 = (inp[0]) ? node24814 : node24801;
													assign node24801 = (inp[10]) ? node24807 : node24802;
														assign node24802 = (inp[11]) ? node24804 : 4'b1000;
															assign node24804 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node24807 = (inp[1]) ? node24811 : node24808;
															assign node24808 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node24811 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node24814 = (inp[9]) ? node24830 : node24815;
														assign node24815 = (inp[10]) ? node24823 : node24816;
															assign node24816 = (inp[11]) ? node24820 : node24817;
																assign node24817 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node24820 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node24823 = (inp[1]) ? node24827 : node24824;
																assign node24824 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node24827 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node24830 = (inp[11]) ? 4'b1001 : node24831;
															assign node24831 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node24835 = (inp[9]) ? node24843 : node24836;
													assign node24836 = (inp[11]) ? 4'b1101 : node24837;
														assign node24837 = (inp[1]) ? 4'b1100 : node24838;
															assign node24838 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node24843 = (inp[1]) ? node24849 : node24844;
														assign node24844 = (inp[10]) ? node24846 : 4'b1100;
															assign node24846 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node24849 = (inp[10]) ? node24851 : 4'b1101;
															assign node24851 = (inp[0]) ? 4'b1100 : node24852;
																assign node24852 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node24856 = (inp[11]) ? node24880 : node24857;
												assign node24857 = (inp[9]) ? node24869 : node24858;
													assign node24858 = (inp[4]) ? node24864 : node24859;
														assign node24859 = (inp[1]) ? node24861 : 4'b1010;
															assign node24861 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node24864 = (inp[1]) ? 4'b1010 : node24865;
															assign node24865 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node24869 = (inp[0]) ? node24875 : node24870;
														assign node24870 = (inp[1]) ? 4'b1110 : node24871;
															assign node24871 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node24875 = (inp[4]) ? 4'b1011 : node24876;
															assign node24876 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node24880 = (inp[0]) ? node24888 : node24881;
													assign node24881 = (inp[4]) ? node24885 : node24882;
														assign node24882 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node24885 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node24888 = (inp[1]) ? node24894 : node24889;
														assign node24889 = (inp[4]) ? node24891 : 4'b1010;
															assign node24891 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node24894 = (inp[9]) ? 4'b1110 : node24895;
															assign node24895 = (inp[4]) ? 4'b1011 : 4'b1111;
									assign node24899 = (inp[6]) ? node24987 : node24900;
										assign node24900 = (inp[15]) ? node24942 : node24901;
											assign node24901 = (inp[4]) ? node24917 : node24902;
												assign node24902 = (inp[1]) ? node24914 : node24903;
													assign node24903 = (inp[10]) ? node24909 : node24904;
														assign node24904 = (inp[9]) ? 4'b1111 : node24905;
															assign node24905 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node24909 = (inp[9]) ? 4'b1110 : node24910;
															assign node24910 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node24914 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node24917 = (inp[10]) ? node24931 : node24918;
													assign node24918 = (inp[0]) ? node24924 : node24919;
														assign node24919 = (inp[9]) ? 4'b1101 : node24920;
															assign node24920 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node24924 = (inp[9]) ? node24928 : node24925;
															assign node24925 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node24928 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node24931 = (inp[0]) ? node24937 : node24932;
														assign node24932 = (inp[9]) ? 4'b1100 : node24933;
															assign node24933 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node24937 = (inp[9]) ? 4'b1101 : node24938;
															assign node24938 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node24942 = (inp[1]) ? node24970 : node24943;
												assign node24943 = (inp[4]) ? node24957 : node24944;
													assign node24944 = (inp[0]) ? node24952 : node24945;
														assign node24945 = (inp[11]) ? node24947 : 4'b1010;
															assign node24947 = (inp[9]) ? node24949 : 4'b1010;
																assign node24949 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node24952 = (inp[11]) ? 4'b1011 : node24953;
															assign node24953 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node24957 = (inp[10]) ? node24961 : node24958;
														assign node24958 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node24961 = (inp[9]) ? node24967 : node24962;
															assign node24962 = (inp[11]) ? 4'b1110 : node24963;
																assign node24963 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node24967 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node24970 = (inp[4]) ? node24972 : 4'b1111;
													assign node24972 = (inp[9]) ? node24980 : node24973;
														assign node24973 = (inp[10]) ? 4'b1011 : node24974;
															assign node24974 = (inp[11]) ? 4'b1010 : node24975;
																assign node24975 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node24980 = (inp[10]) ? node24982 : 4'b1011;
															assign node24982 = (inp[0]) ? node24984 : 4'b1010;
																assign node24984 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node24987 = (inp[15]) ? node25027 : node24988;
											assign node24988 = (inp[1]) ? node25012 : node24989;
												assign node24989 = (inp[4]) ? node24999 : node24990;
													assign node24990 = (inp[0]) ? node24992 : 4'b1010;
														assign node24992 = (inp[9]) ? node24996 : node24993;
															assign node24993 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node24996 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node24999 = (inp[11]) ? node25005 : node25000;
														assign node25000 = (inp[9]) ? node25002 : 4'b1110;
															assign node25002 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node25005 = (inp[9]) ? node25009 : node25006;
															assign node25006 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node25009 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node25012 = (inp[4]) ? node25020 : node25013;
													assign node25013 = (inp[0]) ? node25015 : 4'b1011;
														assign node25015 = (inp[9]) ? 4'b1011 : node25016;
															assign node25016 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node25020 = (inp[11]) ? node25024 : node25021;
														assign node25021 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node25024 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node25027 = (inp[4]) ? node25045 : node25028;
												assign node25028 = (inp[1]) ? node25036 : node25029;
													assign node25029 = (inp[11]) ? 4'b1000 : node25030;
														assign node25030 = (inp[0]) ? 4'b1000 : node25031;
															assign node25031 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node25036 = (inp[10]) ? 4'b1100 : node25037;
														assign node25037 = (inp[11]) ? node25041 : node25038;
															assign node25038 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node25041 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node25045 = (inp[1]) ? node25053 : node25046;
													assign node25046 = (inp[0]) ? node25050 : node25047;
														assign node25047 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node25050 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node25053 = (inp[0]) ? node25061 : node25054;
														assign node25054 = (inp[10]) ? node25056 : 4'b1001;
															assign node25056 = (inp[9]) ? 4'b1001 : node25057;
																assign node25057 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node25061 = (inp[10]) ? node25065 : node25062;
															assign node25062 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node25065 = (inp[9]) ? 4'b1000 : 4'b1001;
								assign node25068 = (inp[15]) ? node25232 : node25069;
									assign node25069 = (inp[7]) ? node25141 : node25070;
										assign node25070 = (inp[4]) ? node25104 : node25071;
											assign node25071 = (inp[6]) ? node25091 : node25072;
												assign node25072 = (inp[0]) ? node25076 : node25073;
													assign node25073 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node25076 = (inp[9]) ? node25088 : node25077;
														assign node25077 = (inp[10]) ? node25083 : node25078;
															assign node25078 = (inp[11]) ? node25080 : 4'b1010;
																assign node25080 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node25083 = (inp[11]) ? node25085 : 4'b1011;
																assign node25085 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node25088 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node25091 = (inp[0]) ? node25099 : node25092;
													assign node25092 = (inp[9]) ? node25096 : node25093;
														assign node25093 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node25096 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node25099 = (inp[11]) ? 4'b1000 : node25100;
														assign node25100 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node25104 = (inp[1]) ? node25120 : node25105;
												assign node25105 = (inp[10]) ? node25113 : node25106;
													assign node25106 = (inp[9]) ? node25108 : 4'b1001;
														assign node25108 = (inp[6]) ? node25110 : 4'b1000;
															assign node25110 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node25113 = (inp[0]) ? node25115 : 4'b1000;
														assign node25115 = (inp[9]) ? node25117 : 4'b1001;
															assign node25117 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node25120 = (inp[0]) ? node25130 : node25121;
													assign node25121 = (inp[9]) ? node25123 : 4'b1100;
														assign node25123 = (inp[11]) ? node25127 : node25124;
															assign node25124 = (inp[6]) ? 4'b1101 : 4'b1100;
															assign node25127 = (inp[6]) ? 4'b1100 : 4'b1101;
													assign node25130 = (inp[9]) ? 4'b1101 : node25131;
														assign node25131 = (inp[10]) ? 4'b1101 : node25132;
															assign node25132 = (inp[11]) ? node25136 : node25133;
																assign node25133 = (inp[6]) ? 4'b1100 : 4'b1101;
																assign node25136 = (inp[6]) ? 4'b1101 : 4'b1100;
										assign node25141 = (inp[4]) ? node25189 : node25142;
											assign node25142 = (inp[6]) ? node25168 : node25143;
												assign node25143 = (inp[9]) ? node25153 : node25144;
													assign node25144 = (inp[0]) ? 4'b1100 : node25145;
														assign node25145 = (inp[10]) ? 4'b1101 : node25146;
															assign node25146 = (inp[11]) ? node25148 : 4'b1100;
																assign node25148 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node25153 = (inp[10]) ? node25159 : node25154;
														assign node25154 = (inp[11]) ? 4'b1101 : node25155;
															assign node25155 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node25159 = (inp[0]) ? node25163 : node25160;
															assign node25160 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node25163 = (inp[1]) ? node25165 : 4'b1100;
																assign node25165 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node25168 = (inp[1]) ? node25182 : node25169;
													assign node25169 = (inp[11]) ? node25177 : node25170;
														assign node25170 = (inp[0]) ? node25174 : node25171;
															assign node25171 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node25174 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node25177 = (inp[9]) ? 4'b1111 : node25178;
															assign node25178 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node25182 = (inp[9]) ? node25186 : node25183;
														assign node25183 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node25186 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node25189 = (inp[6]) ? node25219 : node25190;
												assign node25190 = (inp[0]) ? node25204 : node25191;
													assign node25191 = (inp[10]) ? node25195 : node25192;
														assign node25192 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node25195 = (inp[9]) ? node25199 : node25196;
															assign node25196 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node25199 = (inp[1]) ? 4'b1010 : node25200;
																assign node25200 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node25204 = (inp[9]) ? node25212 : node25205;
														assign node25205 = (inp[11]) ? node25209 : node25206;
															assign node25206 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node25209 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node25212 = (inp[11]) ? node25216 : node25213;
															assign node25213 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node25216 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node25219 = (inp[10]) ? node25227 : node25220;
													assign node25220 = (inp[11]) ? 4'b1010 : node25221;
														assign node25221 = (inp[0]) ? 4'b1011 : node25222;
															assign node25222 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node25227 = (inp[9]) ? 4'b1011 : node25228;
														assign node25228 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node25232 = (inp[7]) ? node25290 : node25233;
										assign node25233 = (inp[4]) ? node25263 : node25234;
											assign node25234 = (inp[9]) ? node25252 : node25235;
												assign node25235 = (inp[11]) ? node25247 : node25236;
													assign node25236 = (inp[6]) ? 4'b1010 : node25237;
														assign node25237 = (inp[1]) ? node25243 : node25238;
															assign node25238 = (inp[10]) ? 4'b1011 : node25239;
																assign node25239 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node25243 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node25247 = (inp[6]) ? 4'b1011 : node25248;
														assign node25248 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node25252 = (inp[11]) ? node25260 : node25253;
													assign node25253 = (inp[10]) ? 4'b1011 : node25254;
														assign node25254 = (inp[0]) ? node25256 : 4'b1011;
															assign node25256 = (inp[6]) ? 4'b1011 : 4'b1010;
													assign node25260 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node25263 = (inp[9]) ? node25277 : node25264;
												assign node25264 = (inp[11]) ? node25272 : node25265;
													assign node25265 = (inp[6]) ? 4'b1010 : node25266;
														assign node25266 = (inp[10]) ? node25268 : 4'b1011;
															assign node25268 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node25272 = (inp[6]) ? 4'b1011 : node25273;
														assign node25273 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node25277 = (inp[11]) ? node25285 : node25278;
													assign node25278 = (inp[6]) ? 4'b1011 : node25279;
														assign node25279 = (inp[10]) ? node25281 : 4'b1010;
															assign node25281 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node25285 = (inp[10]) ? 4'b1010 : node25286;
														assign node25286 = (inp[1]) ? 4'b1010 : 4'b1011;
										assign node25290 = (inp[9]) ? node25308 : node25291;
											assign node25291 = (inp[11]) ? node25303 : node25292;
												assign node25292 = (inp[6]) ? 4'b1000 : node25293;
													assign node25293 = (inp[4]) ? node25295 : 4'b1001;
														assign node25295 = (inp[1]) ? node25297 : 4'b1001;
															assign node25297 = (inp[0]) ? node25299 : 4'b1001;
																assign node25299 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node25303 = (inp[6]) ? 4'b1001 : node25304;
													assign node25304 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node25308 = (inp[11]) ? node25320 : node25309;
												assign node25309 = (inp[6]) ? 4'b1001 : node25310;
													assign node25310 = (inp[4]) ? 4'b1001 : node25311;
														assign node25311 = (inp[1]) ? 4'b1001 : node25312;
															assign node25312 = (inp[10]) ? node25314 : 4'b1000;
																assign node25314 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node25320 = (inp[10]) ? 4'b1000 : node25321;
													assign node25321 = (inp[6]) ? 4'b1000 : 4'b1001;
				assign node25325 = (inp[7]) ? node27719 : node25326;
					assign node25326 = (inp[6]) ? node26938 : node25327;
						assign node25327 = (inp[12]) ? node26111 : node25328;
							assign node25328 = (inp[15]) ? node25702 : node25329;
								assign node25329 = (inp[4]) ? node25529 : node25330;
									assign node25330 = (inp[0]) ? node25424 : node25331;
										assign node25331 = (inp[10]) ? node25373 : node25332;
											assign node25332 = (inp[9]) ? node25348 : node25333;
												assign node25333 = (inp[2]) ? node25343 : node25334;
													assign node25334 = (inp[5]) ? node25340 : node25335;
														assign node25335 = (inp[13]) ? 4'b0110 : node25336;
															assign node25336 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25340 = (inp[13]) ? 4'b0011 : 4'b0110;
													assign node25343 = (inp[11]) ? node25345 : 4'b0011;
														assign node25345 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node25348 = (inp[13]) ? node25364 : node25349;
													assign node25349 = (inp[2]) ? node25359 : node25350;
														assign node25350 = (inp[11]) ? node25354 : node25351;
															assign node25351 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node25354 = (inp[5]) ? node25356 : 4'b0110;
																assign node25356 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node25359 = (inp[1]) ? node25361 : 4'b0111;
															assign node25361 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node25364 = (inp[1]) ? node25370 : node25365;
														assign node25365 = (inp[11]) ? node25367 : 4'b0010;
															assign node25367 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25370 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node25373 = (inp[13]) ? node25411 : node25374;
												assign node25374 = (inp[2]) ? node25394 : node25375;
													assign node25375 = (inp[1]) ? node25385 : node25376;
														assign node25376 = (inp[5]) ? node25382 : node25377;
															assign node25377 = (inp[11]) ? 4'b0011 : node25378;
																assign node25378 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node25382 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25385 = (inp[9]) ? node25389 : node25386;
															assign node25386 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25389 = (inp[11]) ? node25391 : 4'b0110;
																assign node25391 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node25394 = (inp[1]) ? node25406 : node25395;
														assign node25395 = (inp[5]) ? node25399 : node25396;
															assign node25396 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25399 = (inp[9]) ? node25403 : node25400;
																assign node25400 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node25403 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node25406 = (inp[9]) ? 4'b0011 : node25407;
															assign node25407 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node25411 = (inp[2]) ? node25419 : node25412;
													assign node25412 = (inp[1]) ? 4'b0010 : node25413;
														assign node25413 = (inp[5]) ? node25415 : 4'b0110;
															assign node25415 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node25419 = (inp[9]) ? 4'b0111 : node25420;
														assign node25420 = (inp[11]) ? 4'b0110 : 4'b0010;
										assign node25424 = (inp[13]) ? node25478 : node25425;
											assign node25425 = (inp[2]) ? node25455 : node25426;
												assign node25426 = (inp[5]) ? node25436 : node25427;
													assign node25427 = (inp[1]) ? 4'b0110 : node25428;
														assign node25428 = (inp[11]) ? node25432 : node25429;
															assign node25429 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node25432 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node25436 = (inp[11]) ? node25446 : node25437;
														assign node25437 = (inp[10]) ? node25439 : 4'b0111;
															assign node25439 = (inp[9]) ? node25443 : node25440;
																assign node25440 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node25443 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25446 = (inp[1]) ? node25452 : node25447;
															assign node25447 = (inp[10]) ? node25449 : 4'b0110;
																assign node25449 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25452 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node25455 = (inp[5]) ? node25465 : node25456;
													assign node25456 = (inp[1]) ? node25458 : 4'b0110;
														assign node25458 = (inp[10]) ? node25462 : node25459;
															assign node25459 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node25462 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node25465 = (inp[9]) ? node25471 : node25466;
														assign node25466 = (inp[10]) ? node25468 : 4'b0010;
															assign node25468 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node25471 = (inp[10]) ? node25473 : 4'b0011;
															assign node25473 = (inp[1]) ? node25475 : 4'b0010;
																assign node25475 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node25478 = (inp[2]) ? node25498 : node25479;
												assign node25479 = (inp[5]) ? node25491 : node25480;
													assign node25480 = (inp[1]) ? 4'b0011 : node25481;
														assign node25481 = (inp[10]) ? 4'b0111 : node25482;
															assign node25482 = (inp[11]) ? node25486 : node25483;
																assign node25483 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node25486 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25491 = (inp[1]) ? node25493 : 4'b0011;
														assign node25493 = (inp[10]) ? node25495 : 4'b0010;
															assign node25495 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node25498 = (inp[1]) ? node25512 : node25499;
													assign node25499 = (inp[5]) ? node25503 : node25500;
														assign node25500 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25503 = (inp[11]) ? 4'b0111 : node25504;
															assign node25504 = (inp[10]) ? node25508 : node25505;
																assign node25505 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node25508 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node25512 = (inp[5]) ? node25526 : node25513;
														assign node25513 = (inp[11]) ? node25519 : node25514;
															assign node25514 = (inp[10]) ? 4'b0111 : node25515;
																assign node25515 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node25519 = (inp[10]) ? node25523 : node25520;
																assign node25520 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node25523 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node25526 = (inp[9]) ? 4'b0111 : 4'b0110;
									assign node25529 = (inp[2]) ? node25631 : node25530;
										assign node25530 = (inp[13]) ? node25584 : node25531;
											assign node25531 = (inp[1]) ? node25559 : node25532;
												assign node25532 = (inp[11]) ? node25546 : node25533;
													assign node25533 = (inp[10]) ? node25539 : node25534;
														assign node25534 = (inp[0]) ? node25536 : 4'b0001;
															assign node25536 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node25539 = (inp[9]) ? node25543 : node25540;
															assign node25540 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node25543 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node25546 = (inp[0]) ? node25552 : node25547;
														assign node25547 = (inp[9]) ? node25549 : 4'b0000;
															assign node25549 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node25552 = (inp[5]) ? node25556 : node25553;
															assign node25553 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node25556 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node25559 = (inp[5]) ? node25571 : node25560;
													assign node25560 = (inp[9]) ? node25562 : 4'b0000;
														assign node25562 = (inp[10]) ? node25566 : node25563;
															assign node25563 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node25566 = (inp[11]) ? node25568 : 4'b0000;
																assign node25568 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node25571 = (inp[9]) ? node25581 : node25572;
														assign node25572 = (inp[10]) ? node25576 : node25573;
															assign node25573 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node25576 = (inp[0]) ? 4'b0101 : node25577;
																assign node25577 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node25581 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node25584 = (inp[1]) ? node25604 : node25585;
												assign node25585 = (inp[0]) ? node25597 : node25586;
													assign node25586 = (inp[9]) ? node25592 : node25587;
														assign node25587 = (inp[10]) ? node25589 : 4'b0101;
															assign node25589 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node25592 = (inp[11]) ? 4'b0100 : node25593;
															assign node25593 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node25597 = (inp[9]) ? node25599 : 4'b0101;
														assign node25599 = (inp[10]) ? 4'b0101 : node25600;
															assign node25600 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node25604 = (inp[5]) ? node25616 : node25605;
													assign node25605 = (inp[10]) ? node25611 : node25606;
														assign node25606 = (inp[9]) ? 4'b0101 : node25607;
															assign node25607 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node25611 = (inp[9]) ? 4'b0100 : node25612;
															assign node25612 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node25616 = (inp[10]) ? node25626 : node25617;
														assign node25617 = (inp[9]) ? node25621 : node25618;
															assign node25618 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node25621 = (inp[11]) ? 4'b0000 : node25622;
																assign node25622 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node25626 = (inp[9]) ? 4'b0001 : node25627;
															assign node25627 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node25631 = (inp[13]) ? node25669 : node25632;
											assign node25632 = (inp[1]) ? node25650 : node25633;
												assign node25633 = (inp[11]) ? node25645 : node25634;
													assign node25634 = (inp[0]) ? 4'b0100 : node25635;
														assign node25635 = (inp[9]) ? node25637 : 4'b0101;
															assign node25637 = (inp[10]) ? node25641 : node25638;
																assign node25638 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node25641 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node25645 = (inp[9]) ? node25647 : 4'b0101;
														assign node25647 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node25650 = (inp[5]) ? node25656 : node25651;
													assign node25651 = (inp[10]) ? 4'b0101 : node25652;
														assign node25652 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node25656 = (inp[11]) ? node25658 : 4'b0001;
														assign node25658 = (inp[0]) ? node25664 : node25659;
															assign node25659 = (inp[9]) ? node25661 : 4'b0000;
																assign node25661 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node25664 = (inp[10]) ? node25666 : 4'b0001;
																assign node25666 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node25669 = (inp[5]) ? node25685 : node25670;
												assign node25670 = (inp[10]) ? node25678 : node25671;
													assign node25671 = (inp[9]) ? 4'b0001 : node25672;
														assign node25672 = (inp[0]) ? node25674 : 4'b0001;
															assign node25674 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node25678 = (inp[9]) ? node25680 : 4'b0001;
														assign node25680 = (inp[0]) ? 4'b0000 : node25681;
															assign node25681 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node25685 = (inp[1]) ? node25697 : node25686;
													assign node25686 = (inp[9]) ? node25688 : 4'b0000;
														assign node25688 = (inp[11]) ? node25692 : node25689;
															assign node25689 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node25692 = (inp[10]) ? node25694 : 4'b0001;
																assign node25694 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node25697 = (inp[9]) ? node25699 : 4'b0101;
														assign node25699 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node25702 = (inp[2]) ? node25912 : node25703;
									assign node25703 = (inp[9]) ? node25803 : node25704;
										assign node25704 = (inp[1]) ? node25744 : node25705;
											assign node25705 = (inp[10]) ? node25729 : node25706;
												assign node25706 = (inp[5]) ? node25718 : node25707;
													assign node25707 = (inp[4]) ? node25715 : node25708;
														assign node25708 = (inp[13]) ? node25712 : node25709;
															assign node25709 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node25712 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node25715 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node25718 = (inp[13]) ? node25724 : node25719;
														assign node25719 = (inp[4]) ? node25721 : 4'b0001;
															assign node25721 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node25724 = (inp[4]) ? 4'b0001 : node25725;
															assign node25725 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node25729 = (inp[4]) ? node25741 : node25730;
													assign node25730 = (inp[13]) ? node25736 : node25731;
														assign node25731 = (inp[5]) ? 4'b0001 : node25732;
															assign node25732 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node25736 = (inp[11]) ? 4'b0101 : node25737;
															assign node25737 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node25741 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node25744 = (inp[10]) ? node25768 : node25745;
												assign node25745 = (inp[5]) ? node25761 : node25746;
													assign node25746 = (inp[11]) ? node25756 : node25747;
														assign node25747 = (inp[0]) ? node25753 : node25748;
															assign node25748 = (inp[13]) ? node25750 : 4'b0001;
																assign node25750 = (inp[4]) ? 4'b0001 : 4'b0100;
															assign node25753 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25756 = (inp[4]) ? node25758 : 4'b0101;
															assign node25758 = (inp[0]) ? 4'b0000 : 4'b0100;
													assign node25761 = (inp[4]) ? 4'b0001 : node25762;
														assign node25762 = (inp[13]) ? node25764 : 4'b0100;
															assign node25764 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node25768 = (inp[5]) ? node25788 : node25769;
													assign node25769 = (inp[0]) ? node25775 : node25770;
														assign node25770 = (inp[4]) ? 4'b0100 : node25771;
															assign node25771 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node25775 = (inp[11]) ? node25783 : node25776;
															assign node25776 = (inp[13]) ? node25780 : node25777;
																assign node25777 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node25780 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node25783 = (inp[13]) ? node25785 : 4'b0001;
																assign node25785 = (inp[4]) ? 4'b0001 : 4'b0100;
													assign node25788 = (inp[4]) ? node25796 : node25789;
														assign node25789 = (inp[13]) ? node25791 : 4'b0101;
															assign node25791 = (inp[11]) ? 4'b0001 : node25792;
																assign node25792 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node25796 = (inp[13]) ? node25800 : node25797;
															assign node25797 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node25800 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node25803 = (inp[5]) ? node25869 : node25804;
											assign node25804 = (inp[4]) ? node25838 : node25805;
												assign node25805 = (inp[13]) ? node25823 : node25806;
													assign node25806 = (inp[0]) ? node25814 : node25807;
														assign node25807 = (inp[11]) ? node25809 : 4'b0000;
															assign node25809 = (inp[10]) ? node25811 : 4'b0000;
																assign node25811 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node25814 = (inp[11]) ? node25818 : node25815;
															assign node25815 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node25818 = (inp[1]) ? 4'b0000 : node25819;
																assign node25819 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node25823 = (inp[11]) ? node25825 : 4'b0100;
														assign node25825 = (inp[0]) ? node25833 : node25826;
															assign node25826 = (inp[10]) ? node25830 : node25827;
																assign node25827 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node25830 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node25833 = (inp[10]) ? node25835 : 4'b0100;
																assign node25835 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node25838 = (inp[13]) ? node25852 : node25839;
													assign node25839 = (inp[10]) ? node25847 : node25840;
														assign node25840 = (inp[1]) ? node25842 : 4'b0100;
															assign node25842 = (inp[11]) ? 4'b0101 : node25843;
																assign node25843 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node25847 = (inp[1]) ? node25849 : 4'b0101;
															assign node25849 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node25852 = (inp[11]) ? node25860 : node25853;
														assign node25853 = (inp[0]) ? 4'b0001 : node25854;
															assign node25854 = (inp[1]) ? 4'b0001 : node25855;
																assign node25855 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node25860 = (inp[0]) ? node25864 : node25861;
															assign node25861 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node25864 = (inp[1]) ? node25866 : 4'b0001;
																assign node25866 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node25869 = (inp[4]) ? node25887 : node25870;
												assign node25870 = (inp[10]) ? node25880 : node25871;
													assign node25871 = (inp[13]) ? node25875 : node25872;
														assign node25872 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node25875 = (inp[1]) ? 4'b0001 : node25876;
															assign node25876 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node25880 = (inp[1]) ? node25882 : 4'b0101;
														assign node25882 = (inp[13]) ? 4'b0000 : node25883;
															assign node25883 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node25887 = (inp[0]) ? node25893 : node25888;
													assign node25888 = (inp[10]) ? node25890 : 4'b0100;
														assign node25890 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node25893 = (inp[13]) ? node25901 : node25894;
														assign node25894 = (inp[1]) ? node25898 : node25895;
															assign node25895 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node25898 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node25901 = (inp[1]) ? node25905 : node25902;
															assign node25902 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node25905 = (inp[10]) ? node25909 : node25906;
																assign node25906 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node25909 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node25912 = (inp[5]) ? node26012 : node25913;
										assign node25913 = (inp[10]) ? node25955 : node25914;
											assign node25914 = (inp[13]) ? node25936 : node25915;
												assign node25915 = (inp[4]) ? node25925 : node25916;
													assign node25916 = (inp[11]) ? 4'b0100 : node25917;
														assign node25917 = (inp[9]) ? node25921 : node25918;
															assign node25918 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node25921 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node25925 = (inp[0]) ? node25931 : node25926;
														assign node25926 = (inp[1]) ? 4'b0001 : node25927;
															assign node25927 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node25931 = (inp[1]) ? 4'b0000 : node25932;
															assign node25932 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node25936 = (inp[4]) ? 4'b0100 : node25937;
													assign node25937 = (inp[11]) ? node25943 : node25938;
														assign node25938 = (inp[9]) ? node25940 : 4'b0000;
															assign node25940 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node25943 = (inp[1]) ? node25949 : node25944;
															assign node25944 = (inp[0]) ? 4'b0000 : node25945;
																assign node25945 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node25949 = (inp[9]) ? node25951 : 4'b0001;
																assign node25951 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node25955 = (inp[0]) ? node25977 : node25956;
												assign node25956 = (inp[4]) ? node25966 : node25957;
													assign node25957 = (inp[13]) ? node25959 : 4'b0100;
														assign node25959 = (inp[1]) ? node25963 : node25960;
															assign node25960 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node25963 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node25966 = (inp[13]) ? node25972 : node25967;
														assign node25967 = (inp[1]) ? 4'b0001 : node25968;
															assign node25968 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node25972 = (inp[9]) ? 4'b0101 : node25973;
															assign node25973 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node25977 = (inp[9]) ? node25993 : node25978;
													assign node25978 = (inp[1]) ? node25986 : node25979;
														assign node25979 = (inp[4]) ? node25983 : node25980;
															assign node25980 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node25983 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node25986 = (inp[13]) ? node25990 : node25987;
															assign node25987 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node25990 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node25993 = (inp[1]) ? node26005 : node25994;
														assign node25994 = (inp[4]) ? node26000 : node25995;
															assign node25995 = (inp[11]) ? 4'b0001 : node25996;
																assign node25996 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node26000 = (inp[13]) ? node26002 : 4'b0001;
																assign node26002 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node26005 = (inp[4]) ? node26009 : node26006;
															assign node26006 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node26009 = (inp[13]) ? 4'b0100 : 4'b0000;
										assign node26012 = (inp[13]) ? node26070 : node26013;
											assign node26013 = (inp[1]) ? node26047 : node26014;
												assign node26014 = (inp[4]) ? node26030 : node26015;
													assign node26015 = (inp[0]) ? node26021 : node26016;
														assign node26016 = (inp[11]) ? 4'b0101 : node26017;
															assign node26017 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node26021 = (inp[11]) ? node26025 : node26022;
															assign node26022 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node26025 = (inp[10]) ? 4'b0100 : node26026;
																assign node26026 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node26030 = (inp[11]) ? node26040 : node26031;
														assign node26031 = (inp[9]) ? 4'b0000 : node26032;
															assign node26032 = (inp[10]) ? node26036 : node26033;
																assign node26033 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node26036 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node26040 = (inp[9]) ? node26044 : node26041;
															assign node26041 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node26044 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node26047 = (inp[4]) ? node26051 : node26048;
													assign node26048 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node26051 = (inp[10]) ? node26061 : node26052;
														assign node26052 = (inp[0]) ? node26054 : 4'b0101;
															assign node26054 = (inp[11]) ? node26058 : node26055;
																assign node26055 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node26058 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node26061 = (inp[9]) ? node26067 : node26062;
															assign node26062 = (inp[11]) ? node26064 : 4'b0100;
																assign node26064 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node26067 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node26070 = (inp[1]) ? node26088 : node26071;
												assign node26071 = (inp[4]) ? node26077 : node26072;
													assign node26072 = (inp[0]) ? node26074 : 4'b0001;
														assign node26074 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node26077 = (inp[9]) ? node26085 : node26078;
														assign node26078 = (inp[10]) ? 4'b0101 : node26079;
															assign node26079 = (inp[0]) ? node26081 : 4'b0100;
																assign node26081 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node26085 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node26088 = (inp[4]) ? node26098 : node26089;
													assign node26089 = (inp[0]) ? node26091 : 4'b0100;
														assign node26091 = (inp[9]) ? node26093 : 4'b0101;
															assign node26093 = (inp[10]) ? 4'b0100 : node26094;
																assign node26094 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node26098 = (inp[10]) ? node26106 : node26099;
														assign node26099 = (inp[9]) ? node26101 : 4'b0001;
															assign node26101 = (inp[0]) ? node26103 : 4'b0000;
																assign node26103 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node26106 = (inp[9]) ? node26108 : 4'b0000;
															assign node26108 = (inp[0]) ? 4'b0000 : 4'b0001;
							assign node26111 = (inp[15]) ? node26501 : node26112;
								assign node26112 = (inp[4]) ? node26324 : node26113;
									assign node26113 = (inp[0]) ? node26229 : node26114;
										assign node26114 = (inp[1]) ? node26170 : node26115;
											assign node26115 = (inp[13]) ? node26135 : node26116;
												assign node26116 = (inp[11]) ? node26124 : node26117;
													assign node26117 = (inp[9]) ? 4'b0101 : node26118;
														assign node26118 = (inp[10]) ? 4'b0100 : node26119;
															assign node26119 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node26124 = (inp[2]) ? node26132 : node26125;
														assign node26125 = (inp[5]) ? 4'b0001 : node26126;
															assign node26126 = (inp[9]) ? 4'b0100 : node26127;
																assign node26127 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node26132 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node26135 = (inp[10]) ? node26155 : node26136;
													assign node26136 = (inp[11]) ? node26146 : node26137;
														assign node26137 = (inp[9]) ? node26141 : node26138;
															assign node26138 = (inp[5]) ? 4'b0000 : 4'b0101;
															assign node26141 = (inp[5]) ? 4'b0100 : node26142;
																assign node26142 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node26146 = (inp[2]) ? node26152 : node26147;
															assign node26147 = (inp[9]) ? node26149 : 4'b0100;
																assign node26149 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node26152 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node26155 = (inp[9]) ? node26165 : node26156;
														assign node26156 = (inp[2]) ? node26160 : node26157;
															assign node26157 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node26160 = (inp[5]) ? node26162 : 4'b0100;
																assign node26162 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node26165 = (inp[2]) ? 4'b0101 : node26166;
															assign node26166 = (inp[5]) ? 4'b0101 : 4'b0001;
											assign node26170 = (inp[13]) ? node26194 : node26171;
												assign node26171 = (inp[2]) ? node26179 : node26172;
													assign node26172 = (inp[11]) ? node26174 : 4'b0000;
														assign node26174 = (inp[5]) ? node26176 : 4'b0000;
															assign node26176 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node26179 = (inp[10]) ? node26189 : node26180;
														assign node26180 = (inp[5]) ? 4'b0100 : node26181;
															assign node26181 = (inp[11]) ? node26185 : node26182;
																assign node26182 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node26185 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node26189 = (inp[9]) ? 4'b0100 : node26190;
															assign node26190 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node26194 = (inp[2]) ? node26214 : node26195;
													assign node26195 = (inp[11]) ? node26201 : node26196;
														assign node26196 = (inp[10]) ? node26198 : 4'b0101;
															assign node26198 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node26201 = (inp[10]) ? node26209 : node26202;
															assign node26202 = (inp[5]) ? node26206 : node26203;
																assign node26203 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node26206 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node26209 = (inp[9]) ? 4'b0101 : node26210;
																assign node26210 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node26214 = (inp[9]) ? node26220 : node26215;
														assign node26215 = (inp[10]) ? node26217 : 4'b0001;
															assign node26217 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node26220 = (inp[10]) ? node26226 : node26221;
															assign node26221 = (inp[11]) ? node26223 : 4'b0000;
																assign node26223 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node26226 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node26229 = (inp[10]) ? node26275 : node26230;
											assign node26230 = (inp[11]) ? node26250 : node26231;
												assign node26231 = (inp[1]) ? node26237 : node26232;
													assign node26232 = (inp[5]) ? 4'b0001 : node26233;
														assign node26233 = (inp[2]) ? 4'b0101 : 4'b0000;
													assign node26237 = (inp[5]) ? node26243 : node26238;
														assign node26238 = (inp[9]) ? node26240 : 4'b0000;
															assign node26240 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node26243 = (inp[13]) ? node26247 : node26244;
															assign node26244 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node26247 = (inp[2]) ? 4'b0000 : 4'b0101;
												assign node26250 = (inp[5]) ? node26266 : node26251;
													assign node26251 = (inp[2]) ? node26257 : node26252;
														assign node26252 = (inp[13]) ? node26254 : 4'b0101;
															assign node26254 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node26257 = (inp[9]) ? node26259 : 4'b0101;
															assign node26259 = (inp[1]) ? node26263 : node26260;
																assign node26260 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node26263 = (inp[13]) ? 4'b0001 : 4'b0100;
													assign node26266 = (inp[2]) ? node26272 : node26267;
														assign node26267 = (inp[13]) ? 4'b0100 : node26268;
															assign node26268 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node26272 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node26275 = (inp[13]) ? node26289 : node26276;
												assign node26276 = (inp[2]) ? node26286 : node26277;
													assign node26277 = (inp[5]) ? node26281 : node26278;
														assign node26278 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node26281 = (inp[9]) ? 4'b0001 : node26282;
															assign node26282 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node26286 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node26289 = (inp[2]) ? node26305 : node26290;
													assign node26290 = (inp[1]) ? node26296 : node26291;
														assign node26291 = (inp[9]) ? 4'b0000 : node26292;
															assign node26292 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node26296 = (inp[9]) ? node26300 : node26297;
															assign node26297 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node26300 = (inp[5]) ? node26302 : 4'b0101;
																assign node26302 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node26305 = (inp[5]) ? node26317 : node26306;
														assign node26306 = (inp[1]) ? node26314 : node26307;
															assign node26307 = (inp[9]) ? node26311 : node26308;
																assign node26308 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node26311 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node26314 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node26317 = (inp[9]) ? node26319 : 4'b0000;
															assign node26319 = (inp[1]) ? node26321 : 4'b0001;
																assign node26321 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node26324 = (inp[10]) ? node26422 : node26325;
										assign node26325 = (inp[13]) ? node26375 : node26326;
											assign node26326 = (inp[2]) ? node26350 : node26327;
												assign node26327 = (inp[1]) ? node26341 : node26328;
													assign node26328 = (inp[5]) ? 4'b0110 : node26329;
														assign node26329 = (inp[9]) ? node26335 : node26330;
															assign node26330 = (inp[0]) ? node26332 : 4'b0010;
																assign node26332 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node26335 = (inp[0]) ? node26337 : 4'b0011;
																assign node26337 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node26341 = (inp[9]) ? node26347 : node26342;
														assign node26342 = (inp[0]) ? 4'b0111 : node26343;
															assign node26343 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node26347 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node26350 = (inp[5]) ? node26364 : node26351;
													assign node26351 = (inp[1]) ? node26357 : node26352;
														assign node26352 = (inp[11]) ? 4'b0111 : node26353;
															assign node26353 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node26357 = (inp[0]) ? node26361 : node26358;
															assign node26358 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node26361 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node26364 = (inp[9]) ? node26370 : node26365;
														assign node26365 = (inp[0]) ? node26367 : 4'b0010;
															assign node26367 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node26370 = (inp[1]) ? node26372 : 4'b0011;
															assign node26372 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node26375 = (inp[2]) ? node26397 : node26376;
												assign node26376 = (inp[1]) ? node26386 : node26377;
													assign node26377 = (inp[5]) ? node26381 : node26378;
														assign node26378 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node26381 = (inp[9]) ? node26383 : 4'b0010;
															assign node26383 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node26386 = (inp[9]) ? 4'b0010 : node26387;
														assign node26387 = (inp[5]) ? node26393 : node26388;
															assign node26388 = (inp[11]) ? node26390 : 4'b0010;
																assign node26390 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node26393 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node26397 = (inp[1]) ? node26413 : node26398;
													assign node26398 = (inp[5]) ? node26410 : node26399;
														assign node26399 = (inp[9]) ? node26405 : node26400;
															assign node26400 = (inp[0]) ? 4'b0010 : node26401;
																assign node26401 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26405 = (inp[11]) ? 4'b0011 : node26406;
																assign node26406 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node26410 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node26413 = (inp[11]) ? node26417 : node26414;
														assign node26414 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node26417 = (inp[9]) ? node26419 : 4'b0110;
															assign node26419 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node26422 = (inp[5]) ? node26464 : node26423;
											assign node26423 = (inp[13]) ? node26441 : node26424;
												assign node26424 = (inp[2]) ? node26432 : node26425;
													assign node26425 = (inp[1]) ? node26429 : node26426;
														assign node26426 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node26429 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node26432 = (inp[1]) ? 4'b0011 : node26433;
														assign node26433 = (inp[11]) ? 4'b0110 : node26434;
															assign node26434 = (inp[0]) ? 4'b0111 : node26435;
																assign node26435 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node26441 = (inp[9]) ? node26455 : node26442;
													assign node26442 = (inp[1]) ? node26450 : node26443;
														assign node26443 = (inp[2]) ? node26445 : 4'b0111;
															assign node26445 = (inp[0]) ? 4'b0011 : node26446;
																assign node26446 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node26450 = (inp[11]) ? node26452 : 4'b0111;
															assign node26452 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node26455 = (inp[0]) ? node26457 : 4'b0010;
														assign node26457 = (inp[11]) ? node26459 : 4'b0010;
															assign node26459 = (inp[1]) ? node26461 : 4'b0110;
																assign node26461 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node26464 = (inp[11]) ? node26482 : node26465;
												assign node26465 = (inp[13]) ? node26471 : node26466;
													assign node26466 = (inp[2]) ? 4'b0011 : node26467;
														assign node26467 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node26471 = (inp[2]) ? node26475 : node26472;
														assign node26472 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node26475 = (inp[9]) ? node26479 : node26476;
															assign node26476 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node26479 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node26482 = (inp[2]) ? node26492 : node26483;
													assign node26483 = (inp[13]) ? node26487 : node26484;
														assign node26484 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node26487 = (inp[9]) ? 4'b0011 : node26488;
															assign node26488 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node26492 = (inp[13]) ? node26496 : node26493;
														assign node26493 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node26496 = (inp[0]) ? node26498 : 4'b0111;
															assign node26498 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node26501 = (inp[0]) ? node26717 : node26502;
									assign node26502 = (inp[9]) ? node26604 : node26503;
										assign node26503 = (inp[13]) ? node26551 : node26504;
											assign node26504 = (inp[2]) ? node26526 : node26505;
												assign node26505 = (inp[5]) ? node26519 : node26506;
													assign node26506 = (inp[1]) ? node26514 : node26507;
														assign node26507 = (inp[10]) ? node26509 : 4'b0110;
															assign node26509 = (inp[11]) ? node26511 : 4'b0111;
																assign node26511 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node26514 = (inp[11]) ? node26516 : 4'b0011;
															assign node26516 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node26519 = (inp[11]) ? 4'b0010 : node26520;
														assign node26520 = (inp[10]) ? node26522 : 4'b0010;
															assign node26522 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node26526 = (inp[1]) ? node26540 : node26527;
													assign node26527 = (inp[5]) ? node26533 : node26528;
														assign node26528 = (inp[10]) ? node26530 : 4'b0010;
															assign node26530 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node26533 = (inp[10]) ? node26537 : node26534;
															assign node26534 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node26537 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node26540 = (inp[5]) ? 4'b0110 : node26541;
														assign node26541 = (inp[4]) ? node26543 : 4'b0110;
															assign node26543 = (inp[11]) ? node26547 : node26544;
																assign node26544 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node26547 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node26551 = (inp[2]) ? node26583 : node26552;
												assign node26552 = (inp[1]) ? node26568 : node26553;
													assign node26553 = (inp[5]) ? node26563 : node26554;
														assign node26554 = (inp[4]) ? node26560 : node26555;
															assign node26555 = (inp[10]) ? node26557 : 4'b0011;
																assign node26557 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26560 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node26563 = (inp[11]) ? node26565 : 4'b0111;
															assign node26565 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node26568 = (inp[10]) ? node26576 : node26569;
														assign node26569 = (inp[4]) ? node26571 : 4'b0111;
															assign node26571 = (inp[11]) ? 4'b0111 : node26572;
																assign node26572 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node26576 = (inp[11]) ? node26578 : 4'b0110;
															assign node26578 = (inp[4]) ? node26580 : 4'b0110;
																assign node26580 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node26583 = (inp[1]) ? node26597 : node26584;
													assign node26584 = (inp[5]) ? node26592 : node26585;
														assign node26585 = (inp[11]) ? node26587 : 4'b0111;
															assign node26587 = (inp[4]) ? node26589 : 4'b0111;
																assign node26589 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node26592 = (inp[11]) ? 4'b0011 : node26593;
															assign node26593 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node26597 = (inp[4]) ? node26601 : node26598;
														assign node26598 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node26601 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node26604 = (inp[1]) ? node26664 : node26605;
											assign node26605 = (inp[10]) ? node26639 : node26606;
												assign node26606 = (inp[4]) ? node26624 : node26607;
													assign node26607 = (inp[11]) ? node26615 : node26608;
														assign node26608 = (inp[5]) ? node26610 : 4'b0111;
															assign node26610 = (inp[2]) ? node26612 : 4'b0111;
																assign node26612 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node26615 = (inp[2]) ? 4'b0111 : node26616;
															assign node26616 = (inp[5]) ? node26620 : node26617;
																assign node26617 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node26620 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node26624 = (inp[13]) ? node26630 : node26625;
														assign node26625 = (inp[2]) ? node26627 : 4'b0010;
															assign node26627 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node26630 = (inp[11]) ? node26636 : node26631;
															assign node26631 = (inp[5]) ? 4'b0010 : node26632;
																assign node26632 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node26636 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node26639 = (inp[2]) ? node26651 : node26640;
													assign node26640 = (inp[11]) ? node26642 : 4'b0010;
														assign node26642 = (inp[13]) ? node26646 : node26643;
															assign node26643 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26646 = (inp[5]) ? node26648 : 4'b0011;
																assign node26648 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node26651 = (inp[11]) ? node26657 : node26652;
														assign node26652 = (inp[13]) ? 4'b0110 : node26653;
															assign node26653 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node26657 = (inp[13]) ? node26661 : node26658;
															assign node26658 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node26661 = (inp[5]) ? 4'b0010 : 4'b0111;
											assign node26664 = (inp[11]) ? node26690 : node26665;
												assign node26665 = (inp[5]) ? node26675 : node26666;
													assign node26666 = (inp[10]) ? 4'b0110 : node26667;
														assign node26667 = (inp[2]) ? node26671 : node26668;
															assign node26668 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node26671 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node26675 = (inp[10]) ? node26679 : node26676;
														assign node26676 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node26679 = (inp[4]) ? node26685 : node26680;
															assign node26680 = (inp[2]) ? 4'b0111 : node26681;
																assign node26681 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node26685 = (inp[13]) ? node26687 : 4'b0011;
																assign node26687 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node26690 = (inp[5]) ? node26710 : node26691;
													assign node26691 = (inp[4]) ? node26701 : node26692;
														assign node26692 = (inp[10]) ? node26698 : node26693;
															assign node26693 = (inp[2]) ? 4'b0011 : node26694;
																assign node26694 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node26698 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node26701 = (inp[2]) ? node26705 : node26702;
															assign node26702 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node26705 = (inp[13]) ? node26707 : 4'b0111;
																assign node26707 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node26710 = (inp[2]) ? node26714 : node26711;
														assign node26711 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node26714 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node26717 = (inp[11]) ? node26823 : node26718;
										assign node26718 = (inp[4]) ? node26774 : node26719;
											assign node26719 = (inp[2]) ? node26753 : node26720;
												assign node26720 = (inp[13]) ? node26734 : node26721;
													assign node26721 = (inp[5]) ? node26729 : node26722;
														assign node26722 = (inp[1]) ? node26726 : node26723;
															assign node26723 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node26726 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node26729 = (inp[10]) ? 4'b0011 : node26730;
															assign node26730 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node26734 = (inp[1]) ? node26746 : node26735;
														assign node26735 = (inp[5]) ? node26741 : node26736;
															assign node26736 = (inp[9]) ? node26738 : 4'b0010;
																assign node26738 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node26741 = (inp[10]) ? 4'b0110 : node26742;
																assign node26742 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node26746 = (inp[10]) ? node26750 : node26747;
															assign node26747 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node26750 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node26753 = (inp[13]) ? node26759 : node26754;
													assign node26754 = (inp[1]) ? 4'b0110 : node26755;
														assign node26755 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node26759 = (inp[1]) ? node26767 : node26760;
														assign node26760 = (inp[5]) ? node26762 : 4'b0110;
															assign node26762 = (inp[10]) ? node26764 : 4'b0010;
																assign node26764 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node26767 = (inp[9]) ? node26771 : node26768;
															assign node26768 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node26771 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node26774 = (inp[2]) ? node26800 : node26775;
												assign node26775 = (inp[1]) ? node26791 : node26776;
													assign node26776 = (inp[9]) ? node26784 : node26777;
														assign node26777 = (inp[10]) ? node26781 : node26778;
															assign node26778 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node26781 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node26784 = (inp[5]) ? node26788 : node26785;
															assign node26785 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node26788 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node26791 = (inp[5]) ? node26793 : 4'b0011;
														assign node26793 = (inp[10]) ? node26797 : node26794;
															assign node26794 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node26797 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node26800 = (inp[13]) ? node26808 : node26801;
													assign node26801 = (inp[5]) ? 4'b0111 : node26802;
														assign node26802 = (inp[1]) ? node26804 : 4'b0010;
															assign node26804 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node26808 = (inp[5]) ? node26818 : node26809;
														assign node26809 = (inp[1]) ? node26813 : node26810;
															assign node26810 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node26813 = (inp[10]) ? node26815 : 4'b0010;
																assign node26815 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node26818 = (inp[9]) ? node26820 : 4'b0011;
															assign node26820 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node26823 = (inp[10]) ? node26883 : node26824;
											assign node26824 = (inp[13]) ? node26854 : node26825;
												assign node26825 = (inp[2]) ? node26843 : node26826;
													assign node26826 = (inp[1]) ? node26834 : node26827;
														assign node26827 = (inp[5]) ? node26829 : 4'b0111;
															assign node26829 = (inp[9]) ? 4'b0011 : node26830;
																assign node26830 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node26834 = (inp[9]) ? node26838 : node26835;
															assign node26835 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node26838 = (inp[5]) ? node26840 : 4'b0010;
																assign node26840 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node26843 = (inp[5]) ? node26851 : node26844;
														assign node26844 = (inp[1]) ? 4'b0110 : node26845;
															assign node26845 = (inp[4]) ? 4'b0010 : node26846;
																assign node26846 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node26851 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node26854 = (inp[2]) ? node26872 : node26855;
													assign node26855 = (inp[1]) ? node26865 : node26856;
														assign node26856 = (inp[5]) ? node26860 : node26857;
															assign node26857 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node26860 = (inp[9]) ? 4'b0111 : node26861;
																assign node26861 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node26865 = (inp[5]) ? 4'b0110 : node26866;
															assign node26866 = (inp[9]) ? 4'b0111 : node26867;
																assign node26867 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node26872 = (inp[1]) ? node26878 : node26873;
														assign node26873 = (inp[5]) ? 4'b0011 : node26874;
															assign node26874 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node26878 = (inp[5]) ? node26880 : 4'b0011;
															assign node26880 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node26883 = (inp[1]) ? node26917 : node26884;
												assign node26884 = (inp[4]) ? node26902 : node26885;
													assign node26885 = (inp[13]) ? node26895 : node26886;
														assign node26886 = (inp[9]) ? node26890 : node26887;
															assign node26887 = (inp[2]) ? 4'b0011 : 4'b0110;
															assign node26890 = (inp[2]) ? node26892 : 4'b0011;
																assign node26892 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node26895 = (inp[9]) ? 4'b0010 : node26896;
															assign node26896 = (inp[2]) ? 4'b0110 : node26897;
																assign node26897 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node26902 = (inp[9]) ? node26914 : node26903;
														assign node26903 = (inp[5]) ? node26909 : node26904;
															assign node26904 = (inp[2]) ? 4'b0010 : node26905;
																assign node26905 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node26909 = (inp[2]) ? node26911 : 4'b0011;
																assign node26911 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node26914 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node26917 = (inp[2]) ? node26925 : node26918;
													assign node26918 = (inp[13]) ? node26920 : 4'b0010;
														assign node26920 = (inp[4]) ? 4'b0110 : node26921;
															assign node26921 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node26925 = (inp[13]) ? node26935 : node26926;
														assign node26926 = (inp[4]) ? node26932 : node26927;
															assign node26927 = (inp[5]) ? node26929 : 4'b0111;
																assign node26929 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node26932 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node26935 = (inp[4]) ? 4'b0010 : 4'b0011;
						assign node26938 = (inp[5]) ? node27342 : node26939;
							assign node26939 = (inp[9]) ? node27153 : node26940;
								assign node26940 = (inp[4]) ? node27094 : node26941;
									assign node26941 = (inp[1]) ? node26991 : node26942;
										assign node26942 = (inp[2]) ? node26968 : node26943;
											assign node26943 = (inp[15]) ? node26957 : node26944;
												assign node26944 = (inp[12]) ? node26950 : node26945;
													assign node26945 = (inp[13]) ? 4'b0110 : node26946;
														assign node26946 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node26950 = (inp[13]) ? node26954 : node26951;
														assign node26951 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node26954 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node26957 = (inp[12]) ? node26961 : node26958;
													assign node26958 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node26961 = (inp[0]) ? node26965 : node26962;
														assign node26962 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node26965 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node26968 = (inp[0]) ? node26980 : node26969;
												assign node26969 = (inp[13]) ? node26973 : node26970;
													assign node26970 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node26973 = (inp[12]) ? node26977 : node26974;
														assign node26974 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node26977 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node26980 = (inp[13]) ? node26984 : node26981;
													assign node26981 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node26984 = (inp[15]) ? node26988 : node26985;
														assign node26985 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node26988 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node26991 = (inp[11]) ? node27033 : node26992;
											assign node26992 = (inp[2]) ? node27012 : node26993;
												assign node26993 = (inp[12]) ? node27003 : node26994;
													assign node26994 = (inp[15]) ? 4'b0110 : node26995;
														assign node26995 = (inp[13]) ? node26999 : node26996;
															assign node26996 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node26999 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node27003 = (inp[13]) ? node27007 : node27004;
														assign node27004 = (inp[15]) ? 4'b0111 : 4'b0011;
														assign node27007 = (inp[15]) ? 4'b0011 : node27008;
															assign node27008 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node27012 = (inp[0]) ? node27024 : node27013;
													assign node27013 = (inp[12]) ? 4'b0111 : node27014;
														assign node27014 = (inp[10]) ? 4'b0111 : node27015;
															assign node27015 = (inp[15]) ? node27019 : node27016;
																assign node27016 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node27019 = (inp[13]) ? 4'b0111 : 4'b0010;
													assign node27024 = (inp[12]) ? node27028 : node27025;
														assign node27025 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node27028 = (inp[15]) ? 4'b0110 : node27029;
															assign node27029 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node27033 = (inp[2]) ? node27059 : node27034;
												assign node27034 = (inp[15]) ? node27046 : node27035;
													assign node27035 = (inp[13]) ? node27041 : node27036;
														assign node27036 = (inp[12]) ? 4'b0011 : node27037;
															assign node27037 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node27041 = (inp[12]) ? 4'b0110 : node27042;
															assign node27042 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node27046 = (inp[10]) ? node27052 : node27047;
														assign node27047 = (inp[12]) ? 4'b0010 : node27048;
															assign node27048 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node27052 = (inp[12]) ? node27056 : node27053;
															assign node27053 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node27056 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node27059 = (inp[10]) ? node27073 : node27060;
													assign node27060 = (inp[13]) ? node27066 : node27061;
														assign node27061 = (inp[15]) ? node27063 : 4'b0111;
															assign node27063 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node27066 = (inp[12]) ? node27070 : node27067;
															assign node27067 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node27070 = (inp[15]) ? 4'b0011 : 4'b0111;
													assign node27073 = (inp[13]) ? node27087 : node27074;
														assign node27074 = (inp[0]) ? node27082 : node27075;
															assign node27075 = (inp[15]) ? node27079 : node27076;
																assign node27076 = (inp[12]) ? 4'b0010 : 4'b0111;
																assign node27079 = (inp[12]) ? 4'b0111 : 4'b0010;
															assign node27082 = (inp[15]) ? node27084 : 4'b0110;
																assign node27084 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node27087 = (inp[15]) ? node27091 : node27088;
															assign node27088 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node27091 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node27094 = (inp[12]) ? node27138 : node27095;
										assign node27095 = (inp[15]) ? node27107 : node27096;
											assign node27096 = (inp[13]) ? node27102 : node27097;
												assign node27097 = (inp[0]) ? node27099 : 4'b0010;
													assign node27099 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node27102 = (inp[0]) ? 4'b0110 : node27103;
													assign node27103 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node27107 = (inp[13]) ? node27131 : node27108;
												assign node27108 = (inp[2]) ? node27122 : node27109;
													assign node27109 = (inp[10]) ? node27117 : node27110;
														assign node27110 = (inp[11]) ? node27112 : 4'b0110;
															assign node27112 = (inp[1]) ? 4'b0111 : node27113;
																assign node27113 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node27117 = (inp[11]) ? 4'b0110 : node27118;
															assign node27118 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node27122 = (inp[10]) ? node27126 : node27123;
														assign node27123 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node27126 = (inp[11]) ? node27128 : 4'b0111;
															assign node27128 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node27131 = (inp[0]) ? node27135 : node27132;
													assign node27132 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node27135 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node27138 = (inp[15]) ? node27150 : node27139;
											assign node27139 = (inp[13]) ? node27145 : node27140;
												assign node27140 = (inp[1]) ? node27142 : 4'b0010;
													assign node27142 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node27145 = (inp[1]) ? 4'b0110 : node27146;
													assign node27146 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node27150 = (inp[13]) ? 4'b0010 : 4'b0110;
								assign node27153 = (inp[4]) ? node27291 : node27154;
									assign node27154 = (inp[0]) ? node27238 : node27155;
										assign node27155 = (inp[2]) ? node27181 : node27156;
											assign node27156 = (inp[15]) ? node27170 : node27157;
												assign node27157 = (inp[12]) ? node27165 : node27158;
													assign node27158 = (inp[13]) ? node27162 : node27159;
														assign node27159 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node27162 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node27165 = (inp[13]) ? 4'b0010 : node27166;
														assign node27166 = (inp[1]) ? 4'b0010 : 4'b0111;
												assign node27170 = (inp[12]) ? node27178 : node27171;
													assign node27171 = (inp[13]) ? node27175 : node27172;
														assign node27172 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node27175 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node27178 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node27181 = (inp[10]) ? node27215 : node27182;
												assign node27182 = (inp[11]) ? node27198 : node27183;
													assign node27183 = (inp[15]) ? node27193 : node27184;
														assign node27184 = (inp[13]) ? 4'b0011 : node27185;
															assign node27185 = (inp[12]) ? node27189 : node27186;
																assign node27186 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node27189 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node27193 = (inp[12]) ? 4'b0010 : node27194;
															assign node27194 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node27198 = (inp[12]) ? node27206 : node27199;
														assign node27199 = (inp[1]) ? 4'b0011 : node27200;
															assign node27200 = (inp[13]) ? node27202 : 4'b0010;
																assign node27202 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node27206 = (inp[13]) ? node27208 : 4'b0110;
															assign node27208 = (inp[1]) ? node27212 : node27209;
																assign node27209 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node27212 = (inp[15]) ? 4'b0010 : 4'b0110;
												assign node27215 = (inp[12]) ? node27225 : node27216;
													assign node27216 = (inp[13]) ? node27220 : node27217;
														assign node27217 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node27220 = (inp[1]) ? 4'b0110 : node27221;
															assign node27221 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node27225 = (inp[15]) ? node27235 : node27226;
														assign node27226 = (inp[11]) ? node27230 : node27227;
															assign node27227 = (inp[1]) ? 4'b0110 : 4'b0011;
															assign node27230 = (inp[1]) ? 4'b0011 : node27231;
																assign node27231 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node27235 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node27238 = (inp[2]) ? node27264 : node27239;
											assign node27239 = (inp[12]) ? node27255 : node27240;
												assign node27240 = (inp[13]) ? node27248 : node27241;
													assign node27241 = (inp[15]) ? node27245 : node27242;
														assign node27242 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node27245 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node27248 = (inp[15]) ? node27252 : node27249;
														assign node27249 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node27252 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node27255 = (inp[13]) ? node27261 : node27256;
													assign node27256 = (inp[15]) ? 4'b0110 : node27257;
														assign node27257 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node27261 = (inp[15]) ? 4'b0010 : 4'b0110;
											assign node27264 = (inp[13]) ? node27278 : node27265;
												assign node27265 = (inp[12]) ? node27273 : node27266;
													assign node27266 = (inp[15]) ? node27270 : node27267;
														assign node27267 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node27270 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node27273 = (inp[1]) ? node27275 : 4'b0111;
														assign node27275 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node27278 = (inp[12]) ? node27286 : node27279;
													assign node27279 = (inp[15]) ? node27283 : node27280;
														assign node27280 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node27283 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node27286 = (inp[1]) ? node27288 : 4'b0010;
														assign node27288 = (inp[15]) ? 4'b0011 : 4'b0111;
									assign node27291 = (inp[12]) ? node27327 : node27292;
										assign node27292 = (inp[15]) ? node27304 : node27293;
											assign node27293 = (inp[13]) ? node27299 : node27294;
												assign node27294 = (inp[1]) ? 4'b0011 : node27295;
													assign node27295 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node27299 = (inp[0]) ? 4'b0111 : node27300;
													assign node27300 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node27304 = (inp[13]) ? node27320 : node27305;
												assign node27305 = (inp[10]) ? node27313 : node27306;
													assign node27306 = (inp[1]) ? node27310 : node27307;
														assign node27307 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node27310 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node27313 = (inp[11]) ? node27315 : 4'b0111;
														assign node27315 = (inp[1]) ? 4'b0110 : node27316;
															assign node27316 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node27320 = (inp[1]) ? node27324 : node27321;
													assign node27321 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node27324 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node27327 = (inp[15]) ? node27339 : node27328;
											assign node27328 = (inp[13]) ? node27334 : node27329;
												assign node27329 = (inp[0]) ? node27331 : 4'b0011;
													assign node27331 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node27334 = (inp[0]) ? 4'b0111 : node27335;
													assign node27335 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node27339 = (inp[13]) ? 4'b0011 : 4'b0111;
							assign node27342 = (inp[9]) ? node27488 : node27343;
								assign node27343 = (inp[4]) ? node27415 : node27344;
									assign node27344 = (inp[2]) ? node27376 : node27345;
										assign node27345 = (inp[12]) ? node27363 : node27346;
											assign node27346 = (inp[13]) ? node27352 : node27347;
												assign node27347 = (inp[1]) ? node27349 : 4'b0010;
													assign node27349 = (inp[15]) ? 4'b0011 : 4'b0110;
												assign node27352 = (inp[1]) ? node27360 : node27353;
													assign node27353 = (inp[15]) ? node27357 : node27354;
														assign node27354 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node27357 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node27360 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node27363 = (inp[15]) ? node27373 : node27364;
												assign node27364 = (inp[1]) ? node27368 : node27365;
													assign node27365 = (inp[13]) ? 4'b0011 : 4'b0110;
													assign node27368 = (inp[13]) ? 4'b0110 : node27369;
														assign node27369 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node27373 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node27376 = (inp[12]) ? node27402 : node27377;
											assign node27377 = (inp[13]) ? node27385 : node27378;
												assign node27378 = (inp[15]) ? node27382 : node27379;
													assign node27379 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node27382 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node27385 = (inp[15]) ? node27391 : node27386;
													assign node27386 = (inp[1]) ? 4'b0010 : node27387;
														assign node27387 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node27391 = (inp[10]) ? node27397 : node27392;
														assign node27392 = (inp[1]) ? node27394 : 4'b0110;
															assign node27394 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node27397 = (inp[0]) ? 4'b0110 : node27398;
															assign node27398 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node27402 = (inp[15]) ? node27412 : node27403;
												assign node27403 = (inp[1]) ? node27407 : node27404;
													assign node27404 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node27407 = (inp[13]) ? 4'b0111 : node27408;
														assign node27408 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node27412 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node27415 = (inp[12]) ? node27473 : node27416;
										assign node27416 = (inp[15]) ? node27428 : node27417;
											assign node27417 = (inp[13]) ? node27423 : node27418;
												assign node27418 = (inp[0]) ? node27420 : 4'b0011;
													assign node27420 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node27423 = (inp[0]) ? 4'b0111 : node27424;
													assign node27424 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node27428 = (inp[13]) ? node27444 : node27429;
												assign node27429 = (inp[2]) ? node27437 : node27430;
													assign node27430 = (inp[0]) ? node27434 : node27431;
														assign node27431 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node27434 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node27437 = (inp[11]) ? node27439 : 4'b0110;
														assign node27439 = (inp[0]) ? 4'b0111 : node27440;
															assign node27440 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node27444 = (inp[10]) ? node27456 : node27445;
													assign node27445 = (inp[11]) ? 4'b0010 : node27446;
														assign node27446 = (inp[2]) ? node27450 : node27447;
															assign node27447 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node27450 = (inp[1]) ? 4'b0010 : node27451;
																assign node27451 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node27456 = (inp[2]) ? node27462 : node27457;
														assign node27457 = (inp[0]) ? 4'b0010 : node27458;
															assign node27458 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node27462 = (inp[11]) ? node27468 : node27463;
															assign node27463 = (inp[1]) ? node27465 : 4'b0011;
																assign node27465 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node27468 = (inp[1]) ? 4'b0011 : node27469;
																assign node27469 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node27473 = (inp[15]) ? node27485 : node27474;
											assign node27474 = (inp[13]) ? node27480 : node27475;
												assign node27475 = (inp[1]) ? node27477 : 4'b0011;
													assign node27477 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node27480 = (inp[0]) ? 4'b0111 : node27481;
													assign node27481 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node27485 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node27488 = (inp[2]) ? node27638 : node27489;
									assign node27489 = (inp[4]) ? node27545 : node27490;
										assign node27490 = (inp[12]) ? node27512 : node27491;
											assign node27491 = (inp[13]) ? node27497 : node27492;
												assign node27492 = (inp[1]) ? node27494 : 4'b0011;
													assign node27494 = (inp[15]) ? 4'b0010 : 4'b0111;
												assign node27497 = (inp[15]) ? node27501 : node27498;
													assign node27498 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node27501 = (inp[10]) ? node27503 : 4'b0111;
														assign node27503 = (inp[11]) ? node27505 : 4'b0110;
															assign node27505 = (inp[1]) ? node27509 : node27506;
																assign node27506 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node27509 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node27512 = (inp[15]) ? node27542 : node27513;
												assign node27513 = (inp[0]) ? node27521 : node27514;
													assign node27514 = (inp[1]) ? node27518 : node27515;
														assign node27515 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node27518 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node27521 = (inp[10]) ? node27529 : node27522;
														assign node27522 = (inp[13]) ? node27526 : node27523;
															assign node27523 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node27526 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node27529 = (inp[11]) ? node27535 : node27530;
															assign node27530 = (inp[1]) ? node27532 : 4'b0111;
																assign node27532 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node27535 = (inp[13]) ? node27539 : node27536;
																assign node27536 = (inp[1]) ? 4'b0010 : 4'b0111;
																assign node27539 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node27542 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node27545 = (inp[10]) ? node27589 : node27546;
											assign node27546 = (inp[0]) ? node27572 : node27547;
												assign node27547 = (inp[1]) ? node27565 : node27548;
													assign node27548 = (inp[11]) ? node27554 : node27549;
														assign node27549 = (inp[15]) ? node27551 : 4'b0010;
															assign node27551 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node27554 = (inp[12]) ? node27562 : node27555;
															assign node27555 = (inp[13]) ? node27559 : node27556;
																assign node27556 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node27559 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node27562 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node27565 = (inp[15]) ? node27569 : node27566;
														assign node27566 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node27569 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node27572 = (inp[13]) ? node27582 : node27573;
													assign node27573 = (inp[15]) ? 4'b0110 : node27574;
														assign node27574 = (inp[12]) ? node27578 : node27575;
															assign node27575 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node27578 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node27582 = (inp[15]) ? node27584 : 4'b0110;
														assign node27584 = (inp[12]) ? 4'b0010 : node27585;
															assign node27585 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node27589 = (inp[12]) ? node27615 : node27590;
												assign node27590 = (inp[0]) ? node27598 : node27591;
													assign node27591 = (inp[13]) ? node27595 : node27592;
														assign node27592 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node27595 = (inp[11]) ? 4'b0011 : 4'b0111;
													assign node27598 = (inp[1]) ? node27610 : node27599;
														assign node27599 = (inp[11]) ? node27605 : node27600;
															assign node27600 = (inp[15]) ? node27602 : 4'b0011;
																assign node27602 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node27605 = (inp[13]) ? 4'b0110 : node27606;
																assign node27606 = (inp[15]) ? 4'b0111 : 4'b0011;
														assign node27610 = (inp[15]) ? node27612 : 4'b0110;
															assign node27612 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node27615 = (inp[0]) ? node27623 : node27616;
													assign node27616 = (inp[13]) ? node27620 : node27617;
														assign node27617 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node27620 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node27623 = (inp[1]) ? node27635 : node27624;
														assign node27624 = (inp[11]) ? node27630 : node27625;
															assign node27625 = (inp[15]) ? node27627 : 4'b0010;
																assign node27627 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node27630 = (inp[13]) ? node27632 : 4'b0110;
																assign node27632 = (inp[15]) ? 4'b0010 : 4'b0110;
														assign node27635 = (inp[13]) ? 4'b0110 : 4'b0011;
									assign node27638 = (inp[12]) ? node27698 : node27639;
										assign node27639 = (inp[13]) ? node27665 : node27640;
											assign node27640 = (inp[15]) ? node27650 : node27641;
												assign node27641 = (inp[4]) ? node27645 : node27642;
													assign node27642 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node27645 = (inp[0]) ? node27647 : 4'b0010;
														assign node27647 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node27650 = (inp[4]) ? node27654 : node27651;
													assign node27651 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node27654 = (inp[11]) ? node27660 : node27655;
														assign node27655 = (inp[1]) ? node27657 : 4'b0110;
															assign node27657 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node27660 = (inp[0]) ? node27662 : 4'b0111;
															assign node27662 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node27665 = (inp[4]) ? node27683 : node27666;
												assign node27666 = (inp[1]) ? node27678 : node27667;
													assign node27667 = (inp[11]) ? node27673 : node27668;
														assign node27668 = (inp[15]) ? 4'b0111 : node27669;
															assign node27669 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node27673 = (inp[10]) ? 4'b0110 : node27674;
															assign node27674 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node27678 = (inp[15]) ? node27680 : 4'b0011;
														assign node27680 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node27683 = (inp[15]) ? node27689 : node27684;
													assign node27684 = (inp[10]) ? 4'b0110 : node27685;
														assign node27685 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node27689 = (inp[10]) ? node27693 : node27690;
														assign node27690 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node27693 = (inp[0]) ? 4'b0011 : node27694;
															assign node27694 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node27698 = (inp[13]) ? node27710 : node27699;
											assign node27699 = (inp[15]) ? 4'b0110 : node27700;
												assign node27700 = (inp[4]) ? node27704 : node27701;
													assign node27701 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node27704 = (inp[1]) ? node27706 : 4'b0010;
														assign node27706 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node27710 = (inp[15]) ? 4'b0010 : node27711;
												assign node27711 = (inp[1]) ? 4'b0110 : node27712;
													assign node27712 = (inp[4]) ? node27714 : 4'b0011;
														assign node27714 = (inp[0]) ? 4'b0110 : 4'b0111;
					assign node27719 = (inp[6]) ? node29257 : node27720;
						assign node27720 = (inp[12]) ? node28486 : node27721;
							assign node27721 = (inp[15]) ? node28069 : node27722;
								assign node27722 = (inp[4]) ? node27910 : node27723;
									assign node27723 = (inp[11]) ? node27801 : node27724;
										assign node27724 = (inp[1]) ? node27756 : node27725;
											assign node27725 = (inp[2]) ? node27743 : node27726;
												assign node27726 = (inp[9]) ? node27734 : node27727;
													assign node27727 = (inp[10]) ? node27729 : 4'b0001;
														assign node27729 = (inp[5]) ? 4'b0100 : node27730;
															assign node27730 = (inp[0]) ? 4'b0001 : 4'b0101;
													assign node27734 = (inp[13]) ? node27740 : node27735;
														assign node27735 = (inp[10]) ? node27737 : 4'b0000;
															assign node27737 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node27740 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node27743 = (inp[13]) ? node27747 : node27744;
													assign node27744 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node27747 = (inp[5]) ? 4'b0000 : node27748;
														assign node27748 = (inp[0]) ? 4'b0100 : node27749;
															assign node27749 = (inp[10]) ? 4'b0101 : node27750;
																assign node27750 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node27756 = (inp[10]) ? node27774 : node27757;
												assign node27757 = (inp[2]) ? node27767 : node27758;
													assign node27758 = (inp[13]) ? node27764 : node27759;
														assign node27759 = (inp[0]) ? 4'b0000 : node27760;
															assign node27760 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node27764 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node27767 = (inp[13]) ? node27771 : node27768;
														assign node27768 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node27771 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node27774 = (inp[5]) ? node27792 : node27775;
													assign node27775 = (inp[9]) ? node27785 : node27776;
														assign node27776 = (inp[0]) ? node27778 : 4'b0100;
															assign node27778 = (inp[13]) ? node27782 : node27779;
																assign node27779 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node27782 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node27785 = (inp[13]) ? node27789 : node27786;
															assign node27786 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node27789 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node27792 = (inp[9]) ? node27798 : node27793;
														assign node27793 = (inp[0]) ? 4'b0000 : node27794;
															assign node27794 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node27798 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node27801 = (inp[10]) ? node27865 : node27802;
											assign node27802 = (inp[1]) ? node27836 : node27803;
												assign node27803 = (inp[13]) ? node27821 : node27804;
													assign node27804 = (inp[2]) ? node27814 : node27805;
														assign node27805 = (inp[5]) ? node27809 : node27806;
															assign node27806 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node27809 = (inp[0]) ? node27811 : 4'b0000;
																assign node27811 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node27814 = (inp[5]) ? node27818 : node27815;
															assign node27815 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node27818 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node27821 = (inp[0]) ? node27827 : node27822;
														assign node27822 = (inp[2]) ? node27824 : 4'b0001;
															assign node27824 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node27827 = (inp[5]) ? node27833 : node27828;
															assign node27828 = (inp[9]) ? 4'b0101 : node27829;
																assign node27829 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node27833 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node27836 = (inp[5]) ? node27846 : node27837;
													assign node27837 = (inp[9]) ? 4'b0101 : node27838;
														assign node27838 = (inp[13]) ? node27842 : node27839;
															assign node27839 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node27842 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node27846 = (inp[0]) ? node27862 : node27847;
														assign node27847 = (inp[2]) ? node27855 : node27848;
															assign node27848 = (inp[13]) ? node27852 : node27849;
																assign node27849 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node27852 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node27855 = (inp[13]) ? node27859 : node27856;
																assign node27856 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node27859 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node27862 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node27865 = (inp[0]) ? node27887 : node27866;
												assign node27866 = (inp[5]) ? node27882 : node27867;
													assign node27867 = (inp[1]) ? node27871 : node27868;
														assign node27868 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node27871 = (inp[13]) ? node27875 : node27872;
															assign node27872 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node27875 = (inp[2]) ? node27879 : node27876;
																assign node27876 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node27879 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node27882 = (inp[9]) ? 4'b0101 : node27883;
														assign node27883 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node27887 = (inp[1]) ? node27897 : node27888;
													assign node27888 = (inp[5]) ? node27890 : 4'b0101;
														assign node27890 = (inp[13]) ? 4'b0001 : node27891;
															assign node27891 = (inp[2]) ? 4'b0100 : node27892;
																assign node27892 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node27897 = (inp[2]) ? node27901 : node27898;
														assign node27898 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node27901 = (inp[13]) ? node27905 : node27902;
															assign node27902 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node27905 = (inp[9]) ? 4'b0000 : node27906;
																assign node27906 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node27910 = (inp[10]) ? node27994 : node27911;
										assign node27911 = (inp[9]) ? node27951 : node27912;
											assign node27912 = (inp[2]) ? node27932 : node27913;
												assign node27913 = (inp[13]) ? node27925 : node27914;
													assign node27914 = (inp[1]) ? 4'b0010 : node27915;
														assign node27915 = (inp[5]) ? node27921 : node27916;
															assign node27916 = (inp[11]) ? 4'b0111 : node27917;
																assign node27917 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node27921 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node27925 = (inp[1]) ? node27929 : node27926;
														assign node27926 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node27929 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node27932 = (inp[13]) ? node27938 : node27933;
													assign node27933 = (inp[11]) ? node27935 : 4'b0010;
														assign node27935 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node27938 = (inp[5]) ? node27942 : node27939;
														assign node27939 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node27942 = (inp[1]) ? node27948 : node27943;
															assign node27943 = (inp[0]) ? node27945 : 4'b0010;
																assign node27945 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node27948 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node27951 = (inp[13]) ? node27973 : node27952;
												assign node27952 = (inp[2]) ? node27962 : node27953;
													assign node27953 = (inp[0]) ? node27955 : 4'b0111;
														assign node27955 = (inp[1]) ? node27959 : node27956;
															assign node27956 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node27959 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node27962 = (inp[5]) ? node27968 : node27963;
														assign node27963 = (inp[1]) ? 4'b0110 : node27964;
															assign node27964 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node27968 = (inp[0]) ? node27970 : 4'b0110;
															assign node27970 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node27973 = (inp[2]) ? node27985 : node27974;
													assign node27974 = (inp[5]) ? node27978 : node27975;
														assign node27975 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node27978 = (inp[1]) ? node27982 : node27979;
															assign node27979 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node27982 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node27985 = (inp[5]) ? node27989 : node27986;
														assign node27986 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node27989 = (inp[11]) ? node27991 : 4'b0011;
															assign node27991 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node27994 = (inp[2]) ? node28040 : node27995;
											assign node27995 = (inp[13]) ? node28023 : node27996;
												assign node27996 = (inp[5]) ? node28006 : node27997;
													assign node27997 = (inp[1]) ? node28003 : node27998;
														assign node27998 = (inp[9]) ? node28000 : 4'b0110;
															assign node28000 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node28003 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node28006 = (inp[0]) ? node28018 : node28007;
														assign node28007 = (inp[9]) ? node28013 : node28008;
															assign node28008 = (inp[1]) ? 4'b0011 : node28009;
																assign node28009 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node28013 = (inp[1]) ? 4'b0010 : node28014;
																assign node28014 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node28018 = (inp[9]) ? node28020 : 4'b0010;
															assign node28020 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node28023 = (inp[5]) ? node28031 : node28024;
													assign node28024 = (inp[1]) ? node28026 : 4'b0011;
														assign node28026 = (inp[9]) ? node28028 : 4'b0111;
															assign node28028 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node28031 = (inp[1]) ? 4'b0110 : node28032;
														assign node28032 = (inp[9]) ? 4'b0110 : node28033;
															assign node28033 = (inp[0]) ? node28035 : 4'b0111;
																assign node28035 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node28040 = (inp[1]) ? node28056 : node28041;
												assign node28041 = (inp[9]) ? node28049 : node28042;
													assign node28042 = (inp[13]) ? node28046 : node28043;
														assign node28043 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node28046 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node28049 = (inp[13]) ? 4'b0110 : node28050;
														assign node28050 = (inp[5]) ? node28052 : 4'b0011;
															assign node28052 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node28056 = (inp[13]) ? node28066 : node28057;
													assign node28057 = (inp[0]) ? 4'b0111 : node28058;
														assign node28058 = (inp[11]) ? node28062 : node28059;
															assign node28059 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node28062 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node28066 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node28069 = (inp[0]) ? node28281 : node28070;
									assign node28070 = (inp[11]) ? node28162 : node28071;
										assign node28071 = (inp[5]) ? node28115 : node28072;
											assign node28072 = (inp[4]) ? node28086 : node28073;
												assign node28073 = (inp[1]) ? 4'b0110 : node28074;
													assign node28074 = (inp[2]) ? node28082 : node28075;
														assign node28075 = (inp[13]) ? 4'b0110 : node28076;
															assign node28076 = (inp[10]) ? node28078 : 4'b0010;
																assign node28078 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node28082 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node28086 = (inp[2]) ? node28098 : node28087;
													assign node28087 = (inp[10]) ? node28089 : 4'b0010;
														assign node28089 = (inp[9]) ? node28095 : node28090;
															assign node28090 = (inp[1]) ? node28092 : 4'b0111;
																assign node28092 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node28095 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node28098 = (inp[10]) ? node28108 : node28099;
														assign node28099 = (inp[1]) ? node28105 : node28100;
															assign node28100 = (inp[13]) ? node28102 : 4'b0011;
																assign node28102 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node28105 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node28108 = (inp[9]) ? node28110 : 4'b0111;
															assign node28110 = (inp[1]) ? 4'b0111 : node28111;
																assign node28111 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node28115 = (inp[4]) ? node28145 : node28116;
												assign node28116 = (inp[1]) ? node28132 : node28117;
													assign node28117 = (inp[9]) ? node28123 : node28118;
														assign node28118 = (inp[13]) ? 4'b0110 : node28119;
															assign node28119 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node28123 = (inp[2]) ? node28129 : node28124;
															assign node28124 = (inp[10]) ? node28126 : 4'b0110;
																assign node28126 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node28129 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node28132 = (inp[9]) ? 4'b0110 : node28133;
														assign node28133 = (inp[13]) ? node28141 : node28134;
															assign node28134 = (inp[2]) ? node28138 : node28135;
																assign node28135 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node28138 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node28141 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node28145 = (inp[10]) ? node28153 : node28146;
													assign node28146 = (inp[1]) ? node28148 : 4'b0110;
														assign node28148 = (inp[2]) ? 4'b0110 : node28149;
															assign node28149 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node28153 = (inp[13]) ? 4'b0011 : node28154;
														assign node28154 = (inp[2]) ? node28158 : node28155;
															assign node28155 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node28158 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node28162 = (inp[1]) ? node28226 : node28163;
											assign node28163 = (inp[5]) ? node28193 : node28164;
												assign node28164 = (inp[2]) ? node28180 : node28165;
													assign node28165 = (inp[9]) ? node28171 : node28166;
														assign node28166 = (inp[4]) ? node28168 : 4'b0111;
															assign node28168 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node28171 = (inp[4]) ? node28175 : node28172;
															assign node28172 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node28175 = (inp[10]) ? 4'b0110 : node28176;
																assign node28176 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node28180 = (inp[4]) ? node28184 : node28181;
														assign node28181 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node28184 = (inp[13]) ? node28186 : 4'b0011;
															assign node28186 = (inp[10]) ? node28190 : node28187;
																assign node28187 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node28190 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node28193 = (inp[10]) ? node28211 : node28194;
													assign node28194 = (inp[9]) ? node28198 : node28195;
														assign node28195 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node28198 = (inp[13]) ? node28206 : node28199;
															assign node28199 = (inp[4]) ? node28203 : node28200;
																assign node28200 = (inp[2]) ? 4'b0011 : 4'b0110;
																assign node28203 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node28206 = (inp[4]) ? 4'b0110 : node28207;
																assign node28207 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node28211 = (inp[9]) ? node28217 : node28212;
														assign node28212 = (inp[4]) ? 4'b0110 : node28213;
															assign node28213 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node28217 = (inp[4]) ? 4'b0111 : node28218;
															assign node28218 = (inp[13]) ? node28222 : node28219;
																assign node28219 = (inp[2]) ? 4'b0010 : 4'b0111;
																assign node28222 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node28226 = (inp[13]) ? node28256 : node28227;
												assign node28227 = (inp[4]) ? node28243 : node28228;
													assign node28228 = (inp[2]) ? node28234 : node28229;
														assign node28229 = (inp[10]) ? 4'b0111 : node28230;
															assign node28230 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node28234 = (inp[5]) ? node28240 : node28235;
															assign node28235 = (inp[9]) ? 4'b0010 : node28236;
																assign node28236 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node28240 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node28243 = (inp[2]) ? node28249 : node28244;
														assign node28244 = (inp[9]) ? node28246 : 4'b0011;
															assign node28246 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node28249 = (inp[9]) ? node28253 : node28250;
															assign node28250 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node28253 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node28256 = (inp[4]) ? node28270 : node28257;
													assign node28257 = (inp[2]) ? node28261 : node28258;
														assign node28258 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node28261 = (inp[9]) ? node28263 : 4'b0110;
															assign node28263 = (inp[10]) ? node28267 : node28264;
																assign node28264 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node28267 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node28270 = (inp[2]) ? node28276 : node28271;
														assign node28271 = (inp[10]) ? node28273 : 4'b0110;
															assign node28273 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node28276 = (inp[9]) ? 4'b0010 : node28277;
															assign node28277 = (inp[10]) ? 4'b0011 : 4'b0010;
									assign node28281 = (inp[5]) ? node28381 : node28282;
										assign node28282 = (inp[1]) ? node28344 : node28283;
											assign node28283 = (inp[10]) ? node28319 : node28284;
												assign node28284 = (inp[9]) ? node28304 : node28285;
													assign node28285 = (inp[11]) ? node28295 : node28286;
														assign node28286 = (inp[13]) ? node28288 : 4'b0110;
															assign node28288 = (inp[2]) ? node28292 : node28289;
																assign node28289 = (inp[4]) ? 4'b0010 : 4'b0111;
																assign node28292 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node28295 = (inp[2]) ? node28301 : node28296;
															assign node28296 = (inp[4]) ? 4'b0011 : node28297;
																assign node28297 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node28301 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node28304 = (inp[11]) ? node28308 : node28305;
														assign node28305 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node28308 = (inp[4]) ? node28312 : node28309;
															assign node28309 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node28312 = (inp[2]) ? node28316 : node28313;
																assign node28313 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node28316 = (inp[13]) ? 4'b0110 : 4'b0010;
												assign node28319 = (inp[4]) ? node28335 : node28320;
													assign node28320 = (inp[11]) ? node28330 : node28321;
														assign node28321 = (inp[9]) ? node28323 : 4'b0110;
															assign node28323 = (inp[2]) ? node28327 : node28324;
																assign node28324 = (inp[13]) ? 4'b0111 : 4'b0010;
																assign node28327 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node28330 = (inp[13]) ? node28332 : 4'b0111;
															assign node28332 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node28335 = (inp[11]) ? node28339 : node28336;
														assign node28336 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node28339 = (inp[2]) ? node28341 : 4'b0010;
															assign node28341 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node28344 = (inp[4]) ? node28362 : node28345;
												assign node28345 = (inp[2]) ? node28357 : node28346;
													assign node28346 = (inp[13]) ? node28350 : node28347;
														assign node28347 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node28350 = (inp[11]) ? node28352 : 4'b0011;
															assign node28352 = (inp[10]) ? 4'b0010 : node28353;
																assign node28353 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node28357 = (inp[13]) ? node28359 : 4'b0010;
														assign node28359 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node28362 = (inp[13]) ? node28370 : node28363;
													assign node28363 = (inp[2]) ? node28365 : 4'b0011;
														assign node28365 = (inp[9]) ? 4'b0111 : node28366;
															assign node28366 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node28370 = (inp[2]) ? node28378 : node28371;
														assign node28371 = (inp[10]) ? node28375 : node28372;
															assign node28372 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node28375 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node28378 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node28381 = (inp[4]) ? node28449 : node28382;
											assign node28382 = (inp[13]) ? node28414 : node28383;
												assign node28383 = (inp[2]) ? node28399 : node28384;
													assign node28384 = (inp[1]) ? node28392 : node28385;
														assign node28385 = (inp[10]) ? node28389 : node28386;
															assign node28386 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node28389 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node28392 = (inp[11]) ? 4'b0110 : node28393;
															assign node28393 = (inp[10]) ? node28395 : 4'b0110;
																assign node28395 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node28399 = (inp[9]) ? node28401 : 4'b0010;
														assign node28401 = (inp[1]) ? node28409 : node28402;
															assign node28402 = (inp[11]) ? node28406 : node28403;
																assign node28403 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node28406 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node28409 = (inp[10]) ? node28411 : 4'b0010;
																assign node28411 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node28414 = (inp[2]) ? node28440 : node28415;
													assign node28415 = (inp[9]) ? node28425 : node28416;
														assign node28416 = (inp[1]) ? node28418 : 4'b0010;
															assign node28418 = (inp[10]) ? node28422 : node28419;
																assign node28419 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node28422 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node28425 = (inp[10]) ? node28433 : node28426;
															assign node28426 = (inp[11]) ? node28430 : node28427;
																assign node28427 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node28430 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node28433 = (inp[11]) ? node28437 : node28434;
																assign node28434 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node28437 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node28440 = (inp[1]) ? node28442 : 4'b0111;
														assign node28442 = (inp[10]) ? node28446 : node28443;
															assign node28443 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node28446 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node28449 = (inp[2]) ? node28469 : node28450;
												assign node28450 = (inp[13]) ? node28462 : node28451;
													assign node28451 = (inp[1]) ? node28455 : node28452;
														assign node28452 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node28455 = (inp[9]) ? node28457 : 4'b0010;
															assign node28457 = (inp[10]) ? node28459 : 4'b0011;
																assign node28459 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node28462 = (inp[1]) ? 4'b0110 : node28463;
														assign node28463 = (inp[10]) ? node28465 : 4'b0111;
															assign node28465 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node28469 = (inp[13]) ? node28471 : 4'b0110;
													assign node28471 = (inp[10]) ? node28479 : node28472;
														assign node28472 = (inp[9]) ? node28476 : node28473;
															assign node28473 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node28476 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node28479 = (inp[9]) ? node28483 : node28480;
															assign node28480 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node28483 = (inp[1]) ? 4'b0010 : 4'b0011;
							assign node28486 = (inp[15]) ? node28846 : node28487;
								assign node28487 = (inp[4]) ? node28653 : node28488;
									assign node28488 = (inp[13]) ? node28574 : node28489;
										assign node28489 = (inp[2]) ? node28531 : node28490;
											assign node28490 = (inp[1]) ? node28520 : node28491;
												assign node28491 = (inp[0]) ? node28509 : node28492;
													assign node28492 = (inp[11]) ? node28498 : node28493;
														assign node28493 = (inp[10]) ? node28495 : 4'b0111;
															assign node28495 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node28498 = (inp[5]) ? node28504 : node28499;
															assign node28499 = (inp[9]) ? node28501 : 4'b0110;
																assign node28501 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node28504 = (inp[10]) ? 4'b0111 : node28505;
																assign node28505 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node28509 = (inp[11]) ? node28515 : node28510;
														assign node28510 = (inp[5]) ? node28512 : 4'b0110;
															assign node28512 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node28515 = (inp[9]) ? 4'b0110 : node28516;
															assign node28516 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node28520 = (inp[5]) ? node28528 : node28521;
													assign node28521 = (inp[11]) ? node28523 : 4'b0111;
														assign node28523 = (inp[10]) ? node28525 : 4'b0110;
															assign node28525 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node28528 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node28531 = (inp[1]) ? node28551 : node28532;
												assign node28532 = (inp[0]) ? node28542 : node28533;
													assign node28533 = (inp[11]) ? 4'b0010 : node28534;
														assign node28534 = (inp[5]) ? node28536 : 4'b0010;
															assign node28536 = (inp[9]) ? node28538 : 4'b0011;
																assign node28538 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node28542 = (inp[11]) ? node28546 : node28543;
														assign node28543 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node28546 = (inp[9]) ? node28548 : 4'b0011;
															assign node28548 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node28551 = (inp[5]) ? node28561 : node28552;
													assign node28552 = (inp[11]) ? node28554 : 4'b0010;
														assign node28554 = (inp[10]) ? node28558 : node28555;
															assign node28555 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node28558 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node28561 = (inp[9]) ? node28567 : node28562;
														assign node28562 = (inp[10]) ? 4'b0110 : node28563;
															assign node28563 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node28567 = (inp[11]) ? node28571 : node28568;
															assign node28568 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node28571 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node28574 = (inp[2]) ? node28614 : node28575;
											assign node28575 = (inp[5]) ? node28591 : node28576;
												assign node28576 = (inp[9]) ? node28582 : node28577;
													assign node28577 = (inp[0]) ? node28579 : 4'b0011;
														assign node28579 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node28582 = (inp[10]) ? node28588 : node28583;
														assign node28583 = (inp[11]) ? node28585 : 4'b0010;
															assign node28585 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node28588 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node28591 = (inp[1]) ? node28601 : node28592;
													assign node28592 = (inp[9]) ? node28594 : 4'b0011;
														assign node28594 = (inp[11]) ? node28598 : node28595;
															assign node28595 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node28598 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node28601 = (inp[10]) ? node28609 : node28602;
														assign node28602 = (inp[0]) ? 4'b0111 : node28603;
															assign node28603 = (inp[11]) ? 4'b0110 : node28604;
																assign node28604 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node28609 = (inp[9]) ? 4'b0111 : node28610;
															assign node28610 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node28614 = (inp[1]) ? node28628 : node28615;
												assign node28615 = (inp[10]) ? node28623 : node28616;
													assign node28616 = (inp[9]) ? 4'b0110 : node28617;
														assign node28617 = (inp[0]) ? node28619 : 4'b0111;
															assign node28619 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node28623 = (inp[9]) ? node28625 : 4'b0110;
														assign node28625 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node28628 = (inp[5]) ? node28636 : node28629;
													assign node28629 = (inp[9]) ? 4'b0110 : node28630;
														assign node28630 = (inp[10]) ? node28632 : 4'b0111;
															assign node28632 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node28636 = (inp[9]) ? node28646 : node28637;
														assign node28637 = (inp[10]) ? node28641 : node28638;
															assign node28638 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node28641 = (inp[11]) ? 4'b0011 : node28642;
																assign node28642 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node28646 = (inp[0]) ? 4'b0011 : node28647;
															assign node28647 = (inp[10]) ? 4'b0011 : node28648;
																assign node28648 = (inp[11]) ? 4'b0011 : 4'b0010;
									assign node28653 = (inp[0]) ? node28755 : node28654;
										assign node28654 = (inp[2]) ? node28698 : node28655;
											assign node28655 = (inp[13]) ? node28675 : node28656;
												assign node28656 = (inp[1]) ? node28668 : node28657;
													assign node28657 = (inp[5]) ? node28665 : node28658;
														assign node28658 = (inp[11]) ? node28660 : 4'b0100;
															assign node28660 = (inp[9]) ? node28662 : 4'b0101;
																assign node28662 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node28665 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node28668 = (inp[9]) ? node28672 : node28669;
														assign node28669 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node28672 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node28675 = (inp[1]) ? node28691 : node28676;
													assign node28676 = (inp[5]) ? node28686 : node28677;
														assign node28677 = (inp[9]) ? node28679 : 4'b0001;
															assign node28679 = (inp[10]) ? node28683 : node28680;
																assign node28680 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node28683 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node28686 = (inp[9]) ? 4'b0101 : node28687;
															assign node28687 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node28691 = (inp[9]) ? 4'b0100 : node28692;
														assign node28692 = (inp[10]) ? 4'b0100 : node28693;
															assign node28693 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node28698 = (inp[13]) ? node28730 : node28699;
												assign node28699 = (inp[1]) ? node28711 : node28700;
													assign node28700 = (inp[5]) ? node28706 : node28701;
														assign node28701 = (inp[9]) ? 4'b0000 : node28702;
															assign node28702 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node28706 = (inp[9]) ? node28708 : 4'b0100;
															assign node28708 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node28711 = (inp[9]) ? node28719 : node28712;
														assign node28712 = (inp[5]) ? node28714 : 4'b0100;
															assign node28714 = (inp[10]) ? 4'b0101 : node28715;
																assign node28715 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node28719 = (inp[5]) ? node28725 : node28720;
															assign node28720 = (inp[10]) ? 4'b0101 : node28721;
																assign node28721 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node28725 = (inp[11]) ? 4'b0100 : node28726;
																assign node28726 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node28730 = (inp[1]) ? node28742 : node28731;
													assign node28731 = (inp[5]) ? node28739 : node28732;
														assign node28732 = (inp[9]) ? node28736 : node28733;
															assign node28733 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node28736 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node28739 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node28742 = (inp[9]) ? node28750 : node28743;
														assign node28743 = (inp[10]) ? node28747 : node28744;
															assign node28744 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node28747 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node28750 = (inp[10]) ? 4'b0000 : node28751;
															assign node28751 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node28755 = (inp[13]) ? node28815 : node28756;
											assign node28756 = (inp[2]) ? node28786 : node28757;
												assign node28757 = (inp[5]) ? node28775 : node28758;
													assign node28758 = (inp[1]) ? node28772 : node28759;
														assign node28759 = (inp[11]) ? node28765 : node28760;
															assign node28760 = (inp[10]) ? 4'b0101 : node28761;
																assign node28761 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node28765 = (inp[9]) ? node28769 : node28766;
																assign node28766 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node28769 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node28772 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node28775 = (inp[1]) ? node28781 : node28776;
														assign node28776 = (inp[9]) ? node28778 : 4'b0000;
															assign node28778 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node28781 = (inp[9]) ? 4'b0001 : node28782;
															assign node28782 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node28786 = (inp[1]) ? node28802 : node28787;
													assign node28787 = (inp[5]) ? node28795 : node28788;
														assign node28788 = (inp[9]) ? node28792 : node28789;
															assign node28789 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node28792 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node28795 = (inp[10]) ? node28797 : 4'b0100;
															assign node28797 = (inp[9]) ? node28799 : 4'b0101;
																assign node28799 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node28802 = (inp[11]) ? node28810 : node28803;
														assign node28803 = (inp[10]) ? node28807 : node28804;
															assign node28804 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node28807 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node28810 = (inp[9]) ? 4'b0101 : node28811;
															assign node28811 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node28815 = (inp[2]) ? node28831 : node28816;
												assign node28816 = (inp[1]) ? node28824 : node28817;
													assign node28817 = (inp[5]) ? 4'b0101 : node28818;
														assign node28818 = (inp[9]) ? node28820 : 4'b0000;
															assign node28820 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node28824 = (inp[9]) ? node28828 : node28825;
														assign node28825 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node28828 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node28831 = (inp[1]) ? node28841 : node28832;
													assign node28832 = (inp[5]) ? 4'b0001 : node28833;
														assign node28833 = (inp[9]) ? 4'b0101 : node28834;
															assign node28834 = (inp[11]) ? node28836 : 4'b0101;
																assign node28836 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node28841 = (inp[10]) ? 4'b0001 : node28842;
														assign node28842 = (inp[9]) ? 4'b0001 : 4'b0000;
								assign node28846 = (inp[5]) ? node29078 : node28847;
									assign node28847 = (inp[0]) ? node28967 : node28848;
										assign node28848 = (inp[10]) ? node28906 : node28849;
											assign node28849 = (inp[9]) ? node28877 : node28850;
												assign node28850 = (inp[4]) ? node28868 : node28851;
													assign node28851 = (inp[13]) ? node28859 : node28852;
														assign node28852 = (inp[11]) ? node28856 : node28853;
															assign node28853 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node28856 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node28859 = (inp[2]) ? node28865 : node28860;
															assign node28860 = (inp[1]) ? 4'b0100 : node28861;
																assign node28861 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node28865 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node28868 = (inp[13]) ? 4'b0001 : node28869;
														assign node28869 = (inp[1]) ? node28873 : node28870;
															assign node28870 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node28873 = (inp[11]) ? 4'b0100 : 4'b0001;
												assign node28877 = (inp[11]) ? node28889 : node28878;
													assign node28878 = (inp[13]) ? node28880 : 4'b0100;
														assign node28880 = (inp[2]) ? node28886 : node28881;
															assign node28881 = (inp[1]) ? node28883 : 4'b0000;
																assign node28883 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node28886 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node28889 = (inp[1]) ? node28895 : node28890;
														assign node28890 = (inp[2]) ? node28892 : 4'b0000;
															assign node28892 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node28895 = (inp[2]) ? node28899 : node28896;
															assign node28896 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node28899 = (inp[13]) ? node28903 : node28900;
																assign node28900 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node28903 = (inp[4]) ? 4'b0001 : 4'b0000;
											assign node28906 = (inp[9]) ? node28936 : node28907;
												assign node28907 = (inp[11]) ? node28927 : node28908;
													assign node28908 = (inp[4]) ? node28920 : node28909;
														assign node28909 = (inp[2]) ? node28913 : node28910;
															assign node28910 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node28913 = (inp[13]) ? node28917 : node28914;
																assign node28914 = (inp[1]) ? 4'b0100 : 4'b0001;
																assign node28917 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node28920 = (inp[13]) ? node28922 : 4'b0000;
															assign node28922 = (inp[2]) ? 4'b0100 : node28923;
																assign node28923 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node28927 = (inp[4]) ? node28931 : node28928;
														assign node28928 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node28931 = (inp[2]) ? 4'b0101 : node28932;
															assign node28932 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node28936 = (inp[11]) ? node28946 : node28937;
													assign node28937 = (inp[2]) ? node28943 : node28938;
														assign node28938 = (inp[4]) ? 4'b0101 : node28939;
															assign node28939 = (inp[1]) ? 4'b0100 : 4'b0001;
														assign node28943 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node28946 = (inp[4]) ? node28958 : node28947;
														assign node28947 = (inp[2]) ? node28953 : node28948;
															assign node28948 = (inp[13]) ? 4'b0100 : node28949;
																assign node28949 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node28953 = (inp[13]) ? 4'b0001 : node28954;
																assign node28954 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node28958 = (inp[13]) ? node28962 : node28959;
															assign node28959 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node28962 = (inp[1]) ? node28964 : 4'b0100;
																assign node28964 = (inp[2]) ? 4'b0000 : 4'b0100;
										assign node28967 = (inp[13]) ? node29013 : node28968;
											assign node28968 = (inp[2]) ? node28996 : node28969;
												assign node28969 = (inp[1]) ? node28989 : node28970;
													assign node28970 = (inp[4]) ? node28980 : node28971;
														assign node28971 = (inp[11]) ? node28973 : 4'b0101;
															assign node28973 = (inp[10]) ? node28977 : node28974;
																assign node28974 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node28977 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node28980 = (inp[9]) ? 4'b0100 : node28981;
															assign node28981 = (inp[10]) ? node28985 : node28982;
																assign node28982 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node28985 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node28989 = (inp[10]) ? node28993 : node28990;
														assign node28990 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node28993 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node28996 = (inp[1]) ? node29006 : node28997;
													assign node28997 = (inp[9]) ? 4'b0001 : node28998;
														assign node28998 = (inp[10]) ? node29000 : 4'b0001;
															assign node29000 = (inp[11]) ? node29002 : 4'b0000;
																assign node29002 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node29006 = (inp[11]) ? node29008 : 4'b0101;
														assign node29008 = (inp[10]) ? node29010 : 4'b0101;
															assign node29010 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node29013 = (inp[10]) ? node29051 : node29014;
												assign node29014 = (inp[9]) ? node29034 : node29015;
													assign node29015 = (inp[4]) ? node29025 : node29016;
														assign node29016 = (inp[1]) ? node29022 : node29017;
															assign node29017 = (inp[11]) ? node29019 : 4'b0101;
																assign node29019 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node29022 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node29025 = (inp[2]) ? node29031 : node29026;
															assign node29026 = (inp[1]) ? 4'b0100 : node29027;
																assign node29027 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node29031 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node29034 = (inp[1]) ? node29044 : node29035;
														assign node29035 = (inp[2]) ? node29039 : node29036;
															assign node29036 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node29039 = (inp[4]) ? 4'b0101 : node29040;
																assign node29040 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node29044 = (inp[2]) ? 4'b0001 : node29045;
															assign node29045 = (inp[4]) ? 4'b0101 : node29046;
																assign node29046 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node29051 = (inp[9]) ? node29063 : node29052;
													assign node29052 = (inp[4]) ? node29058 : node29053;
														assign node29053 = (inp[2]) ? node29055 : 4'b0001;
															assign node29055 = (inp[11]) ? 4'b0001 : 4'b0100;
														assign node29058 = (inp[2]) ? node29060 : 4'b0101;
															assign node29060 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node29063 = (inp[4]) ? node29071 : node29064;
														assign node29064 = (inp[2]) ? node29068 : node29065;
															assign node29065 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node29068 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node29071 = (inp[1]) ? 4'b0100 : node29072;
															assign node29072 = (inp[2]) ? 4'b0100 : node29073;
																assign node29073 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node29078 = (inp[11]) ? node29168 : node29079;
										assign node29079 = (inp[4]) ? node29127 : node29080;
											assign node29080 = (inp[0]) ? node29104 : node29081;
												assign node29081 = (inp[9]) ? node29095 : node29082;
													assign node29082 = (inp[10]) ? node29090 : node29083;
														assign node29083 = (inp[2]) ? node29087 : node29084;
															assign node29084 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node29087 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node29090 = (inp[2]) ? 4'b0000 : node29091;
															assign node29091 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node29095 = (inp[2]) ? node29099 : node29096;
														assign node29096 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node29099 = (inp[13]) ? 4'b0001 : node29100;
															assign node29100 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node29104 = (inp[2]) ? node29116 : node29105;
													assign node29105 = (inp[13]) ? node29111 : node29106;
														assign node29106 = (inp[1]) ? node29108 : 4'b0001;
															assign node29108 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node29111 = (inp[10]) ? node29113 : 4'b0101;
															assign node29113 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node29116 = (inp[13]) ? node29122 : node29117;
														assign node29117 = (inp[9]) ? 4'b0100 : node29118;
															assign node29118 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node29122 = (inp[10]) ? node29124 : 4'b0000;
															assign node29124 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node29127 = (inp[13]) ? node29139 : node29128;
												assign node29128 = (inp[2]) ? node29136 : node29129;
													assign node29129 = (inp[10]) ? node29133 : node29130;
														assign node29130 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node29133 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node29136 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node29139 = (inp[2]) ? node29153 : node29140;
													assign node29140 = (inp[0]) ? node29148 : node29141;
														assign node29141 = (inp[1]) ? node29143 : 4'b0100;
															assign node29143 = (inp[10]) ? node29145 : 4'b0101;
																assign node29145 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29148 = (inp[9]) ? node29150 : 4'b0100;
															assign node29150 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node29153 = (inp[9]) ? node29161 : node29154;
														assign node29154 = (inp[10]) ? node29158 : node29155;
															assign node29155 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node29158 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node29161 = (inp[0]) ? node29165 : node29162;
															assign node29162 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node29165 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node29168 = (inp[4]) ? node29212 : node29169;
											assign node29169 = (inp[2]) ? node29191 : node29170;
												assign node29170 = (inp[13]) ? node29184 : node29171;
													assign node29171 = (inp[0]) ? node29177 : node29172;
														assign node29172 = (inp[10]) ? node29174 : 4'b0000;
															assign node29174 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node29177 = (inp[10]) ? node29181 : node29178;
															assign node29178 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node29181 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node29184 = (inp[0]) ? 4'b0100 : node29185;
														assign node29185 = (inp[1]) ? node29187 : 4'b0101;
															assign node29187 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node29191 = (inp[13]) ? node29199 : node29192;
													assign node29192 = (inp[1]) ? node29194 : 4'b0100;
														assign node29194 = (inp[9]) ? node29196 : 4'b0101;
															assign node29196 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node29199 = (inp[1]) ? node29205 : node29200;
														assign node29200 = (inp[0]) ? 4'b0001 : node29201;
															assign node29201 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node29205 = (inp[9]) ? node29209 : node29206;
															assign node29206 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node29209 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node29212 = (inp[13]) ? node29230 : node29213;
												assign node29213 = (inp[2]) ? node29223 : node29214;
													assign node29214 = (inp[0]) ? node29216 : 4'b0001;
														assign node29216 = (inp[10]) ? node29220 : node29217;
															assign node29217 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node29220 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node29223 = (inp[10]) ? node29227 : node29224;
														assign node29224 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29227 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node29230 = (inp[2]) ? node29242 : node29231;
													assign node29231 = (inp[1]) ? node29237 : node29232;
														assign node29232 = (inp[9]) ? 4'b0101 : node29233;
															assign node29233 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node29237 = (inp[0]) ? 4'b0100 : node29238;
															assign node29238 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node29242 = (inp[1]) ? node29250 : node29243;
														assign node29243 = (inp[0]) ? 4'b0000 : node29244;
															assign node29244 = (inp[9]) ? 4'b0000 : node29245;
																assign node29245 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node29250 = (inp[0]) ? node29252 : 4'b0001;
															assign node29252 = (inp[9]) ? 4'b0001 : node29253;
																assign node29253 = (inp[10]) ? 4'b0001 : 4'b0000;
						assign node29257 = (inp[13]) ? node29715 : node29258;
							assign node29258 = (inp[4]) ? node29524 : node29259;
								assign node29259 = (inp[12]) ? node29381 : node29260;
									assign node29260 = (inp[1]) ? node29310 : node29261;
										assign node29261 = (inp[15]) ? node29293 : node29262;
											assign node29262 = (inp[0]) ? node29286 : node29263;
												assign node29263 = (inp[11]) ? node29275 : node29264;
													assign node29264 = (inp[5]) ? node29270 : node29265;
														assign node29265 = (inp[9]) ? node29267 : 4'b0100;
															assign node29267 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node29270 = (inp[9]) ? node29272 : 4'b0101;
															assign node29272 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node29275 = (inp[5]) ? node29279 : node29276;
														assign node29276 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node29279 = (inp[2]) ? node29283 : node29280;
															assign node29280 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node29283 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node29286 = (inp[2]) ? node29290 : node29287;
													assign node29287 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node29290 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node29293 = (inp[5]) ? node29301 : node29294;
												assign node29294 = (inp[2]) ? node29298 : node29295;
													assign node29295 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node29298 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node29301 = (inp[9]) ? node29303 : 4'b0001;
													assign node29303 = (inp[2]) ? node29307 : node29304;
														assign node29304 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node29307 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node29310 = (inp[15]) ? node29358 : node29311;
											assign node29311 = (inp[10]) ? node29331 : node29312;
												assign node29312 = (inp[2]) ? node29324 : node29313;
													assign node29313 = (inp[9]) ? node29319 : node29314;
														assign node29314 = (inp[0]) ? node29316 : 4'b0000;
															assign node29316 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node29319 = (inp[0]) ? node29321 : 4'b0001;
															assign node29321 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node29324 = (inp[9]) ? 4'b0000 : node29325;
														assign node29325 = (inp[5]) ? node29327 : 4'b0001;
															assign node29327 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node29331 = (inp[5]) ? node29341 : node29332;
													assign node29332 = (inp[11]) ? node29334 : 4'b0000;
														assign node29334 = (inp[0]) ? node29336 : 4'b0000;
															assign node29336 = (inp[9]) ? 4'b0001 : node29337;
																assign node29337 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node29341 = (inp[0]) ? node29351 : node29342;
														assign node29342 = (inp[11]) ? node29344 : 4'b0001;
															assign node29344 = (inp[9]) ? node29348 : node29345;
																assign node29345 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node29348 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node29351 = (inp[2]) ? node29355 : node29352;
															assign node29352 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node29355 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node29358 = (inp[9]) ? node29370 : node29359;
												assign node29359 = (inp[2]) ? node29365 : node29360;
													assign node29360 = (inp[0]) ? node29362 : 4'b0001;
														assign node29362 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node29365 = (inp[5]) ? node29367 : 4'b0000;
														assign node29367 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node29370 = (inp[2]) ? node29376 : node29371;
													assign node29371 = (inp[0]) ? node29373 : 4'b0000;
														assign node29373 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node29376 = (inp[0]) ? node29378 : 4'b0001;
														assign node29378 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node29381 = (inp[1]) ? node29435 : node29382;
										assign node29382 = (inp[15]) ? node29412 : node29383;
											assign node29383 = (inp[10]) ? node29393 : node29384;
												assign node29384 = (inp[5]) ? node29386 : 4'b0000;
													assign node29386 = (inp[9]) ? node29390 : node29387;
														assign node29387 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node29390 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node29393 = (inp[2]) ? node29399 : node29394;
													assign node29394 = (inp[9]) ? 4'b0001 : node29395;
														assign node29395 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node29399 = (inp[9]) ? node29405 : node29400;
														assign node29400 = (inp[0]) ? 4'b0001 : node29401;
															assign node29401 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node29405 = (inp[11]) ? 4'b0000 : node29406;
															assign node29406 = (inp[0]) ? 4'b0000 : node29407;
																assign node29407 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node29412 = (inp[9]) ? node29424 : node29413;
												assign node29413 = (inp[0]) ? node29421 : node29414;
													assign node29414 = (inp[2]) ? node29418 : node29415;
														assign node29415 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node29418 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node29421 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node29424 = (inp[11]) ? 4'b0100 : node29425;
													assign node29425 = (inp[2]) ? node29429 : node29426;
														assign node29426 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node29429 = (inp[5]) ? 4'b0100 : node29430;
															assign node29430 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node29435 = (inp[0]) ? node29481 : node29436;
											assign node29436 = (inp[9]) ? node29452 : node29437;
												assign node29437 = (inp[11]) ? node29439 : 4'b0101;
													assign node29439 = (inp[10]) ? node29447 : node29440;
														assign node29440 = (inp[15]) ? node29442 : 4'b0101;
															assign node29442 = (inp[2]) ? 4'b0101 : node29443;
																assign node29443 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node29447 = (inp[15]) ? 4'b0100 : node29448;
															assign node29448 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node29452 = (inp[10]) ? node29466 : node29453;
													assign node29453 = (inp[15]) ? node29455 : 4'b0101;
														assign node29455 = (inp[11]) ? node29461 : node29456;
															assign node29456 = (inp[2]) ? 4'b0101 : node29457;
																assign node29457 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node29461 = (inp[2]) ? 4'b0100 : node29462;
																assign node29462 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node29466 = (inp[5]) ? node29476 : node29467;
														assign node29467 = (inp[11]) ? 4'b0101 : node29468;
															assign node29468 = (inp[2]) ? node29472 : node29469;
																assign node29469 = (inp[15]) ? 4'b0100 : 4'b0101;
																assign node29472 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node29476 = (inp[15]) ? node29478 : 4'b0100;
															assign node29478 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node29481 = (inp[10]) ? node29503 : node29482;
												assign node29482 = (inp[2]) ? node29496 : node29483;
													assign node29483 = (inp[5]) ? node29491 : node29484;
														assign node29484 = (inp[9]) ? node29488 : node29485;
															assign node29485 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node29488 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node29491 = (inp[15]) ? 4'b0100 : node29492;
															assign node29492 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node29496 = (inp[15]) ? node29500 : node29497;
														assign node29497 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29500 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node29503 = (inp[9]) ? node29515 : node29504;
													assign node29504 = (inp[11]) ? node29512 : node29505;
														assign node29505 = (inp[5]) ? node29507 : 4'b0100;
															assign node29507 = (inp[2]) ? node29509 : 4'b0101;
																assign node29509 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node29512 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node29515 = (inp[5]) ? node29519 : node29516;
														assign node29516 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node29519 = (inp[11]) ? node29521 : 4'b0100;
															assign node29521 = (inp[15]) ? 4'b0101 : 4'b0100;
								assign node29524 = (inp[0]) ? node29592 : node29525;
									assign node29525 = (inp[10]) ? node29569 : node29526;
										assign node29526 = (inp[5]) ? node29546 : node29527;
											assign node29527 = (inp[9]) ? node29539 : node29528;
												assign node29528 = (inp[15]) ? node29534 : node29529;
													assign node29529 = (inp[1]) ? 4'b0100 : node29530;
														assign node29530 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node29534 = (inp[1]) ? 4'b0101 : node29535;
														assign node29535 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node29539 = (inp[15]) ? node29541 : 4'b0101;
													assign node29541 = (inp[1]) ? 4'b0100 : node29542;
														assign node29542 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node29546 = (inp[9]) ? node29558 : node29547;
												assign node29547 = (inp[12]) ? node29553 : node29548;
													assign node29548 = (inp[1]) ? node29550 : 4'b0100;
														assign node29550 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node29553 = (inp[15]) ? 4'b0101 : node29554;
														assign node29554 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node29558 = (inp[12]) ? node29564 : node29559;
													assign node29559 = (inp[1]) ? node29561 : 4'b0101;
														assign node29561 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node29564 = (inp[1]) ? node29566 : 4'b0100;
														assign node29566 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node29569 = (inp[15]) ? node29581 : node29570;
											assign node29570 = (inp[9]) ? node29576 : node29571;
												assign node29571 = (inp[12]) ? node29573 : 4'b0100;
													assign node29573 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node29576 = (inp[12]) ? node29578 : 4'b0101;
													assign node29578 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node29581 = (inp[9]) ? node29587 : node29582;
												assign node29582 = (inp[12]) ? 4'b0101 : node29583;
													assign node29583 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node29587 = (inp[1]) ? 4'b0100 : node29588;
													assign node29588 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node29592 = (inp[1]) ? node29664 : node29593;
										assign node29593 = (inp[2]) ? node29621 : node29594;
											assign node29594 = (inp[12]) ? node29614 : node29595;
												assign node29595 = (inp[11]) ? node29609 : node29596;
													assign node29596 = (inp[10]) ? node29602 : node29597;
														assign node29597 = (inp[5]) ? node29599 : 4'b0100;
															assign node29599 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29602 = (inp[5]) ? 4'b0100 : node29603;
															assign node29603 = (inp[15]) ? 4'b0101 : node29604;
																assign node29604 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node29609 = (inp[9]) ? 4'b0100 : node29610;
														assign node29610 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node29614 = (inp[9]) ? node29618 : node29615;
													assign node29615 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node29618 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node29621 = (inp[11]) ? node29645 : node29622;
												assign node29622 = (inp[15]) ? node29640 : node29623;
													assign node29623 = (inp[10]) ? node29631 : node29624;
														assign node29624 = (inp[9]) ? node29628 : node29625;
															assign node29625 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node29628 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node29631 = (inp[5]) ? 4'b0100 : node29632;
															assign node29632 = (inp[12]) ? node29636 : node29633;
																assign node29633 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node29636 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node29640 = (inp[10]) ? node29642 : 4'b0100;
														assign node29642 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node29645 = (inp[12]) ? node29657 : node29646;
													assign node29646 = (inp[5]) ? node29650 : node29647;
														assign node29647 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node29650 = (inp[10]) ? node29652 : 4'b0101;
															assign node29652 = (inp[15]) ? node29654 : 4'b0100;
																assign node29654 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node29657 = (inp[15]) ? node29661 : node29658;
														assign node29658 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29661 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node29664 = (inp[2]) ? node29694 : node29665;
											assign node29665 = (inp[10]) ? node29687 : node29666;
												assign node29666 = (inp[12]) ? node29680 : node29667;
													assign node29667 = (inp[5]) ? 4'b0101 : node29668;
														assign node29668 = (inp[11]) ? node29674 : node29669;
															assign node29669 = (inp[15]) ? node29671 : 4'b0101;
																assign node29671 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node29674 = (inp[9]) ? node29676 : 4'b0100;
																assign node29676 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node29680 = (inp[9]) ? node29684 : node29681;
														assign node29681 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node29684 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node29687 = (inp[9]) ? node29691 : node29688;
													assign node29688 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node29691 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node29694 = (inp[10]) ? node29708 : node29695;
												assign node29695 = (inp[5]) ? node29701 : node29696;
													assign node29696 = (inp[9]) ? node29698 : 4'b0101;
														assign node29698 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node29701 = (inp[15]) ? node29705 : node29702;
														assign node29702 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29705 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node29708 = (inp[9]) ? node29712 : node29709;
													assign node29709 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node29712 = (inp[15]) ? 4'b0100 : 4'b0101;
							assign node29715 = (inp[4]) ? node30005 : node29716;
								assign node29716 = (inp[12]) ? node29880 : node29717;
									assign node29717 = (inp[15]) ? node29787 : node29718;
										assign node29718 = (inp[1]) ? node29752 : node29719;
											assign node29719 = (inp[11]) ? node29737 : node29720;
												assign node29720 = (inp[5]) ? node29732 : node29721;
													assign node29721 = (inp[0]) ? node29727 : node29722;
														assign node29722 = (inp[2]) ? node29724 : 4'b0001;
															assign node29724 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node29727 = (inp[9]) ? 4'b0000 : node29728;
															assign node29728 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node29732 = (inp[9]) ? 4'b0001 : node29733;
														assign node29733 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node29737 = (inp[2]) ? node29741 : node29738;
													assign node29738 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node29741 = (inp[9]) ? node29747 : node29742;
														assign node29742 = (inp[0]) ? 4'b0001 : node29743;
															assign node29743 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node29747 = (inp[0]) ? 4'b0000 : node29748;
															assign node29748 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node29752 = (inp[10]) ? node29772 : node29753;
												assign node29753 = (inp[9]) ? node29763 : node29754;
													assign node29754 = (inp[11]) ? node29756 : 4'b0100;
														assign node29756 = (inp[2]) ? node29760 : node29757;
															assign node29757 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node29760 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node29763 = (inp[2]) ? node29767 : node29764;
														assign node29764 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node29767 = (inp[0]) ? 4'b0100 : node29768;
															assign node29768 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node29772 = (inp[0]) ? node29780 : node29773;
													assign node29773 = (inp[2]) ? node29775 : 4'b0101;
														assign node29775 = (inp[9]) ? 4'b0101 : node29776;
															assign node29776 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node29780 = (inp[2]) ? node29784 : node29781;
														assign node29781 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29784 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node29787 = (inp[11]) ? node29839 : node29788;
											assign node29788 = (inp[0]) ? node29816 : node29789;
												assign node29789 = (inp[2]) ? node29797 : node29790;
													assign node29790 = (inp[9]) ? 4'b0101 : node29791;
														assign node29791 = (inp[1]) ? 4'b0100 : node29792;
															assign node29792 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node29797 = (inp[1]) ? node29807 : node29798;
														assign node29798 = (inp[10]) ? 4'b0100 : node29799;
															assign node29799 = (inp[5]) ? node29803 : node29800;
																assign node29800 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node29803 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node29807 = (inp[10]) ? 4'b0101 : node29808;
															assign node29808 = (inp[5]) ? node29812 : node29809;
																assign node29809 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node29812 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node29816 = (inp[10]) ? node29830 : node29817;
													assign node29817 = (inp[9]) ? node29825 : node29818;
														assign node29818 = (inp[1]) ? node29822 : node29819;
															assign node29819 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node29822 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node29825 = (inp[1]) ? node29827 : 4'b0100;
															assign node29827 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node29830 = (inp[9]) ? node29832 : 4'b0100;
														assign node29832 = (inp[1]) ? node29836 : node29833;
															assign node29833 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node29836 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node29839 = (inp[1]) ? node29863 : node29840;
												assign node29840 = (inp[10]) ? node29850 : node29841;
													assign node29841 = (inp[2]) ? node29845 : node29842;
														assign node29842 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node29845 = (inp[9]) ? node29847 : 4'b0100;
															assign node29847 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node29850 = (inp[0]) ? 4'b0101 : node29851;
														assign node29851 = (inp[2]) ? node29857 : node29852;
															assign node29852 = (inp[9]) ? 4'b0100 : node29853;
																assign node29853 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node29857 = (inp[5]) ? 4'b0101 : node29858;
																assign node29858 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node29863 = (inp[5]) ? node29875 : node29864;
													assign node29864 = (inp[9]) ? 4'b0101 : node29865;
														assign node29865 = (inp[10]) ? 4'b0101 : node29866;
															assign node29866 = (inp[2]) ? node29870 : node29867;
																assign node29867 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node29870 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node29875 = (inp[9]) ? node29877 : 4'b0101;
														assign node29877 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node29880 = (inp[1]) ? node29920 : node29881;
										assign node29881 = (inp[15]) ? node29897 : node29882;
											assign node29882 = (inp[9]) ? node29888 : node29883;
												assign node29883 = (inp[2]) ? node29885 : 4'b0101;
													assign node29885 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node29888 = (inp[2]) ? node29894 : node29889;
													assign node29889 = (inp[0]) ? node29891 : 4'b0100;
														assign node29891 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node29894 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node29897 = (inp[9]) ? node29909 : node29898;
												assign node29898 = (inp[2]) ? node29904 : node29899;
													assign node29899 = (inp[0]) ? 4'b0000 : node29900;
														assign node29900 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node29904 = (inp[5]) ? 4'b0001 : node29905;
														assign node29905 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node29909 = (inp[2]) ? node29915 : node29910;
													assign node29910 = (inp[5]) ? 4'b0001 : node29911;
														assign node29911 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node29915 = (inp[5]) ? 4'b0000 : node29916;
														assign node29916 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node29920 = (inp[10]) ? node29952 : node29921;
											assign node29921 = (inp[5]) ? node29935 : node29922;
												assign node29922 = (inp[11]) ? node29924 : 4'b0000;
													assign node29924 = (inp[9]) ? node29930 : node29925;
														assign node29925 = (inp[2]) ? node29927 : 4'b0000;
															assign node29927 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node29930 = (inp[2]) ? 4'b0001 : node29931;
															assign node29931 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node29935 = (inp[11]) ? node29945 : node29936;
													assign node29936 = (inp[15]) ? 4'b0001 : node29937;
														assign node29937 = (inp[9]) ? node29941 : node29938;
															assign node29938 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node29941 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node29945 = (inp[2]) ? node29949 : node29946;
														assign node29946 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node29949 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node29952 = (inp[11]) ? node29990 : node29953;
												assign node29953 = (inp[15]) ? node29975 : node29954;
													assign node29954 = (inp[0]) ? node29968 : node29955;
														assign node29955 = (inp[9]) ? node29963 : node29956;
															assign node29956 = (inp[5]) ? node29960 : node29957;
																assign node29957 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node29960 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node29963 = (inp[5]) ? node29965 : 4'b0000;
																assign node29965 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node29968 = (inp[2]) ? node29972 : node29969;
															assign node29969 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node29972 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node29975 = (inp[9]) ? node29981 : node29976;
														assign node29976 = (inp[5]) ? 4'b0000 : node29977;
															assign node29977 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node29981 = (inp[0]) ? node29987 : node29982;
															assign node29982 = (inp[2]) ? 4'b0001 : node29983;
																assign node29983 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node29987 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node29990 = (inp[15]) ? node29998 : node29991;
													assign node29991 = (inp[5]) ? 4'b0001 : node29992;
														assign node29992 = (inp[9]) ? node29994 : 4'b0001;
															assign node29994 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node29998 = (inp[0]) ? 4'b0001 : node29999;
														assign node29999 = (inp[9]) ? node30001 : 4'b0000;
															assign node30001 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node30005 = (inp[9]) ? node30019 : node30006;
									assign node30006 = (inp[1]) ? 4'b0001 : node30007;
										assign node30007 = (inp[12]) ? node30013 : node30008;
											assign node30008 = (inp[15]) ? 4'b0000 : node30009;
												assign node30009 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node30013 = (inp[0]) ? 4'b0001 : node30014;
												assign node30014 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node30019 = (inp[1]) ? 4'b0000 : node30020;
										assign node30020 = (inp[12]) ? node30026 : node30021;
											assign node30021 = (inp[0]) ? 4'b0001 : node30022;
												assign node30022 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node30026 = (inp[15]) ? 4'b0000 : node30027;
												assign node30027 = (inp[0]) ? 4'b0000 : 4'b0001;
			assign node30032 = (inp[6]) ? node33348 : node30033;
				assign node30033 = (inp[12]) ? node31529 : node30034;
					assign node30034 = (inp[14]) ? node30848 : node30035;
						assign node30035 = (inp[15]) ? node30571 : node30036;
							assign node30036 = (inp[7]) ? node30260 : node30037;
								assign node30037 = (inp[2]) ? node30159 : node30038;
									assign node30038 = (inp[4]) ? node30086 : node30039;
										assign node30039 = (inp[9]) ? node30063 : node30040;
											assign node30040 = (inp[10]) ? node30052 : node30041;
												assign node30041 = (inp[13]) ? node30047 : node30042;
													assign node30042 = (inp[1]) ? node30044 : 4'b0000;
														assign node30044 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node30047 = (inp[1]) ? node30049 : 4'b0001;
														assign node30049 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node30052 = (inp[13]) ? node30058 : node30053;
													assign node30053 = (inp[1]) ? node30055 : 4'b0001;
														assign node30055 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node30058 = (inp[11]) ? node30060 : 4'b0000;
														assign node30060 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node30063 = (inp[13]) ? node30075 : node30064;
												assign node30064 = (inp[10]) ? node30070 : node30065;
													assign node30065 = (inp[11]) ? node30067 : 4'b0000;
														assign node30067 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node30070 = (inp[11]) ? node30072 : 4'b0001;
														assign node30072 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node30075 = (inp[10]) ? node30081 : node30076;
													assign node30076 = (inp[1]) ? node30078 : 4'b0001;
														assign node30078 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node30081 = (inp[11]) ? node30083 : 4'b0000;
														assign node30083 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node30086 = (inp[5]) ? node30108 : node30087;
											assign node30087 = (inp[10]) ? node30099 : node30088;
												assign node30088 = (inp[13]) ? node30094 : node30089;
													assign node30089 = (inp[11]) ? node30091 : 4'b0000;
														assign node30091 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node30094 = (inp[11]) ? node30096 : 4'b0001;
														assign node30096 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node30099 = (inp[1]) ? node30101 : 4'b0000;
													assign node30101 = (inp[11]) ? node30105 : node30102;
														assign node30102 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node30105 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node30108 = (inp[0]) ? node30132 : node30109;
												assign node30109 = (inp[9]) ? node30115 : node30110;
													assign node30110 = (inp[11]) ? node30112 : 4'b0101;
														assign node30112 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node30115 = (inp[1]) ? node30127 : node30116;
														assign node30116 = (inp[10]) ? node30122 : node30117;
															assign node30117 = (inp[11]) ? 4'b0101 : node30118;
																assign node30118 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node30122 = (inp[11]) ? 4'b0100 : node30123;
																assign node30123 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node30127 = (inp[13]) ? node30129 : 4'b0101;
															assign node30129 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node30132 = (inp[11]) ? node30146 : node30133;
													assign node30133 = (inp[10]) ? node30141 : node30134;
														assign node30134 = (inp[9]) ? 4'b0101 : node30135;
															assign node30135 = (inp[1]) ? node30137 : 4'b0100;
																assign node30137 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node30141 = (inp[1]) ? node30143 : 4'b0101;
															assign node30143 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node30146 = (inp[9]) ? 4'b0100 : node30147;
														assign node30147 = (inp[1]) ? node30153 : node30148;
															assign node30148 = (inp[10]) ? node30150 : 4'b0100;
																assign node30150 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node30153 = (inp[10]) ? 4'b0100 : node30154;
																assign node30154 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node30159 = (inp[5]) ? node30219 : node30160;
										assign node30160 = (inp[4]) ? node30190 : node30161;
											assign node30161 = (inp[9]) ? node30175 : node30162;
												assign node30162 = (inp[1]) ? node30164 : 4'b0100;
													assign node30164 = (inp[13]) ? node30170 : node30165;
														assign node30165 = (inp[0]) ? 4'b0101 : node30166;
															assign node30166 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node30170 = (inp[11]) ? 4'b0100 : node30171;
															assign node30171 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node30175 = (inp[11]) ? node30181 : node30176;
													assign node30176 = (inp[10]) ? node30178 : 4'b0100;
														assign node30178 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node30181 = (inp[10]) ? node30183 : 4'b0101;
														assign node30183 = (inp[1]) ? node30187 : node30184;
															assign node30184 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node30187 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node30190 = (inp[1]) ? node30198 : node30191;
												assign node30191 = (inp[10]) ? node30195 : node30192;
													assign node30192 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node30195 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node30198 = (inp[13]) ? node30210 : node30199;
													assign node30199 = (inp[9]) ? node30201 : 4'b0101;
														assign node30201 = (inp[0]) ? node30203 : 4'b0101;
															assign node30203 = (inp[10]) ? node30207 : node30204;
																assign node30204 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node30207 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node30210 = (inp[0]) ? 4'b0101 : node30211;
														assign node30211 = (inp[10]) ? node30215 : node30212;
															assign node30212 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node30215 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node30219 = (inp[4]) ? node30239 : node30220;
											assign node30220 = (inp[10]) ? node30228 : node30221;
												assign node30221 = (inp[13]) ? node30225 : node30222;
													assign node30222 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node30225 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node30228 = (inp[13]) ? node30234 : node30229;
													assign node30229 = (inp[1]) ? node30231 : 4'b0101;
														assign node30231 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node30234 = (inp[1]) ? node30236 : 4'b0100;
														assign node30236 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node30239 = (inp[13]) ? node30251 : node30240;
												assign node30240 = (inp[10]) ? node30246 : node30241;
													assign node30241 = (inp[11]) ? node30243 : 4'b0000;
														assign node30243 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node30246 = (inp[11]) ? node30248 : 4'b0001;
														assign node30248 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node30251 = (inp[10]) ? node30257 : node30252;
													assign node30252 = (inp[1]) ? node30254 : 4'b0001;
														assign node30254 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node30257 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node30260 = (inp[2]) ? node30406 : node30261;
									assign node30261 = (inp[4]) ? node30333 : node30262;
										assign node30262 = (inp[11]) ? node30278 : node30263;
											assign node30263 = (inp[10]) ? node30271 : node30264;
												assign node30264 = (inp[5]) ? node30268 : node30265;
													assign node30265 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node30268 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node30271 = (inp[13]) ? node30275 : node30272;
													assign node30272 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node30275 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node30278 = (inp[9]) ? node30308 : node30279;
												assign node30279 = (inp[10]) ? node30295 : node30280;
													assign node30280 = (inp[0]) ? node30290 : node30281;
														assign node30281 = (inp[5]) ? 4'b0101 : node30282;
															assign node30282 = (inp[1]) ? node30286 : node30283;
																assign node30283 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node30286 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node30290 = (inp[13]) ? 4'b0101 : node30291;
															assign node30291 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node30295 = (inp[5]) ? node30301 : node30296;
														assign node30296 = (inp[0]) ? node30298 : 4'b0100;
															assign node30298 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node30301 = (inp[0]) ? node30303 : 4'b0101;
															assign node30303 = (inp[13]) ? 4'b0100 : node30304;
																assign node30304 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node30308 = (inp[5]) ? node30320 : node30309;
													assign node30309 = (inp[13]) ? node30313 : node30310;
														assign node30310 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node30313 = (inp[1]) ? node30317 : node30314;
															assign node30314 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node30317 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node30320 = (inp[13]) ? node30328 : node30321;
														assign node30321 = (inp[10]) ? node30325 : node30322;
															assign node30322 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node30325 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node30328 = (inp[1]) ? node30330 : 4'b0100;
															assign node30330 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node30333 = (inp[5]) ? node30373 : node30334;
											assign node30334 = (inp[9]) ? node30352 : node30335;
												assign node30335 = (inp[1]) ? node30343 : node30336;
													assign node30336 = (inp[10]) ? node30340 : node30337;
														assign node30337 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node30340 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node30343 = (inp[11]) ? node30345 : 4'b0100;
														assign node30345 = (inp[10]) ? node30349 : node30346;
															assign node30346 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node30349 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node30352 = (inp[0]) ? node30364 : node30353;
													assign node30353 = (inp[13]) ? 4'b0100 : node30354;
														assign node30354 = (inp[1]) ? node30356 : 4'b0100;
															assign node30356 = (inp[11]) ? node30360 : node30357;
																assign node30357 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node30360 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node30364 = (inp[13]) ? node30366 : 4'b0101;
														assign node30366 = (inp[1]) ? node30368 : 4'b0100;
															assign node30368 = (inp[11]) ? 4'b0101 : node30369;
																assign node30369 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node30373 = (inp[0]) ? node30391 : node30374;
												assign node30374 = (inp[9]) ? node30382 : node30375;
													assign node30375 = (inp[10]) ? node30379 : node30376;
														assign node30376 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node30379 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node30382 = (inp[11]) ? 4'b0001 : node30383;
														assign node30383 = (inp[13]) ? node30387 : node30384;
															assign node30384 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node30387 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node30391 = (inp[13]) ? node30395 : node30392;
													assign node30392 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node30395 = (inp[10]) ? node30401 : node30396;
														assign node30396 = (inp[1]) ? node30398 : 4'b0001;
															assign node30398 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node30401 = (inp[1]) ? node30403 : 4'b0000;
															assign node30403 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node30406 = (inp[5]) ? node30490 : node30407;
										assign node30407 = (inp[1]) ? node30453 : node30408;
											assign node30408 = (inp[0]) ? node30432 : node30409;
												assign node30409 = (inp[10]) ? node30425 : node30410;
													assign node30410 = (inp[13]) ? node30418 : node30411;
														assign node30411 = (inp[4]) ? node30415 : node30412;
															assign node30412 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node30415 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node30418 = (inp[4]) ? node30422 : node30419;
															assign node30419 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node30422 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node30425 = (inp[11]) ? node30427 : 4'b0001;
														assign node30427 = (inp[13]) ? 4'b0001 : node30428;
															assign node30428 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node30432 = (inp[10]) ? node30442 : node30433;
													assign node30433 = (inp[9]) ? 4'b0001 : node30434;
														assign node30434 = (inp[13]) ? node30436 : 4'b0001;
															assign node30436 = (inp[11]) ? node30438 : 4'b0000;
																assign node30438 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node30442 = (inp[13]) ? 4'b0000 : node30443;
														assign node30443 = (inp[9]) ? node30449 : node30444;
															assign node30444 = (inp[11]) ? node30446 : 4'b0000;
																assign node30446 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node30449 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node30453 = (inp[11]) ? node30467 : node30454;
												assign node30454 = (inp[13]) ? node30462 : node30455;
													assign node30455 = (inp[10]) ? node30459 : node30456;
														assign node30456 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node30459 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node30462 = (inp[10]) ? 4'b0000 : node30463;
														assign node30463 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node30467 = (inp[10]) ? node30475 : node30468;
													assign node30468 = (inp[4]) ? node30472 : node30469;
														assign node30469 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node30472 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node30475 = (inp[9]) ? node30481 : node30476;
														assign node30476 = (inp[13]) ? 4'b0001 : node30477;
															assign node30477 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node30481 = (inp[0]) ? node30483 : 4'b0000;
															assign node30483 = (inp[4]) ? node30487 : node30484;
																assign node30484 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node30487 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node30490 = (inp[4]) ? node30514 : node30491;
											assign node30491 = (inp[10]) ? node30503 : node30492;
												assign node30492 = (inp[13]) ? node30498 : node30493;
													assign node30493 = (inp[1]) ? 4'b0000 : node30494;
														assign node30494 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node30498 = (inp[11]) ? 4'b0001 : node30499;
														assign node30499 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node30503 = (inp[13]) ? node30509 : node30504;
													assign node30504 = (inp[11]) ? 4'b0001 : node30505;
														assign node30505 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node30509 = (inp[11]) ? 4'b0000 : node30510;
														assign node30510 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node30514 = (inp[9]) ? node30548 : node30515;
												assign node30515 = (inp[1]) ? node30533 : node30516;
													assign node30516 = (inp[11]) ? node30524 : node30517;
														assign node30517 = (inp[0]) ? node30519 : 4'b0100;
															assign node30519 = (inp[13]) ? node30521 : 4'b0101;
																assign node30521 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node30524 = (inp[0]) ? node30526 : 4'b0101;
															assign node30526 = (inp[10]) ? node30530 : node30527;
																assign node30527 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node30530 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node30533 = (inp[13]) ? node30541 : node30534;
														assign node30534 = (inp[11]) ? node30538 : node30535;
															assign node30535 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node30538 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node30541 = (inp[11]) ? node30545 : node30542;
															assign node30542 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node30545 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node30548 = (inp[0]) ? 4'b0100 : node30549;
													assign node30549 = (inp[1]) ? node30559 : node30550;
														assign node30550 = (inp[11]) ? node30554 : node30551;
															assign node30551 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node30554 = (inp[13]) ? 4'b0100 : node30555;
																assign node30555 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node30559 = (inp[13]) ? node30565 : node30560;
															assign node30560 = (inp[10]) ? node30562 : 4'b0101;
																assign node30562 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node30565 = (inp[11]) ? 4'b0100 : node30566;
																assign node30566 = (inp[10]) ? 4'b0101 : 4'b0100;
							assign node30571 = (inp[10]) ? node30711 : node30572;
								assign node30572 = (inp[1]) ? node30644 : node30573;
									assign node30573 = (inp[7]) ? node30589 : node30574;
										assign node30574 = (inp[4]) ? node30578 : node30575;
											assign node30575 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node30578 = (inp[2]) ? node30584 : node30579;
												assign node30579 = (inp[11]) ? node30581 : 4'b0110;
													assign node30581 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node30584 = (inp[5]) ? 4'b0010 : node30585;
													assign node30585 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node30589 = (inp[4]) ? node30633 : node30590;
											assign node30590 = (inp[2]) ? node30612 : node30591;
												assign node30591 = (inp[13]) ? node30605 : node30592;
													assign node30592 = (inp[9]) ? node30598 : node30593;
														assign node30593 = (inp[11]) ? 4'b0010 : node30594;
															assign node30594 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node30598 = (inp[11]) ? node30602 : node30599;
															assign node30599 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node30602 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node30605 = (inp[11]) ? node30609 : node30606;
														assign node30606 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node30609 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node30612 = (inp[0]) ? node30620 : node30613;
													assign node30613 = (inp[11]) ? node30617 : node30614;
														assign node30614 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node30617 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node30620 = (inp[9]) ? node30628 : node30621;
														assign node30621 = (inp[13]) ? node30623 : 4'b0111;
															assign node30623 = (inp[11]) ? 4'b0110 : node30624;
																assign node30624 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node30628 = (inp[5]) ? 4'b0110 : node30629;
															assign node30629 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node30633 = (inp[2]) ? node30639 : node30634;
												assign node30634 = (inp[11]) ? node30636 : 4'b0110;
													assign node30636 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node30639 = (inp[11]) ? 4'b0010 : node30640;
													assign node30640 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node30644 = (inp[7]) ? node30660 : node30645;
										assign node30645 = (inp[4]) ? node30649 : node30646;
											assign node30646 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node30649 = (inp[2]) ? node30655 : node30650;
												assign node30650 = (inp[11]) ? node30652 : 4'b0111;
													assign node30652 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node30655 = (inp[5]) ? 4'b0011 : node30656;
													assign node30656 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node30660 = (inp[4]) ? node30700 : node30661;
											assign node30661 = (inp[2]) ? node30679 : node30662;
												assign node30662 = (inp[0]) ? node30672 : node30663;
													assign node30663 = (inp[9]) ? 4'b0010 : node30664;
														assign node30664 = (inp[11]) ? node30668 : node30665;
															assign node30665 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node30668 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node30672 = (inp[5]) ? node30676 : node30673;
														assign node30673 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node30676 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node30679 = (inp[9]) ? node30691 : node30680;
													assign node30680 = (inp[13]) ? 4'b0110 : node30681;
														assign node30681 = (inp[0]) ? 4'b0111 : node30682;
															assign node30682 = (inp[5]) ? node30686 : node30683;
																assign node30683 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node30686 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node30691 = (inp[13]) ? node30693 : 4'b0111;
														assign node30693 = (inp[11]) ? node30697 : node30694;
															assign node30694 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node30697 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node30700 = (inp[2]) ? node30706 : node30701;
												assign node30701 = (inp[5]) ? 4'b0111 : node30702;
													assign node30702 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node30706 = (inp[11]) ? 4'b0011 : node30707;
													assign node30707 = (inp[5]) ? 4'b0010 : 4'b0011;
								assign node30711 = (inp[1]) ? node30773 : node30712;
									assign node30712 = (inp[7]) ? node30728 : node30713;
										assign node30713 = (inp[4]) ? node30717 : node30714;
											assign node30714 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node30717 = (inp[2]) ? node30723 : node30718;
												assign node30718 = (inp[5]) ? node30720 : 4'b0111;
													assign node30720 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node30723 = (inp[5]) ? 4'b0011 : node30724;
													assign node30724 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node30728 = (inp[4]) ? node30762 : node30729;
											assign node30729 = (inp[2]) ? node30737 : node30730;
												assign node30730 = (inp[11]) ? node30734 : node30731;
													assign node30731 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node30734 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node30737 = (inp[0]) ? node30745 : node30738;
													assign node30738 = (inp[5]) ? node30742 : node30739;
														assign node30739 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node30742 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node30745 = (inp[13]) ? node30753 : node30746;
														assign node30746 = (inp[9]) ? node30748 : 4'b0111;
															assign node30748 = (inp[5]) ? 4'b0110 : node30749;
																assign node30749 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node30753 = (inp[9]) ? 4'b0111 : node30754;
															assign node30754 = (inp[11]) ? node30758 : node30755;
																assign node30755 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node30758 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node30762 = (inp[2]) ? node30768 : node30763;
												assign node30763 = (inp[5]) ? 4'b0111 : node30764;
													assign node30764 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node30768 = (inp[11]) ? 4'b0011 : node30769;
													assign node30769 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node30773 = (inp[7]) ? node30789 : node30774;
										assign node30774 = (inp[4]) ? node30778 : node30775;
											assign node30775 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node30778 = (inp[2]) ? node30784 : node30779;
												assign node30779 = (inp[11]) ? node30781 : 4'b0110;
													assign node30781 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node30784 = (inp[11]) ? 4'b0010 : node30785;
													assign node30785 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node30789 = (inp[13]) ? node30813 : node30790;
											assign node30790 = (inp[5]) ? node30804 : node30791;
												assign node30791 = (inp[11]) ? node30799 : node30792;
													assign node30792 = (inp[4]) ? node30796 : node30793;
														assign node30793 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node30796 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node30799 = (inp[2]) ? 4'b0010 : node30800;
														assign node30800 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node30804 = (inp[11]) ? node30810 : node30805;
													assign node30805 = (inp[0]) ? 4'b0011 : node30806;
														assign node30806 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node30810 = (inp[0]) ? 4'b0110 : 4'b0010;
											assign node30813 = (inp[4]) ? node30837 : node30814;
												assign node30814 = (inp[2]) ? node30822 : node30815;
													assign node30815 = (inp[9]) ? 4'b0011 : node30816;
														assign node30816 = (inp[11]) ? 4'b0010 : node30817;
															assign node30817 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node30822 = (inp[9]) ? node30832 : node30823;
														assign node30823 = (inp[0]) ? node30827 : node30824;
															assign node30824 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node30827 = (inp[11]) ? node30829 : 4'b0111;
																assign node30829 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node30832 = (inp[11]) ? node30834 : 4'b0110;
															assign node30834 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node30837 = (inp[2]) ? node30843 : node30838;
													assign node30838 = (inp[11]) ? node30840 : 4'b0110;
														assign node30840 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node30843 = (inp[11]) ? 4'b0010 : node30844;
														assign node30844 = (inp[5]) ? 4'b0011 : 4'b0010;
						assign node30848 = (inp[1]) ? node31274 : node30849;
							assign node30849 = (inp[10]) ? node31065 : node30850;
								assign node30850 = (inp[15]) ? node30978 : node30851;
									assign node30851 = (inp[7]) ? node30907 : node30852;
										assign node30852 = (inp[2]) ? node30888 : node30853;
											assign node30853 = (inp[5]) ? node30871 : node30854;
												assign node30854 = (inp[9]) ? node30864 : node30855;
													assign node30855 = (inp[0]) ? node30861 : node30856;
														assign node30856 = (inp[13]) ? node30858 : 4'b0010;
															assign node30858 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node30861 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node30864 = (inp[13]) ? node30868 : node30865;
														assign node30865 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node30868 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node30871 = (inp[4]) ? node30881 : node30872;
													assign node30872 = (inp[9]) ? node30874 : 4'b0111;
														assign node30874 = (inp[0]) ? node30878 : node30875;
															assign node30875 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node30878 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node30881 = (inp[11]) ? node30885 : node30882;
														assign node30882 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node30885 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node30888 = (inp[5]) ? node30896 : node30889;
												assign node30889 = (inp[13]) ? node30893 : node30890;
													assign node30890 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node30893 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node30896 = (inp[4]) ? node30904 : node30897;
													assign node30897 = (inp[9]) ? node30899 : 4'b0010;
														assign node30899 = (inp[11]) ? 4'b0011 : node30900;
															assign node30900 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node30904 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node30907 = (inp[2]) ? node30943 : node30908;
											assign node30908 = (inp[4]) ? node30920 : node30909;
												assign node30909 = (inp[5]) ? node30917 : node30910;
													assign node30910 = (inp[11]) ? node30914 : node30911;
														assign node30911 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node30914 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node30917 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node30920 = (inp[9]) ? node30928 : node30921;
													assign node30921 = (inp[11]) ? node30925 : node30922;
														assign node30922 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node30925 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node30928 = (inp[5]) ? node30936 : node30929;
														assign node30929 = (inp[0]) ? 4'b0110 : node30930;
															assign node30930 = (inp[13]) ? node30932 : 4'b0110;
																assign node30932 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node30936 = (inp[11]) ? node30940 : node30937;
															assign node30937 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node30940 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node30943 = (inp[5]) ? node30961 : node30944;
												assign node30944 = (inp[13]) ? node30952 : node30945;
													assign node30945 = (inp[4]) ? node30949 : node30946;
														assign node30946 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node30949 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node30952 = (inp[0]) ? 4'b0010 : node30953;
														assign node30953 = (inp[4]) ? node30957 : node30954;
															assign node30954 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node30957 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node30961 = (inp[4]) ? node30969 : node30962;
													assign node30962 = (inp[11]) ? node30966 : node30963;
														assign node30963 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node30966 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node30969 = (inp[9]) ? node30971 : 4'b0011;
														assign node30971 = (inp[0]) ? node30975 : node30972;
															assign node30972 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node30975 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node30978 = (inp[7]) ? node31050 : node30979;
										assign node30979 = (inp[13]) ? node31017 : node30980;
											assign node30980 = (inp[11]) ? node31004 : node30981;
												assign node30981 = (inp[5]) ? node30995 : node30982;
													assign node30982 = (inp[0]) ? node30990 : node30983;
														assign node30983 = (inp[9]) ? 4'b0010 : node30984;
															assign node30984 = (inp[4]) ? node30986 : 4'b0110;
																assign node30986 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node30990 = (inp[9]) ? 4'b0110 : node30991;
															assign node30991 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node30995 = (inp[9]) ? node31001 : node30996;
														assign node30996 = (inp[2]) ? 4'b0111 : node30997;
															assign node30997 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node31001 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node31004 = (inp[5]) ? node31010 : node31005;
													assign node31005 = (inp[2]) ? 4'b0110 : node31006;
														assign node31006 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node31010 = (inp[0]) ? node31012 : 4'b0110;
														assign node31012 = (inp[2]) ? node31014 : 4'b0110;
															assign node31014 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node31017 = (inp[9]) ? node31031 : node31018;
												assign node31018 = (inp[2]) ? node31026 : node31019;
													assign node31019 = (inp[4]) ? 4'b0110 : node31020;
														assign node31020 = (inp[5]) ? 4'b0010 : node31021;
															assign node31021 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node31026 = (inp[4]) ? 4'b0010 : node31027;
														assign node31027 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node31031 = (inp[4]) ? node31039 : node31032;
													assign node31032 = (inp[2]) ? node31034 : 4'b0010;
														assign node31034 = (inp[5]) ? node31036 : 4'b0110;
															assign node31036 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node31039 = (inp[2]) ? 4'b0011 : node31040;
														assign node31040 = (inp[0]) ? node31044 : node31041;
															assign node31041 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node31044 = (inp[5]) ? node31046 : 4'b0111;
																assign node31046 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node31050 = (inp[4]) ? node31062 : node31051;
											assign node31051 = (inp[2]) ? node31057 : node31052;
												assign node31052 = (inp[11]) ? node31054 : 4'b0010;
													assign node31054 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node31057 = (inp[5]) ? 4'b0110 : node31058;
													assign node31058 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node31062 = (inp[2]) ? 4'b0010 : 4'b0110;
								assign node31065 = (inp[15]) ? node31223 : node31066;
									assign node31066 = (inp[9]) ? node31146 : node31067;
										assign node31067 = (inp[13]) ? node31105 : node31068;
											assign node31068 = (inp[11]) ? node31090 : node31069;
												assign node31069 = (inp[5]) ? node31083 : node31070;
													assign node31070 = (inp[0]) ? node31078 : node31071;
														assign node31071 = (inp[7]) ? node31075 : node31072;
															assign node31072 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node31075 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node31078 = (inp[4]) ? node31080 : 4'b0111;
															assign node31080 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node31083 = (inp[4]) ? node31085 : 4'b0010;
														assign node31085 = (inp[7]) ? node31087 : 4'b0010;
															assign node31087 = (inp[0]) ? 4'b0111 : 4'b0011;
												assign node31090 = (inp[2]) ? node31098 : node31091;
													assign node31091 = (inp[7]) ? 4'b0110 : node31092;
														assign node31092 = (inp[5]) ? node31094 : 4'b0010;
															assign node31094 = (inp[4]) ? 4'b0011 : 4'b0110;
													assign node31098 = (inp[4]) ? 4'b0010 : node31099;
														assign node31099 = (inp[5]) ? 4'b0110 : node31100;
															assign node31100 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node31105 = (inp[2]) ? node31129 : node31106;
												assign node31106 = (inp[11]) ? node31116 : node31107;
													assign node31107 = (inp[5]) ? node31109 : 4'b0010;
														assign node31109 = (inp[4]) ? node31113 : node31110;
															assign node31110 = (inp[7]) ? 4'b0011 : 4'b0110;
															assign node31113 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node31116 = (inp[4]) ? 4'b0111 : node31117;
														assign node31117 = (inp[0]) ? node31123 : node31118;
															assign node31118 = (inp[7]) ? 4'b0011 : node31119;
																assign node31119 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node31123 = (inp[5]) ? node31125 : 4'b0111;
																assign node31125 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node31129 = (inp[5]) ? node31139 : node31130;
													assign node31130 = (inp[7]) ? node31134 : node31131;
														assign node31131 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node31134 = (inp[4]) ? 4'b0011 : node31135;
															assign node31135 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node31139 = (inp[4]) ? 4'b0110 : node31140;
														assign node31140 = (inp[7]) ? 4'b0110 : node31141;
															assign node31141 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node31146 = (inp[11]) ? node31180 : node31147;
											assign node31147 = (inp[13]) ? node31163 : node31148;
												assign node31148 = (inp[2]) ? node31152 : node31149;
													assign node31149 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node31152 = (inp[7]) ? node31160 : node31153;
														assign node31153 = (inp[4]) ? node31157 : node31154;
															assign node31154 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node31157 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node31160 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node31163 = (inp[7]) ? node31173 : node31164;
													assign node31164 = (inp[2]) ? node31168 : node31165;
														assign node31165 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node31168 = (inp[4]) ? node31170 : 4'b0110;
															assign node31170 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node31173 = (inp[2]) ? 4'b0010 : node31174;
														assign node31174 = (inp[4]) ? 4'b0110 : node31175;
															assign node31175 = (inp[5]) ? 4'b0011 : 4'b0110;
											assign node31180 = (inp[2]) ? node31198 : node31181;
												assign node31181 = (inp[13]) ? node31193 : node31182;
													assign node31182 = (inp[7]) ? node31188 : node31183;
														assign node31183 = (inp[5]) ? node31185 : 4'b0010;
															assign node31185 = (inp[0]) ? 4'b0011 : 4'b0110;
														assign node31188 = (inp[4]) ? 4'b0110 : node31189;
															assign node31189 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node31193 = (inp[4]) ? node31195 : 4'b0011;
														assign node31195 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node31198 = (inp[7]) ? node31214 : node31199;
													assign node31199 = (inp[4]) ? node31207 : node31200;
														assign node31200 = (inp[13]) ? node31204 : node31201;
															assign node31201 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node31204 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node31207 = (inp[5]) ? node31211 : node31208;
															assign node31208 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node31211 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node31214 = (inp[13]) ? node31218 : node31215;
														assign node31215 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node31218 = (inp[5]) ? node31220 : 4'b0010;
															assign node31220 = (inp[0]) ? 4'b0011 : 4'b0111;
									assign node31223 = (inp[7]) ? node31259 : node31224;
										assign node31224 = (inp[4]) ? node31236 : node31225;
											assign node31225 = (inp[2]) ? node31231 : node31226;
												assign node31226 = (inp[5]) ? 4'b0011 : node31227;
													assign node31227 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node31231 = (inp[5]) ? node31233 : 4'b0111;
													assign node31233 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node31236 = (inp[2]) ? node31244 : node31237;
												assign node31237 = (inp[11]) ? node31241 : node31238;
													assign node31238 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node31241 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node31244 = (inp[0]) ? node31252 : node31245;
													assign node31245 = (inp[11]) ? node31249 : node31246;
														assign node31246 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node31249 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node31252 = (inp[5]) ? node31256 : node31253;
														assign node31253 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node31256 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node31259 = (inp[4]) ? node31271 : node31260;
											assign node31260 = (inp[2]) ? node31266 : node31261;
												assign node31261 = (inp[11]) ? node31263 : 4'b0011;
													assign node31263 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node31266 = (inp[5]) ? 4'b0111 : node31267;
													assign node31267 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node31271 = (inp[2]) ? 4'b0011 : 4'b0111;
							assign node31274 = (inp[10]) ? node31396 : node31275;
								assign node31275 = (inp[15]) ? node31347 : node31276;
									assign node31276 = (inp[13]) ? node31312 : node31277;
										assign node31277 = (inp[7]) ? node31297 : node31278;
											assign node31278 = (inp[2]) ? node31284 : node31279;
												assign node31279 = (inp[5]) ? node31281 : 4'b0010;
													assign node31281 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node31284 = (inp[4]) ? node31290 : node31285;
													assign node31285 = (inp[5]) ? 4'b0011 : node31286;
														assign node31286 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node31290 = (inp[11]) ? node31294 : node31291;
														assign node31291 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node31294 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node31297 = (inp[2]) ? node31305 : node31298;
												assign node31298 = (inp[4]) ? 4'b0110 : node31299;
													assign node31299 = (inp[5]) ? node31301 : 4'b0110;
														assign node31301 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node31305 = (inp[5]) ? node31309 : node31306;
													assign node31306 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node31309 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node31312 = (inp[2]) ? node31326 : node31313;
											assign node31313 = (inp[7]) ? node31319 : node31314;
												assign node31314 = (inp[5]) ? node31316 : 4'b0011;
													assign node31316 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node31319 = (inp[5]) ? node31321 : 4'b0111;
													assign node31321 = (inp[4]) ? 4'b0111 : node31322;
														assign node31322 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node31326 = (inp[7]) ? node31342 : node31327;
												assign node31327 = (inp[4]) ? node31333 : node31328;
													assign node31328 = (inp[5]) ? 4'b0010 : node31329;
														assign node31329 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node31333 = (inp[0]) ? node31335 : 4'b0111;
														assign node31335 = (inp[5]) ? node31339 : node31336;
															assign node31336 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node31339 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node31342 = (inp[4]) ? 4'b0011 : node31343;
													assign node31343 = (inp[5]) ? 4'b0111 : 4'b0010;
									assign node31347 = (inp[7]) ? node31381 : node31348;
										assign node31348 = (inp[4]) ? node31360 : node31349;
											assign node31349 = (inp[2]) ? node31355 : node31350;
												assign node31350 = (inp[5]) ? 4'b0011 : node31351;
													assign node31351 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node31355 = (inp[11]) ? 4'b0111 : node31356;
													assign node31356 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node31360 = (inp[2]) ? node31368 : node31361;
												assign node31361 = (inp[11]) ? node31365 : node31362;
													assign node31362 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node31365 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node31368 = (inp[9]) ? node31374 : node31369;
													assign node31369 = (inp[11]) ? 4'b0010 : node31370;
														assign node31370 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node31374 = (inp[11]) ? node31378 : node31375;
														assign node31375 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node31378 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node31381 = (inp[4]) ? node31393 : node31382;
											assign node31382 = (inp[2]) ? node31388 : node31383;
												assign node31383 = (inp[5]) ? node31385 : 4'b0011;
													assign node31385 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node31388 = (inp[5]) ? 4'b0111 : node31389;
													assign node31389 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node31393 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node31396 = (inp[15]) ? node31472 : node31397;
									assign node31397 = (inp[13]) ? node31437 : node31398;
										assign node31398 = (inp[5]) ? node31418 : node31399;
											assign node31399 = (inp[2]) ? node31403 : node31400;
												assign node31400 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node31403 = (inp[7]) ? node31415 : node31404;
													assign node31404 = (inp[9]) ? node31406 : 4'b0111;
														assign node31406 = (inp[0]) ? node31410 : node31407;
															assign node31407 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node31410 = (inp[11]) ? node31412 : 4'b0111;
																assign node31412 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node31415 = (inp[4]) ? 4'b0011 : 4'b0010;
											assign node31418 = (inp[7]) ? node31428 : node31419;
												assign node31419 = (inp[4]) ? node31423 : node31420;
													assign node31420 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node31423 = (inp[2]) ? node31425 : 4'b0010;
														assign node31425 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node31428 = (inp[4]) ? node31434 : node31429;
													assign node31429 = (inp[2]) ? 4'b0111 : node31430;
														assign node31430 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node31434 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node31437 = (inp[7]) ? node31459 : node31438;
											assign node31438 = (inp[2]) ? node31444 : node31439;
												assign node31439 = (inp[5]) ? node31441 : 4'b0010;
													assign node31441 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node31444 = (inp[4]) ? node31450 : node31445;
													assign node31445 = (inp[5]) ? 4'b0011 : node31446;
														assign node31446 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node31450 = (inp[9]) ? node31452 : 4'b0110;
														assign node31452 = (inp[11]) ? node31456 : node31453;
															assign node31453 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node31456 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node31459 = (inp[2]) ? node31467 : node31460;
												assign node31460 = (inp[4]) ? 4'b0110 : node31461;
													assign node31461 = (inp[5]) ? node31463 : 4'b0110;
														assign node31463 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node31467 = (inp[4]) ? 4'b0010 : node31468;
													assign node31468 = (inp[5]) ? 4'b0110 : 4'b0011;
									assign node31472 = (inp[7]) ? node31514 : node31473;
										assign node31473 = (inp[4]) ? node31485 : node31474;
											assign node31474 = (inp[2]) ? node31480 : node31475;
												assign node31475 = (inp[5]) ? 4'b0010 : node31476;
													assign node31476 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node31480 = (inp[5]) ? node31482 : 4'b0110;
													assign node31482 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node31485 = (inp[2]) ? node31501 : node31486;
												assign node31486 = (inp[9]) ? node31494 : node31487;
													assign node31487 = (inp[11]) ? node31491 : node31488;
														assign node31488 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node31491 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node31494 = (inp[5]) ? node31498 : node31495;
														assign node31495 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node31498 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node31501 = (inp[0]) ? node31509 : node31502;
													assign node31502 = (inp[5]) ? node31506 : node31503;
														assign node31503 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node31506 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node31509 = (inp[11]) ? 4'b0010 : node31510;
														assign node31510 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node31514 = (inp[4]) ? node31526 : node31515;
											assign node31515 = (inp[2]) ? node31521 : node31516;
												assign node31516 = (inp[11]) ? node31518 : 4'b0010;
													assign node31518 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node31521 = (inp[5]) ? 4'b0110 : node31522;
													assign node31522 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node31526 = (inp[2]) ? 4'b0010 : 4'b0110;
					assign node31529 = (inp[14]) ? node32511 : node31530;
						assign node31530 = (inp[15]) ? node32170 : node31531;
							assign node31531 = (inp[4]) ? node31893 : node31532;
								assign node31532 = (inp[5]) ? node31736 : node31533;
									assign node31533 = (inp[1]) ? node31629 : node31534;
										assign node31534 = (inp[0]) ? node31584 : node31535;
											assign node31535 = (inp[11]) ? node31555 : node31536;
												assign node31536 = (inp[9]) ? node31548 : node31537;
													assign node31537 = (inp[2]) ? node31541 : node31538;
														assign node31538 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node31541 = (inp[7]) ? node31543 : 4'b0110;
															assign node31543 = (inp[10]) ? node31545 : 4'b0011;
																assign node31545 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node31548 = (inp[7]) ? node31552 : node31549;
														assign node31549 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node31552 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node31555 = (inp[10]) ? node31569 : node31556;
													assign node31556 = (inp[9]) ? node31564 : node31557;
														assign node31557 = (inp[2]) ? node31561 : node31558;
															assign node31558 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node31561 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node31564 = (inp[7]) ? node31566 : 4'b0111;
															assign node31566 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node31569 = (inp[9]) ? node31573 : node31570;
														assign node31570 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node31573 = (inp[7]) ? node31581 : node31574;
															assign node31574 = (inp[2]) ? node31578 : node31575;
																assign node31575 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node31578 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node31581 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node31584 = (inp[9]) ? node31606 : node31585;
												assign node31585 = (inp[13]) ? node31595 : node31586;
													assign node31586 = (inp[10]) ? node31588 : 4'b0110;
														assign node31588 = (inp[7]) ? node31592 : node31589;
															assign node31589 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node31592 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node31595 = (inp[10]) ? node31603 : node31596;
														assign node31596 = (inp[7]) ? node31600 : node31597;
															assign node31597 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node31600 = (inp[2]) ? 4'b0010 : 4'b0111;
														assign node31603 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node31606 = (inp[13]) ? node31620 : node31607;
													assign node31607 = (inp[10]) ? node31615 : node31608;
														assign node31608 = (inp[2]) ? node31612 : node31609;
															assign node31609 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node31612 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node31615 = (inp[7]) ? node31617 : 4'b0111;
															assign node31617 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node31620 = (inp[2]) ? 4'b0110 : node31621;
														assign node31621 = (inp[11]) ? node31625 : node31622;
															assign node31622 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node31625 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node31629 = (inp[9]) ? node31695 : node31630;
											assign node31630 = (inp[13]) ? node31664 : node31631;
												assign node31631 = (inp[0]) ? node31645 : node31632;
													assign node31632 = (inp[11]) ? node31636 : node31633;
														assign node31633 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node31636 = (inp[2]) ? node31642 : node31637;
															assign node31637 = (inp[7]) ? 4'b0110 : node31638;
																assign node31638 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node31642 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node31645 = (inp[7]) ? node31657 : node31646;
														assign node31646 = (inp[2]) ? node31654 : node31647;
															assign node31647 = (inp[10]) ? node31651 : node31648;
																assign node31648 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node31651 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node31654 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node31657 = (inp[2]) ? node31661 : node31658;
															assign node31658 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node31661 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node31664 = (inp[7]) ? node31680 : node31665;
													assign node31665 = (inp[2]) ? node31671 : node31666;
														assign node31666 = (inp[11]) ? 4'b0010 : node31667;
															assign node31667 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node31671 = (inp[0]) ? 4'b0110 : node31672;
															assign node31672 = (inp[11]) ? node31676 : node31673;
																assign node31673 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node31676 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node31680 = (inp[2]) ? node31682 : 4'b0110;
														assign node31682 = (inp[0]) ? node31690 : node31683;
															assign node31683 = (inp[10]) ? node31687 : node31684;
																assign node31684 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node31687 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node31690 = (inp[10]) ? node31692 : 4'b0010;
																assign node31692 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node31695 = (inp[10]) ? node31717 : node31696;
												assign node31696 = (inp[7]) ? node31708 : node31697;
													assign node31697 = (inp[2]) ? node31703 : node31698;
														assign node31698 = (inp[11]) ? node31700 : 4'b0010;
															assign node31700 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node31703 = (inp[11]) ? 4'b0110 : node31704;
															assign node31704 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node31708 = (inp[2]) ? node31710 : 4'b0111;
														assign node31710 = (inp[0]) ? node31712 : 4'b0011;
															assign node31712 = (inp[11]) ? node31714 : 4'b0010;
																assign node31714 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node31717 = (inp[11]) ? node31725 : node31718;
													assign node31718 = (inp[13]) ? node31722 : node31719;
														assign node31719 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node31722 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node31725 = (inp[13]) ? node31733 : node31726;
														assign node31726 = (inp[7]) ? node31730 : node31727;
															assign node31727 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node31730 = (inp[2]) ? 4'b0010 : 4'b0111;
														assign node31733 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node31736 = (inp[0]) ? node31820 : node31737;
										assign node31737 = (inp[1]) ? node31773 : node31738;
											assign node31738 = (inp[7]) ? node31752 : node31739;
												assign node31739 = (inp[2]) ? node31747 : node31740;
													assign node31740 = (inp[11]) ? 4'b0010 : node31741;
														assign node31741 = (inp[13]) ? node31743 : 4'b0011;
															assign node31743 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node31747 = (inp[10]) ? 4'b0110 : node31748;
														assign node31748 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node31752 = (inp[2]) ? node31764 : node31753;
													assign node31753 = (inp[9]) ? 4'b0110 : node31754;
														assign node31754 = (inp[11]) ? 4'b0110 : node31755;
															assign node31755 = (inp[10]) ? node31759 : node31756;
																assign node31756 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node31759 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node31764 = (inp[9]) ? node31766 : 4'b0010;
														assign node31766 = (inp[11]) ? 4'b0011 : node31767;
															assign node31767 = (inp[13]) ? 4'b0010 : node31768;
																assign node31768 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node31773 = (inp[11]) ? node31797 : node31774;
												assign node31774 = (inp[13]) ? node31788 : node31775;
													assign node31775 = (inp[10]) ? node31781 : node31776;
														assign node31776 = (inp[2]) ? node31778 : 4'b0111;
															assign node31778 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node31781 = (inp[2]) ? node31785 : node31782;
															assign node31782 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node31785 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node31788 = (inp[10]) ? node31792 : node31789;
														assign node31789 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node31792 = (inp[2]) ? 4'b0111 : node31793;
															assign node31793 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node31797 = (inp[13]) ? node31811 : node31798;
													assign node31798 = (inp[9]) ? 4'b0010 : node31799;
														assign node31799 = (inp[10]) ? node31803 : node31800;
															assign node31800 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node31803 = (inp[7]) ? node31807 : node31804;
																assign node31804 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node31807 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node31811 = (inp[9]) ? 4'b0111 : node31812;
														assign node31812 = (inp[10]) ? node31814 : 4'b0110;
															assign node31814 = (inp[2]) ? node31816 : 4'b0010;
																assign node31816 = (inp[7]) ? 4'b0010 : 4'b0110;
										assign node31820 = (inp[13]) ? node31860 : node31821;
											assign node31821 = (inp[2]) ? node31843 : node31822;
												assign node31822 = (inp[7]) ? node31832 : node31823;
													assign node31823 = (inp[1]) ? node31825 : 4'b0010;
														assign node31825 = (inp[11]) ? node31829 : node31826;
															assign node31826 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node31829 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node31832 = (inp[1]) ? 4'b0110 : node31833;
														assign node31833 = (inp[9]) ? node31835 : 4'b0111;
															assign node31835 = (inp[10]) ? node31839 : node31836;
																assign node31836 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node31839 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node31843 = (inp[7]) ? node31851 : node31844;
													assign node31844 = (inp[9]) ? node31846 : 4'b0110;
														assign node31846 = (inp[10]) ? 4'b0111 : node31847;
															assign node31847 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node31851 = (inp[10]) ? node31857 : node31852;
														assign node31852 = (inp[11]) ? 4'b0010 : node31853;
															assign node31853 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node31857 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node31860 = (inp[10]) ? node31880 : node31861;
												assign node31861 = (inp[1]) ? node31867 : node31862;
													assign node31862 = (inp[2]) ? node31864 : 4'b0011;
														assign node31864 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node31867 = (inp[11]) ? node31873 : node31868;
														assign node31868 = (inp[9]) ? 4'b0010 : node31869;
															assign node31869 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node31873 = (inp[9]) ? node31875 : 4'b0011;
															assign node31875 = (inp[2]) ? node31877 : 4'b0110;
																assign node31877 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node31880 = (inp[7]) ? node31888 : node31881;
													assign node31881 = (inp[2]) ? 4'b0110 : node31882;
														assign node31882 = (inp[9]) ? 4'b0010 : node31883;
															assign node31883 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node31888 = (inp[2]) ? node31890 : 4'b0111;
														assign node31890 = (inp[11]) ? 4'b0010 : 4'b0011;
								assign node31893 = (inp[5]) ? node32043 : node31894;
									assign node31894 = (inp[10]) ? node31966 : node31895;
										assign node31895 = (inp[13]) ? node31939 : node31896;
											assign node31896 = (inp[0]) ? node31912 : node31897;
												assign node31897 = (inp[1]) ? node31905 : node31898;
													assign node31898 = (inp[2]) ? node31902 : node31899;
														assign node31899 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node31902 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node31905 = (inp[2]) ? node31909 : node31906;
														assign node31906 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node31909 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node31912 = (inp[9]) ? node31920 : node31913;
													assign node31913 = (inp[7]) ? node31917 : node31914;
														assign node31914 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node31917 = (inp[2]) ? 4'b0110 : 4'b0011;
													assign node31920 = (inp[1]) ? node31928 : node31921;
														assign node31921 = (inp[2]) ? node31923 : 4'b0011;
															assign node31923 = (inp[7]) ? 4'b0110 : node31924;
																assign node31924 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node31928 = (inp[7]) ? node31934 : node31929;
															assign node31929 = (inp[2]) ? 4'b0011 : node31930;
																assign node31930 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node31934 = (inp[2]) ? 4'b0110 : node31935;
																assign node31935 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node31939 = (inp[11]) ? node31951 : node31940;
												assign node31940 = (inp[2]) ? node31948 : node31941;
													assign node31941 = (inp[7]) ? node31945 : node31942;
														assign node31942 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node31945 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node31948 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node31951 = (inp[1]) ? node31959 : node31952;
													assign node31952 = (inp[2]) ? node31956 : node31953;
														assign node31953 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node31956 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node31959 = (inp[0]) ? 4'b0010 : node31960;
														assign node31960 = (inp[7]) ? node31962 : 4'b0010;
															assign node31962 = (inp[9]) ? 4'b0010 : 4'b0111;
										assign node31966 = (inp[9]) ? node32000 : node31967;
											assign node31967 = (inp[2]) ? node31987 : node31968;
												assign node31968 = (inp[7]) ? node31976 : node31969;
													assign node31969 = (inp[13]) ? node31971 : 4'b0111;
														assign node31971 = (inp[1]) ? node31973 : 4'b0110;
															assign node31973 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node31976 = (inp[13]) ? node31982 : node31977;
														assign node31977 = (inp[11]) ? 4'b0010 : node31978;
															assign node31978 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node31982 = (inp[11]) ? 4'b0011 : node31983;
															assign node31983 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node31987 = (inp[7]) ? node31991 : node31988;
													assign node31988 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node31991 = (inp[0]) ? node31993 : 4'b0111;
														assign node31993 = (inp[1]) ? node31995 : 4'b0111;
															assign node31995 = (inp[13]) ? node31997 : 4'b0110;
																assign node31997 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node32000 = (inp[1]) ? node32018 : node32001;
												assign node32001 = (inp[13]) ? node32009 : node32002;
													assign node32002 = (inp[7]) ? 4'b0010 : node32003;
														assign node32003 = (inp[2]) ? node32005 : 4'b0111;
															assign node32005 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node32009 = (inp[7]) ? node32015 : node32010;
														assign node32010 = (inp[2]) ? node32012 : 4'b0110;
															assign node32012 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node32015 = (inp[2]) ? 4'b0110 : 4'b0011;
												assign node32018 = (inp[13]) ? node32034 : node32019;
													assign node32019 = (inp[11]) ? node32029 : node32020;
														assign node32020 = (inp[0]) ? node32024 : node32021;
															assign node32021 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node32024 = (inp[7]) ? 4'b0110 : node32025;
																assign node32025 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node32029 = (inp[7]) ? node32031 : 4'b0111;
															assign node32031 = (inp[2]) ? 4'b0111 : 4'b0010;
													assign node32034 = (inp[11]) ? 4'b0011 : node32035;
														assign node32035 = (inp[7]) ? node32039 : node32036;
															assign node32036 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node32039 = (inp[2]) ? 4'b0111 : 4'b0010;
									assign node32043 = (inp[1]) ? node32115 : node32044;
										assign node32044 = (inp[10]) ? node32062 : node32045;
											assign node32045 = (inp[13]) ? node32053 : node32046;
												assign node32046 = (inp[2]) ? node32050 : node32047;
													assign node32047 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node32050 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node32053 = (inp[2]) ? node32059 : node32054;
													assign node32054 = (inp[7]) ? node32056 : 4'b0010;
														assign node32056 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node32059 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node32062 = (inp[11]) ? node32082 : node32063;
												assign node32063 = (inp[13]) ? node32075 : node32064;
													assign node32064 = (inp[0]) ? node32070 : node32065;
														assign node32065 = (inp[9]) ? 4'b0010 : node32066;
															assign node32066 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node32070 = (inp[7]) ? node32072 : 4'b0111;
															assign node32072 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node32075 = (inp[7]) ? node32079 : node32076;
														assign node32076 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node32079 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node32082 = (inp[0]) ? node32102 : node32083;
													assign node32083 = (inp[9]) ? node32089 : node32084;
														assign node32084 = (inp[2]) ? 4'b0011 : node32085;
															assign node32085 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node32089 = (inp[13]) ? node32095 : node32090;
															assign node32090 = (inp[2]) ? 4'b0111 : node32091;
																assign node32091 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node32095 = (inp[2]) ? node32099 : node32096;
																assign node32096 = (inp[7]) ? 4'b0111 : 4'b0011;
																assign node32099 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node32102 = (inp[2]) ? node32108 : node32103;
														assign node32103 = (inp[13]) ? 4'b0111 : node32104;
															assign node32104 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node32108 = (inp[7]) ? node32112 : node32109;
															assign node32109 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node32112 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node32115 = (inp[11]) ? node32143 : node32116;
											assign node32116 = (inp[2]) ? node32128 : node32117;
												assign node32117 = (inp[7]) ? node32121 : node32118;
													assign node32118 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node32121 = (inp[13]) ? node32125 : node32122;
														assign node32122 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node32125 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node32128 = (inp[7]) ? node32136 : node32129;
													assign node32129 = (inp[9]) ? 4'b0110 : node32130;
														assign node32130 = (inp[10]) ? 4'b0111 : node32131;
															assign node32131 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node32136 = (inp[10]) ? node32140 : node32137;
														assign node32137 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node32140 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node32143 = (inp[2]) ? node32153 : node32144;
												assign node32144 = (inp[7]) ? 4'b0111 : node32145;
													assign node32145 = (inp[9]) ? node32147 : 4'b0010;
														assign node32147 = (inp[0]) ? node32149 : 4'b0011;
															assign node32149 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node32153 = (inp[7]) ? node32163 : node32154;
													assign node32154 = (inp[9]) ? node32160 : node32155;
														assign node32155 = (inp[13]) ? 4'b0111 : node32156;
															assign node32156 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node32160 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node32163 = (inp[13]) ? node32167 : node32164;
														assign node32164 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node32167 = (inp[10]) ? 4'b0010 : 4'b0011;
							assign node32170 = (inp[13]) ? node32278 : node32171;
								assign node32171 = (inp[2]) ? node32211 : node32172;
									assign node32172 = (inp[5]) ? node32196 : node32173;
										assign node32173 = (inp[10]) ? node32185 : node32174;
											assign node32174 = (inp[7]) ? node32180 : node32175;
												assign node32175 = (inp[4]) ? node32177 : 4'b0000;
													assign node32177 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node32180 = (inp[4]) ? node32182 : 4'b0001;
													assign node32182 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node32185 = (inp[7]) ? node32191 : node32186;
												assign node32186 = (inp[11]) ? node32188 : 4'b0001;
													assign node32188 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node32191 = (inp[4]) ? node32193 : 4'b0000;
													assign node32193 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node32196 = (inp[7]) ? node32204 : node32197;
											assign node32197 = (inp[4]) ? node32201 : node32198;
												assign node32198 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node32201 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node32204 = (inp[10]) ? node32208 : node32205;
												assign node32205 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node32208 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node32211 = (inp[5]) ? node32235 : node32212;
										assign node32212 = (inp[10]) ? node32224 : node32213;
											assign node32213 = (inp[7]) ? node32219 : node32214;
												assign node32214 = (inp[4]) ? node32216 : 4'b0100;
													assign node32216 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node32219 = (inp[11]) ? 4'b0101 : node32220;
													assign node32220 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node32224 = (inp[7]) ? node32230 : node32225;
												assign node32225 = (inp[11]) ? 4'b0101 : node32226;
													assign node32226 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node32230 = (inp[11]) ? 4'b0100 : node32231;
													assign node32231 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node32235 = (inp[0]) ? node32271 : node32236;
											assign node32236 = (inp[1]) ? node32256 : node32237;
												assign node32237 = (inp[9]) ? node32245 : node32238;
													assign node32238 = (inp[10]) ? node32242 : node32239;
														assign node32239 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node32242 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node32245 = (inp[7]) ? node32247 : 4'b0000;
														assign node32247 = (inp[4]) ? 4'b0000 : node32248;
															assign node32248 = (inp[10]) ? node32252 : node32249;
																assign node32249 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node32252 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node32256 = (inp[9]) ? node32264 : node32257;
													assign node32257 = (inp[4]) ? node32259 : 4'b0001;
														assign node32259 = (inp[11]) ? node32261 : 4'b0001;
															assign node32261 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node32264 = (inp[10]) ? node32268 : node32265;
														assign node32265 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node32268 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node32271 = (inp[10]) ? node32275 : node32272;
												assign node32272 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node32275 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node32278 = (inp[0]) ? node32412 : node32279;
									assign node32279 = (inp[7]) ? node32359 : node32280;
										assign node32280 = (inp[10]) ? node32310 : node32281;
											assign node32281 = (inp[4]) ? node32297 : node32282;
												assign node32282 = (inp[11]) ? node32292 : node32283;
													assign node32283 = (inp[1]) ? node32289 : node32284;
														assign node32284 = (inp[2]) ? 4'b0100 : node32285;
															assign node32285 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node32289 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node32292 = (inp[2]) ? 4'b0001 : node32293;
														assign node32293 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node32297 = (inp[5]) ? node32305 : node32298;
													assign node32298 = (inp[2]) ? node32302 : node32299;
														assign node32299 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node32302 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node32305 = (inp[2]) ? node32307 : 4'b0101;
														assign node32307 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node32310 = (inp[4]) ? node32340 : node32311;
												assign node32311 = (inp[1]) ? node32333 : node32312;
													assign node32312 = (inp[11]) ? node32326 : node32313;
														assign node32313 = (inp[9]) ? node32321 : node32314;
															assign node32314 = (inp[5]) ? node32318 : node32315;
																assign node32315 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node32318 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node32321 = (inp[2]) ? 4'b0101 : node32322;
																assign node32322 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node32326 = (inp[2]) ? node32330 : node32327;
															assign node32327 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node32330 = (inp[5]) ? 4'b0000 : 4'b0101;
													assign node32333 = (inp[11]) ? node32335 : 4'b0001;
														assign node32335 = (inp[2]) ? 4'b0101 : node32336;
															assign node32336 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node32340 = (inp[1]) ? node32348 : node32341;
													assign node32341 = (inp[5]) ? 4'b0001 : node32342;
														assign node32342 = (inp[2]) ? node32344 : 4'b0001;
															assign node32344 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node32348 = (inp[5]) ? node32356 : node32349;
														assign node32349 = (inp[2]) ? node32353 : node32350;
															assign node32350 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node32353 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node32356 = (inp[2]) ? 4'b0000 : 4'b0100;
										assign node32359 = (inp[10]) ? node32399 : node32360;
											assign node32360 = (inp[9]) ? node32376 : node32361;
												assign node32361 = (inp[1]) ? node32371 : node32362;
													assign node32362 = (inp[2]) ? node32368 : node32363;
														assign node32363 = (inp[5]) ? 4'b0101 : node32364;
															assign node32364 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node32368 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node32371 = (inp[4]) ? 4'b0101 : node32372;
														assign node32372 = (inp[5]) ? 4'b0100 : 4'b0001;
												assign node32376 = (inp[4]) ? node32382 : node32377;
													assign node32377 = (inp[5]) ? 4'b0100 : node32378;
														assign node32378 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node32382 = (inp[1]) ? node32394 : node32383;
														assign node32383 = (inp[2]) ? node32389 : node32384;
															assign node32384 = (inp[5]) ? 4'b0101 : node32385;
																assign node32385 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node32389 = (inp[5]) ? node32391 : 4'b0101;
																assign node32391 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node32394 = (inp[2]) ? node32396 : 4'b0000;
															assign node32396 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node32399 = (inp[5]) ? node32405 : node32400;
												assign node32400 = (inp[2]) ? 4'b0100 : node32401;
													assign node32401 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node32405 = (inp[2]) ? node32409 : node32406;
													assign node32406 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node32409 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node32412 = (inp[10]) ? node32470 : node32413;
										assign node32413 = (inp[7]) ? node32441 : node32414;
											assign node32414 = (inp[4]) ? node32428 : node32415;
												assign node32415 = (inp[9]) ? node32421 : node32416;
													assign node32416 = (inp[5]) ? 4'b0001 : node32417;
														assign node32417 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node32421 = (inp[5]) ? node32425 : node32422;
														assign node32422 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node32425 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node32428 = (inp[11]) ? node32434 : node32429;
													assign node32429 = (inp[9]) ? node32431 : 4'b0000;
														assign node32431 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node32434 = (inp[2]) ? node32438 : node32435;
														assign node32435 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node32438 = (inp[5]) ? 4'b0001 : 4'b0100;
											assign node32441 = (inp[1]) ? node32457 : node32442;
												assign node32442 = (inp[11]) ? node32450 : node32443;
													assign node32443 = (inp[5]) ? node32445 : 4'b0001;
														assign node32445 = (inp[2]) ? 4'b0000 : node32446;
															assign node32446 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node32450 = (inp[5]) ? node32454 : node32451;
														assign node32451 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node32454 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node32457 = (inp[2]) ? node32465 : node32458;
													assign node32458 = (inp[5]) ? node32462 : node32459;
														assign node32459 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node32462 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node32465 = (inp[5]) ? node32467 : 4'b0101;
														assign node32467 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node32470 = (inp[11]) ? node32494 : node32471;
											assign node32471 = (inp[5]) ? node32489 : node32472;
												assign node32472 = (inp[2]) ? node32476 : node32473;
													assign node32473 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node32476 = (inp[1]) ? node32484 : node32477;
														assign node32477 = (inp[7]) ? node32481 : node32478;
															assign node32478 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node32481 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node32484 = (inp[4]) ? 4'b0101 : node32485;
															assign node32485 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node32489 = (inp[2]) ? 4'b0001 : node32490;
													assign node32490 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node32494 = (inp[5]) ? node32506 : node32495;
												assign node32495 = (inp[2]) ? node32503 : node32496;
													assign node32496 = (inp[4]) ? node32500 : node32497;
														assign node32497 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node32500 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node32503 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node32506 = (inp[2]) ? 4'b0000 : node32507;
													assign node32507 = (inp[4]) ? 4'b0100 : 4'b0101;
						assign node32511 = (inp[2]) ? node33005 : node32512;
							assign node32512 = (inp[15]) ? node32776 : node32513;
								assign node32513 = (inp[7]) ? node32621 : node32514;
									assign node32514 = (inp[4]) ? node32578 : node32515;
										assign node32515 = (inp[5]) ? node32559 : node32516;
											assign node32516 = (inp[0]) ? node32536 : node32517;
												assign node32517 = (inp[1]) ? node32527 : node32518;
													assign node32518 = (inp[9]) ? 4'b0101 : node32519;
														assign node32519 = (inp[13]) ? node32521 : 4'b0100;
															assign node32521 = (inp[10]) ? node32523 : 4'b0101;
																assign node32523 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node32527 = (inp[9]) ? 4'b0100 : node32528;
														assign node32528 = (inp[13]) ? node32532 : node32529;
															assign node32529 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node32532 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node32536 = (inp[10]) ? node32548 : node32537;
													assign node32537 = (inp[9]) ? 4'b0100 : node32538;
														assign node32538 = (inp[1]) ? node32544 : node32539;
															assign node32539 = (inp[11]) ? 4'b0100 : node32540;
																assign node32540 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node32544 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node32548 = (inp[13]) ? node32554 : node32549;
														assign node32549 = (inp[11]) ? 4'b0100 : node32550;
															assign node32550 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node32554 = (inp[1]) ? 4'b0101 : node32555;
															assign node32555 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node32559 = (inp[10]) ? node32567 : node32560;
												assign node32560 = (inp[13]) ? node32562 : 4'b0000;
													assign node32562 = (inp[11]) ? node32564 : 4'b0001;
														assign node32564 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node32567 = (inp[13]) ? node32573 : node32568;
													assign node32568 = (inp[1]) ? node32570 : 4'b0001;
														assign node32570 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node32573 = (inp[11]) ? node32575 : 4'b0000;
														assign node32575 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node32578 = (inp[10]) ? node32602 : node32579;
											assign node32579 = (inp[5]) ? node32591 : node32580;
												assign node32580 = (inp[13]) ? node32586 : node32581;
													assign node32581 = (inp[1]) ? node32583 : 4'b0000;
														assign node32583 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node32586 = (inp[1]) ? node32588 : 4'b0001;
														assign node32588 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node32591 = (inp[13]) ? node32597 : node32592;
													assign node32592 = (inp[11]) ? node32594 : 4'b0001;
														assign node32594 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node32597 = (inp[11]) ? node32599 : 4'b0000;
														assign node32599 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node32602 = (inp[13]) ? node32610 : node32603;
												assign node32603 = (inp[5]) ? 4'b0000 : node32604;
													assign node32604 = (inp[11]) ? node32606 : 4'b0001;
														assign node32606 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node32610 = (inp[5]) ? node32616 : node32611;
													assign node32611 = (inp[1]) ? node32613 : 4'b0000;
														assign node32613 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node32616 = (inp[11]) ? node32618 : 4'b0001;
														assign node32618 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node32621 = (inp[4]) ? node32699 : node32622;
										assign node32622 = (inp[5]) ? node32652 : node32623;
											assign node32623 = (inp[13]) ? node32631 : node32624;
												assign node32624 = (inp[10]) ? 4'b0001 : node32625;
													assign node32625 = (inp[1]) ? 4'b0000 : node32626;
														assign node32626 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node32631 = (inp[9]) ? node32643 : node32632;
													assign node32632 = (inp[11]) ? 4'b0001 : node32633;
														assign node32633 = (inp[0]) ? 4'b0000 : node32634;
															assign node32634 = (inp[10]) ? node32638 : node32635;
																assign node32635 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node32638 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node32643 = (inp[10]) ? node32647 : node32644;
														assign node32644 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node32647 = (inp[1]) ? 4'b0000 : node32648;
															assign node32648 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node32652 = (inp[9]) ? node32674 : node32653;
												assign node32653 = (inp[13]) ? node32665 : node32654;
													assign node32654 = (inp[10]) ? node32660 : node32655;
														assign node32655 = (inp[11]) ? 4'b0101 : node32656;
															assign node32656 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node32660 = (inp[11]) ? 4'b0100 : node32661;
															assign node32661 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node32665 = (inp[10]) ? node32669 : node32666;
														assign node32666 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node32669 = (inp[11]) ? 4'b0101 : node32670;
															assign node32670 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node32674 = (inp[0]) ? node32690 : node32675;
													assign node32675 = (inp[11]) ? 4'b0100 : node32676;
														assign node32676 = (inp[1]) ? node32682 : node32677;
															assign node32677 = (inp[10]) ? 4'b0101 : node32678;
																assign node32678 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node32682 = (inp[13]) ? node32686 : node32683;
																assign node32683 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node32686 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node32690 = (inp[11]) ? 4'b0101 : node32691;
														assign node32691 = (inp[10]) ? node32695 : node32692;
															assign node32692 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node32695 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node32699 = (inp[5]) ? node32735 : node32700;
											assign node32700 = (inp[9]) ? node32712 : node32701;
												assign node32701 = (inp[10]) ? node32703 : 4'b0101;
													assign node32703 = (inp[13]) ? node32707 : node32704;
														assign node32704 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node32707 = (inp[1]) ? 4'b0100 : node32708;
															assign node32708 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node32712 = (inp[10]) ? node32724 : node32713;
													assign node32713 = (inp[13]) ? node32719 : node32714;
														assign node32714 = (inp[11]) ? 4'b0100 : node32715;
															assign node32715 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node32719 = (inp[1]) ? 4'b0101 : node32720;
															assign node32720 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node32724 = (inp[13]) ? node32730 : node32725;
														assign node32725 = (inp[11]) ? 4'b0101 : node32726;
															assign node32726 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node32730 = (inp[0]) ? 4'b0100 : node32731;
															assign node32731 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node32735 = (inp[9]) ? node32761 : node32736;
												assign node32736 = (inp[0]) ? node32750 : node32737;
													assign node32737 = (inp[13]) ? node32741 : node32738;
														assign node32738 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node32741 = (inp[1]) ? node32747 : node32742;
															assign node32742 = (inp[10]) ? node32744 : 4'b0100;
																assign node32744 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node32747 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node32750 = (inp[1]) ? node32756 : node32751;
														assign node32751 = (inp[11]) ? 4'b0100 : node32752;
															assign node32752 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node32756 = (inp[11]) ? 4'b0101 : node32757;
															assign node32757 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node32761 = (inp[13]) ? node32767 : node32762;
													assign node32762 = (inp[10]) ? node32764 : 4'b0100;
														assign node32764 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node32767 = (inp[10]) ? node32771 : node32768;
														assign node32768 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node32771 = (inp[11]) ? 4'b0100 : node32772;
															assign node32772 = (inp[0]) ? 4'b0100 : 4'b0101;
								assign node32776 = (inp[13]) ? node32864 : node32777;
									assign node32777 = (inp[11]) ? node32797 : node32778;
										assign node32778 = (inp[10]) ? node32786 : node32779;
											assign node32779 = (inp[7]) ? node32781 : 4'b0100;
												assign node32781 = (inp[4]) ? 4'b0101 : node32782;
													assign node32782 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node32786 = (inp[7]) ? node32792 : node32787;
												assign node32787 = (inp[5]) ? node32789 : 4'b0101;
													assign node32789 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node32792 = (inp[4]) ? 4'b0100 : node32793;
													assign node32793 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node32797 = (inp[5]) ? node32841 : node32798;
											assign node32798 = (inp[9]) ? node32816 : node32799;
												assign node32799 = (inp[10]) ? node32809 : node32800;
													assign node32800 = (inp[0]) ? node32802 : 4'b0100;
														assign node32802 = (inp[1]) ? 4'b0100 : node32803;
															assign node32803 = (inp[4]) ? 4'b0100 : node32804;
																assign node32804 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node32809 = (inp[4]) ? node32813 : node32810;
														assign node32810 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node32813 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node32816 = (inp[10]) ? node32826 : node32817;
													assign node32817 = (inp[1]) ? 4'b0101 : node32818;
														assign node32818 = (inp[7]) ? node32822 : node32819;
															assign node32819 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node32822 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node32826 = (inp[1]) ? node32836 : node32827;
														assign node32827 = (inp[0]) ? node32829 : 4'b0100;
															assign node32829 = (inp[7]) ? node32833 : node32830;
																assign node32830 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node32833 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node32836 = (inp[4]) ? 4'b0101 : node32837;
															assign node32837 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node32841 = (inp[0]) ? node32849 : node32842;
												assign node32842 = (inp[10]) ? node32846 : node32843;
													assign node32843 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node32846 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node32849 = (inp[1]) ? node32857 : node32850;
													assign node32850 = (inp[4]) ? node32854 : node32851;
														assign node32851 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node32854 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node32857 = (inp[9]) ? node32859 : 4'b0101;
														assign node32859 = (inp[4]) ? node32861 : 4'b0101;
															assign node32861 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node32864 = (inp[0]) ? node32918 : node32865;
										assign node32865 = (inp[9]) ? node32895 : node32866;
											assign node32866 = (inp[7]) ? node32880 : node32867;
												assign node32867 = (inp[11]) ? node32873 : node32868;
													assign node32868 = (inp[5]) ? 4'b0101 : node32869;
														assign node32869 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node32873 = (inp[4]) ? 4'b0100 : node32874;
														assign node32874 = (inp[5]) ? 4'b0100 : node32875;
															assign node32875 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node32880 = (inp[10]) ? node32888 : node32881;
													assign node32881 = (inp[4]) ? 4'b0101 : node32882;
														assign node32882 = (inp[11]) ? 4'b0100 : node32883;
															assign node32883 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node32888 = (inp[4]) ? 4'b0100 : node32889;
														assign node32889 = (inp[11]) ? 4'b0101 : node32890;
															assign node32890 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node32895 = (inp[4]) ? node32907 : node32896;
												assign node32896 = (inp[10]) ? node32900 : node32897;
													assign node32897 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node32900 = (inp[7]) ? 4'b0101 : node32901;
														assign node32901 = (inp[11]) ? node32903 : 4'b0101;
															assign node32903 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node32907 = (inp[10]) ? node32913 : node32908;
													assign node32908 = (inp[5]) ? 4'b0101 : node32909;
														assign node32909 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node32913 = (inp[5]) ? 4'b0100 : node32914;
														assign node32914 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node32918 = (inp[11]) ? node32968 : node32919;
											assign node32919 = (inp[1]) ? node32941 : node32920;
												assign node32920 = (inp[9]) ? node32930 : node32921;
													assign node32921 = (inp[5]) ? 4'b0101 : node32922;
														assign node32922 = (inp[4]) ? 4'b0100 : node32923;
															assign node32923 = (inp[7]) ? 4'b0101 : node32924;
																assign node32924 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node32930 = (inp[4]) ? node32932 : 4'b0100;
														assign node32932 = (inp[5]) ? 4'b0100 : node32933;
															assign node32933 = (inp[7]) ? node32937 : node32934;
																assign node32934 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node32937 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node32941 = (inp[5]) ? node32963 : node32942;
													assign node32942 = (inp[4]) ? node32954 : node32943;
														assign node32943 = (inp[9]) ? node32949 : node32944;
															assign node32944 = (inp[10]) ? 4'b0101 : node32945;
																assign node32945 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node32949 = (inp[10]) ? node32951 : 4'b0101;
																assign node32951 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node32954 = (inp[9]) ? node32958 : node32955;
															assign node32955 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node32958 = (inp[7]) ? node32960 : 4'b0100;
																assign node32960 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node32963 = (inp[4]) ? 4'b0101 : node32964;
														assign node32964 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node32968 = (inp[5]) ? node32998 : node32969;
												assign node32969 = (inp[10]) ? node32993 : node32970;
													assign node32970 = (inp[9]) ? node32980 : node32971;
														assign node32971 = (inp[1]) ? node32973 : 4'b0100;
															assign node32973 = (inp[7]) ? node32977 : node32974;
																assign node32974 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node32977 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node32980 = (inp[1]) ? node32988 : node32981;
															assign node32981 = (inp[4]) ? node32985 : node32982;
																assign node32982 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node32985 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node32988 = (inp[7]) ? node32990 : 4'b0100;
																assign node32990 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node32993 = (inp[7]) ? 4'b0100 : node32994;
														assign node32994 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node32998 = (inp[1]) ? node33000 : 4'b0100;
													assign node33000 = (inp[10]) ? node33002 : 4'b0100;
														assign node33002 = (inp[4]) ? 4'b0100 : 4'b0101;
							assign node33005 = (inp[15]) ? node33321 : node33006;
								assign node33006 = (inp[7]) ? node33144 : node33007;
									assign node33007 = (inp[4]) ? node33089 : node33008;
										assign node33008 = (inp[5]) ? node33060 : node33009;
											assign node33009 = (inp[9]) ? node33035 : node33010;
												assign node33010 = (inp[11]) ? node33018 : node33011;
													assign node33011 = (inp[10]) ? node33013 : 4'b0000;
														assign node33013 = (inp[13]) ? 4'b0000 : node33014;
															assign node33014 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node33018 = (inp[0]) ? node33030 : node33019;
														assign node33019 = (inp[1]) ? node33025 : node33020;
															assign node33020 = (inp[13]) ? 4'b0001 : node33021;
																assign node33021 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node33025 = (inp[13]) ? node33027 : 4'b0001;
																assign node33027 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node33030 = (inp[13]) ? node33032 : 4'b0000;
															assign node33032 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node33035 = (inp[11]) ? node33045 : node33036;
													assign node33036 = (inp[1]) ? 4'b0001 : node33037;
														assign node33037 = (inp[10]) ? node33041 : node33038;
															assign node33038 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33041 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node33045 = (inp[1]) ? node33051 : node33046;
														assign node33046 = (inp[13]) ? 4'b0001 : node33047;
															assign node33047 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node33051 = (inp[0]) ? 4'b0000 : node33052;
															assign node33052 = (inp[13]) ? node33056 : node33053;
																assign node33053 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node33056 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node33060 = (inp[9]) ? node33082 : node33061;
												assign node33061 = (inp[11]) ? node33079 : node33062;
													assign node33062 = (inp[1]) ? node33070 : node33063;
														assign node33063 = (inp[0]) ? 4'b0100 : node33064;
															assign node33064 = (inp[10]) ? node33066 : 4'b0101;
																assign node33066 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node33070 = (inp[0]) ? node33074 : node33071;
															assign node33071 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node33074 = (inp[10]) ? node33076 : 4'b0101;
																assign node33076 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node33079 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node33082 = (inp[10]) ? node33086 : node33083;
													assign node33083 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node33086 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node33089 = (inp[1]) ? node33121 : node33090;
											assign node33090 = (inp[0]) ? node33104 : node33091;
												assign node33091 = (inp[9]) ? 4'b0100 : node33092;
													assign node33092 = (inp[11]) ? node33098 : node33093;
														assign node33093 = (inp[10]) ? 4'b0100 : node33094;
															assign node33094 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node33098 = (inp[13]) ? node33100 : 4'b0101;
															assign node33100 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node33104 = (inp[10]) ? node33114 : node33105;
													assign node33105 = (inp[13]) ? node33107 : 4'b0100;
														assign node33107 = (inp[11]) ? node33111 : node33108;
															assign node33108 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node33111 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node33114 = (inp[9]) ? node33116 : 4'b0100;
														assign node33116 = (inp[13]) ? node33118 : 4'b0101;
															assign node33118 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node33121 = (inp[13]) ? node33137 : node33122;
												assign node33122 = (inp[0]) ? node33130 : node33123;
													assign node33123 = (inp[5]) ? node33127 : node33124;
														assign node33124 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node33127 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node33130 = (inp[11]) ? 4'b0100 : node33131;
														assign node33131 = (inp[5]) ? node33133 : 4'b0100;
															assign node33133 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node33137 = (inp[5]) ? node33141 : node33138;
													assign node33138 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node33141 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node33144 = (inp[4]) ? node33220 : node33145;
										assign node33145 = (inp[5]) ? node33185 : node33146;
											assign node33146 = (inp[1]) ? node33162 : node33147;
												assign node33147 = (inp[0]) ? node33155 : node33148;
													assign node33148 = (inp[10]) ? node33152 : node33149;
														assign node33149 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node33152 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node33155 = (inp[10]) ? node33159 : node33156;
														assign node33156 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node33159 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node33162 = (inp[11]) ? node33168 : node33163;
													assign node33163 = (inp[10]) ? 4'b0101 : node33164;
														assign node33164 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node33168 = (inp[9]) ? node33180 : node33169;
														assign node33169 = (inp[0]) ? node33175 : node33170;
															assign node33170 = (inp[13]) ? node33172 : 4'b0100;
																assign node33172 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node33175 = (inp[10]) ? node33177 : 4'b0101;
																assign node33177 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node33180 = (inp[13]) ? 4'b0101 : node33181;
															assign node33181 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node33185 = (inp[9]) ? node33215 : node33186;
												assign node33186 = (inp[0]) ? node33206 : node33187;
													assign node33187 = (inp[11]) ? node33199 : node33188;
														assign node33188 = (inp[1]) ? node33194 : node33189;
															assign node33189 = (inp[13]) ? node33191 : 4'b0001;
																assign node33191 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node33194 = (inp[10]) ? 4'b0000 : node33195;
																assign node33195 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node33199 = (inp[1]) ? node33201 : 4'b0000;
															assign node33201 = (inp[13]) ? 4'b0001 : node33202;
																assign node33202 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node33206 = (inp[10]) ? 4'b0000 : node33207;
														assign node33207 = (inp[11]) ? node33211 : node33208;
															assign node33208 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33211 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node33215 = (inp[10]) ? 4'b0001 : node33216;
													assign node33216 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node33220 = (inp[11]) ? node33286 : node33221;
											assign node33221 = (inp[9]) ? node33257 : node33222;
												assign node33222 = (inp[13]) ? node33242 : node33223;
													assign node33223 = (inp[5]) ? node33233 : node33224;
														assign node33224 = (inp[0]) ? node33226 : 4'b0001;
															assign node33226 = (inp[10]) ? node33230 : node33227;
																assign node33227 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node33230 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node33233 = (inp[0]) ? 4'b0001 : node33234;
															assign node33234 = (inp[1]) ? node33238 : node33235;
																assign node33235 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node33238 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node33242 = (inp[5]) ? node33250 : node33243;
														assign node33243 = (inp[1]) ? node33247 : node33244;
															assign node33244 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node33247 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node33250 = (inp[10]) ? node33254 : node33251;
															assign node33251 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node33254 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node33257 = (inp[13]) ? node33273 : node33258;
													assign node33258 = (inp[0]) ? node33260 : 4'b0000;
														assign node33260 = (inp[5]) ? node33266 : node33261;
															assign node33261 = (inp[10]) ? 4'b0000 : node33262;
																assign node33262 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node33266 = (inp[1]) ? node33270 : node33267;
																assign node33267 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node33270 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node33273 = (inp[0]) ? node33279 : node33274;
														assign node33274 = (inp[10]) ? 4'b0001 : node33275;
															assign node33275 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node33279 = (inp[1]) ? node33283 : node33280;
															assign node33280 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node33283 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node33286 = (inp[9]) ? node33294 : node33287;
												assign node33287 = (inp[13]) ? node33291 : node33288;
													assign node33288 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node33291 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node33294 = (inp[0]) ? node33314 : node33295;
													assign node33295 = (inp[5]) ? node33301 : node33296;
														assign node33296 = (inp[1]) ? 4'b0001 : node33297;
															assign node33297 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node33301 = (inp[1]) ? node33309 : node33302;
															assign node33302 = (inp[10]) ? node33306 : node33303;
																assign node33303 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node33306 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33309 = (inp[10]) ? node33311 : 4'b0000;
																assign node33311 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node33314 = (inp[13]) ? node33318 : node33315;
														assign node33315 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node33318 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node33321 = (inp[10]) ? node33335 : node33322;
									assign node33322 = (inp[5]) ? 4'b0001 : node33323;
										assign node33323 = (inp[7]) ? node33329 : node33324;
											assign node33324 = (inp[4]) ? 4'b0000 : node33325;
												assign node33325 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node33329 = (inp[4]) ? 4'b0001 : node33330;
												assign node33330 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node33335 = (inp[5]) ? 4'b0000 : node33336;
										assign node33336 = (inp[7]) ? node33342 : node33337;
											assign node33337 = (inp[11]) ? 4'b0001 : node33338;
												assign node33338 = (inp[4]) ? 4'b0001 : 4'b0000;
											assign node33342 = (inp[4]) ? 4'b0000 : node33343;
												assign node33343 = (inp[11]) ? 4'b0000 : 4'b0001;
				assign node33348 = (inp[15]) ? node34460 : node33349;
					assign node33349 = (inp[14]) ? node34139 : node33350;
						assign node33350 = (inp[9]) ? node33742 : node33351;
							assign node33351 = (inp[5]) ? node33529 : node33352;
								assign node33352 = (inp[7]) ? node33432 : node33353;
									assign node33353 = (inp[11]) ? node33399 : node33354;
										assign node33354 = (inp[13]) ? node33378 : node33355;
											assign node33355 = (inp[2]) ? node33363 : node33356;
												assign node33356 = (inp[4]) ? 4'b0010 : node33357;
													assign node33357 = (inp[1]) ? node33359 : 4'b0010;
														assign node33359 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node33363 = (inp[12]) ? node33373 : node33364;
													assign node33364 = (inp[0]) ? node33370 : node33365;
														assign node33365 = (inp[4]) ? 4'b0010 : node33366;
															assign node33366 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node33370 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node33373 = (inp[4]) ? node33375 : 4'b0010;
														assign node33375 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node33378 = (inp[1]) ? node33384 : node33379;
												assign node33379 = (inp[4]) ? node33381 : 4'b0011;
													assign node33381 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node33384 = (inp[10]) ? node33394 : node33385;
													assign node33385 = (inp[12]) ? node33387 : 4'b0011;
														assign node33387 = (inp[2]) ? node33391 : node33388;
															assign node33388 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node33391 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node33394 = (inp[12]) ? 4'b0010 : node33395;
														assign node33395 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node33399 = (inp[13]) ? node33413 : node33400;
											assign node33400 = (inp[1]) ? node33402 : 4'b0011;
												assign node33402 = (inp[4]) ? node33410 : node33403;
													assign node33403 = (inp[0]) ? 4'b0011 : node33404;
														assign node33404 = (inp[10]) ? node33406 : 4'b0010;
															assign node33406 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node33410 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node33413 = (inp[1]) ? node33421 : node33414;
												assign node33414 = (inp[2]) ? node33416 : 4'b0010;
													assign node33416 = (inp[12]) ? 4'b0010 : node33417;
														assign node33417 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node33421 = (inp[12]) ? node33425 : node33422;
													assign node33422 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node33425 = (inp[0]) ? 4'b0011 : node33426;
														assign node33426 = (inp[10]) ? node33428 : 4'b0011;
															assign node33428 = (inp[4]) ? 4'b0011 : 4'b0010;
									assign node33432 = (inp[11]) ? node33482 : node33433;
										assign node33433 = (inp[13]) ? node33461 : node33434;
											assign node33434 = (inp[2]) ? node33442 : node33435;
												assign node33435 = (inp[4]) ? node33437 : 4'b0110;
													assign node33437 = (inp[1]) ? 4'b0110 : node33438;
														assign node33438 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node33442 = (inp[12]) ? node33458 : node33443;
													assign node33443 = (inp[10]) ? node33449 : node33444;
														assign node33444 = (inp[4]) ? 4'b0111 : node33445;
															assign node33445 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node33449 = (inp[0]) ? node33453 : node33450;
															assign node33450 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node33453 = (inp[4]) ? 4'b0110 : node33454;
																assign node33454 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node33458 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node33461 = (inp[2]) ? node33469 : node33462;
												assign node33462 = (inp[12]) ? node33464 : 4'b0111;
													assign node33464 = (inp[4]) ? node33466 : 4'b0111;
														assign node33466 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node33469 = (inp[1]) ? node33477 : node33470;
													assign node33470 = (inp[12]) ? node33474 : node33471;
														assign node33471 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node33474 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node33477 = (inp[12]) ? 4'b0111 : node33478;
														assign node33478 = (inp[4]) ? 4'b0111 : 4'b0110;
										assign node33482 = (inp[13]) ? node33504 : node33483;
											assign node33483 = (inp[1]) ? node33497 : node33484;
												assign node33484 = (inp[0]) ? node33486 : 4'b0110;
													assign node33486 = (inp[2]) ? node33492 : node33487;
														assign node33487 = (inp[10]) ? node33489 : 4'b0111;
															assign node33489 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node33492 = (inp[12]) ? node33494 : 4'b0110;
															assign node33494 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node33497 = (inp[4]) ? 4'b0111 : node33498;
													assign node33498 = (inp[12]) ? 4'b0111 : node33499;
														assign node33499 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node33504 = (inp[2]) ? node33514 : node33505;
												assign node33505 = (inp[10]) ? 4'b0110 : node33506;
													assign node33506 = (inp[12]) ? node33508 : 4'b0110;
														assign node33508 = (inp[1]) ? 4'b0110 : node33509;
															assign node33509 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node33514 = (inp[12]) ? node33524 : node33515;
													assign node33515 = (inp[10]) ? 4'b0111 : node33516;
														assign node33516 = (inp[0]) ? 4'b0110 : node33517;
															assign node33517 = (inp[1]) ? node33519 : 4'b0111;
																assign node33519 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node33524 = (inp[1]) ? 4'b0110 : node33525;
														assign node33525 = (inp[10]) ? 4'b0111 : 4'b0110;
								assign node33529 = (inp[7]) ? node33623 : node33530;
									assign node33530 = (inp[2]) ? node33584 : node33531;
										assign node33531 = (inp[11]) ? node33559 : node33532;
											assign node33532 = (inp[13]) ? node33546 : node33533;
												assign node33533 = (inp[4]) ? node33539 : node33534;
													assign node33534 = (inp[12]) ? node33536 : 4'b0110;
														assign node33536 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node33539 = (inp[1]) ? node33543 : node33540;
														assign node33540 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node33543 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node33546 = (inp[12]) ? node33552 : node33547;
													assign node33547 = (inp[1]) ? node33549 : 4'b0111;
														assign node33549 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node33552 = (inp[4]) ? node33556 : node33553;
														assign node33553 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node33556 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node33559 = (inp[13]) ? node33573 : node33560;
												assign node33560 = (inp[4]) ? node33566 : node33561;
													assign node33561 = (inp[12]) ? node33563 : 4'b0111;
														assign node33563 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node33566 = (inp[1]) ? node33570 : node33567;
														assign node33567 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node33570 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node33573 = (inp[4]) ? node33579 : node33574;
													assign node33574 = (inp[12]) ? node33576 : 4'b0110;
														assign node33576 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node33579 = (inp[1]) ? node33581 : 4'b0111;
														assign node33581 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node33584 = (inp[10]) ? node33606 : node33585;
											assign node33585 = (inp[13]) ? node33595 : node33586;
												assign node33586 = (inp[11]) ? node33588 : 4'b0110;
													assign node33588 = (inp[1]) ? node33590 : 4'b0111;
														assign node33590 = (inp[12]) ? 4'b0111 : node33591;
															assign node33591 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node33595 = (inp[11]) ? node33601 : node33596;
													assign node33596 = (inp[12]) ? 4'b0111 : node33597;
														assign node33597 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node33601 = (inp[1]) ? node33603 : 4'b0110;
														assign node33603 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node33606 = (inp[13]) ? node33612 : node33607;
												assign node33607 = (inp[11]) ? node33609 : 4'b0110;
													assign node33609 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node33612 = (inp[11]) ? node33618 : node33613;
													assign node33613 = (inp[4]) ? 4'b0111 : node33614;
														assign node33614 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node33618 = (inp[0]) ? node33620 : 4'b0110;
														assign node33620 = (inp[4]) ? 4'b0110 : 4'b0111;
									assign node33623 = (inp[2]) ? node33711 : node33624;
										assign node33624 = (inp[0]) ? node33662 : node33625;
											assign node33625 = (inp[1]) ? node33649 : node33626;
												assign node33626 = (inp[4]) ? node33636 : node33627;
													assign node33627 = (inp[13]) ? 4'b0010 : node33628;
														assign node33628 = (inp[12]) ? node33632 : node33629;
															assign node33629 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node33632 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node33636 = (inp[13]) ? node33644 : node33637;
														assign node33637 = (inp[12]) ? node33641 : node33638;
															assign node33638 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node33641 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node33644 = (inp[12]) ? node33646 : 4'b0011;
															assign node33646 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node33649 = (inp[11]) ? node33655 : node33650;
													assign node33650 = (inp[10]) ? node33652 : 4'b0011;
														assign node33652 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node33655 = (inp[12]) ? node33657 : 4'b0010;
														assign node33657 = (inp[13]) ? 4'b0011 : node33658;
															assign node33658 = (inp[4]) ? 4'b0011 : 4'b0010;
											assign node33662 = (inp[12]) ? node33686 : node33663;
												assign node33663 = (inp[10]) ? node33671 : node33664;
													assign node33664 = (inp[4]) ? 4'b0011 : node33665;
														assign node33665 = (inp[11]) ? node33667 : 4'b0011;
															assign node33667 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node33671 = (inp[4]) ? node33679 : node33672;
														assign node33672 = (inp[1]) ? 4'b0011 : node33673;
															assign node33673 = (inp[11]) ? node33675 : 4'b0011;
																assign node33675 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node33679 = (inp[1]) ? node33681 : 4'b0011;
															assign node33681 = (inp[11]) ? 4'b0010 : node33682;
																assign node33682 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node33686 = (inp[4]) ? node33700 : node33687;
													assign node33687 = (inp[1]) ? node33693 : node33688;
														assign node33688 = (inp[10]) ? 4'b0011 : node33689;
															assign node33689 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node33693 = (inp[11]) ? node33697 : node33694;
															assign node33694 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node33697 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node33700 = (inp[13]) ? node33706 : node33701;
														assign node33701 = (inp[1]) ? 4'b0011 : node33702;
															assign node33702 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node33706 = (inp[11]) ? node33708 : 4'b0010;
															assign node33708 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node33711 = (inp[1]) ? node33735 : node33712;
											assign node33712 = (inp[13]) ? node33724 : node33713;
												assign node33713 = (inp[11]) ? node33719 : node33714;
													assign node33714 = (inp[12]) ? 4'b0010 : node33715;
														assign node33715 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node33719 = (inp[4]) ? node33721 : 4'b0011;
														assign node33721 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node33724 = (inp[11]) ? node33730 : node33725;
													assign node33725 = (inp[12]) ? 4'b0011 : node33726;
														assign node33726 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node33730 = (inp[4]) ? node33732 : 4'b0010;
														assign node33732 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node33735 = (inp[11]) ? node33739 : node33736;
												assign node33736 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node33739 = (inp[13]) ? 4'b0010 : 4'b0011;
							assign node33742 = (inp[2]) ? node33960 : node33743;
								assign node33743 = (inp[11]) ? node33869 : node33744;
									assign node33744 = (inp[13]) ? node33816 : node33745;
										assign node33745 = (inp[12]) ? node33769 : node33746;
											assign node33746 = (inp[4]) ? node33760 : node33747;
												assign node33747 = (inp[10]) ? node33753 : node33748;
													assign node33748 = (inp[7]) ? 4'b0110 : node33749;
														assign node33749 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node33753 = (inp[5]) ? node33755 : 4'b0110;
														assign node33755 = (inp[7]) ? node33757 : 4'b0110;
															assign node33757 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node33760 = (inp[5]) ? node33764 : node33761;
													assign node33761 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node33764 = (inp[7]) ? 4'b0010 : node33765;
														assign node33765 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node33769 = (inp[0]) ? node33797 : node33770;
												assign node33770 = (inp[5]) ? node33782 : node33771;
													assign node33771 = (inp[7]) ? node33777 : node33772;
														assign node33772 = (inp[1]) ? node33774 : 4'b0010;
															assign node33774 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node33777 = (inp[4]) ? node33779 : 4'b0110;
															assign node33779 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node33782 = (inp[7]) ? node33792 : node33783;
														assign node33783 = (inp[10]) ? node33787 : node33784;
															assign node33784 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node33787 = (inp[1]) ? node33789 : 4'b0110;
																assign node33789 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node33792 = (inp[1]) ? 4'b0011 : node33793;
															assign node33793 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node33797 = (inp[4]) ? node33809 : node33798;
													assign node33798 = (inp[1]) ? node33802 : node33799;
														assign node33799 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node33802 = (inp[7]) ? node33806 : node33803;
															assign node33803 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node33806 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node33809 = (inp[1]) ? node33811 : 4'b0111;
														assign node33811 = (inp[5]) ? 4'b0110 : node33812;
															assign node33812 = (inp[7]) ? 4'b0110 : 4'b0010;
										assign node33816 = (inp[12]) ? node33842 : node33817;
											assign node33817 = (inp[1]) ? node33835 : node33818;
												assign node33818 = (inp[4]) ? node33828 : node33819;
													assign node33819 = (inp[10]) ? 4'b0111 : node33820;
														assign node33820 = (inp[7]) ? node33824 : node33821;
															assign node33821 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node33824 = (inp[5]) ? 4'b0010 : 4'b0111;
													assign node33828 = (inp[5]) ? node33832 : node33829;
														assign node33829 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node33832 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node33835 = (inp[7]) ? node33839 : node33836;
													assign node33836 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node33839 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node33842 = (inp[5]) ? node33854 : node33843;
												assign node33843 = (inp[7]) ? node33849 : node33844;
													assign node33844 = (inp[1]) ? node33846 : 4'b0011;
														assign node33846 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node33849 = (inp[1]) ? 4'b0111 : node33850;
														assign node33850 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node33854 = (inp[7]) ? node33862 : node33855;
													assign node33855 = (inp[10]) ? node33857 : 4'b0110;
														assign node33857 = (inp[4]) ? 4'b0110 : node33858;
															assign node33858 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node33862 = (inp[4]) ? node33866 : node33863;
														assign node33863 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node33866 = (inp[1]) ? 4'b0011 : 4'b0010;
									assign node33869 = (inp[13]) ? node33913 : node33870;
										assign node33870 = (inp[5]) ? node33886 : node33871;
											assign node33871 = (inp[7]) ? node33879 : node33872;
												assign node33872 = (inp[1]) ? node33874 : 4'b0011;
													assign node33874 = (inp[12]) ? node33876 : 4'b0011;
														assign node33876 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node33879 = (inp[12]) ? node33881 : 4'b0111;
													assign node33881 = (inp[4]) ? node33883 : 4'b0111;
														assign node33883 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node33886 = (inp[7]) ? node33900 : node33887;
												assign node33887 = (inp[4]) ? node33893 : node33888;
													assign node33888 = (inp[0]) ? node33890 : 4'b0111;
														assign node33890 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node33893 = (inp[12]) ? node33897 : node33894;
														assign node33894 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node33897 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node33900 = (inp[4]) ? node33908 : node33901;
													assign node33901 = (inp[12]) ? node33905 : node33902;
														assign node33902 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node33905 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node33908 = (inp[1]) ? 4'b0011 : node33909;
														assign node33909 = (inp[12]) ? 4'b0010 : 4'b0011;
										assign node33913 = (inp[7]) ? node33933 : node33914;
											assign node33914 = (inp[5]) ? node33920 : node33915;
												assign node33915 = (inp[1]) ? node33917 : 4'b0010;
													assign node33917 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node33920 = (inp[4]) ? node33926 : node33921;
													assign node33921 = (inp[1]) ? node33923 : 4'b0110;
														assign node33923 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node33926 = (inp[1]) ? node33930 : node33927;
														assign node33927 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node33930 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node33933 = (inp[5]) ? node33941 : node33934;
												assign node33934 = (inp[4]) ? node33936 : 4'b0110;
													assign node33936 = (inp[1]) ? 4'b0110 : node33937;
														assign node33937 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node33941 = (inp[4]) ? node33955 : node33942;
													assign node33942 = (inp[10]) ? node33950 : node33943;
														assign node33943 = (inp[12]) ? node33947 : node33944;
															assign node33944 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node33947 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node33950 = (inp[1]) ? 4'b0011 : node33951;
															assign node33951 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node33955 = (inp[1]) ? 4'b0010 : node33956;
														assign node33956 = (inp[12]) ? 4'b0011 : 4'b0010;
								assign node33960 = (inp[13]) ? node34052 : node33961;
									assign node33961 = (inp[11]) ? node34005 : node33962;
										assign node33962 = (inp[5]) ? node33990 : node33963;
											assign node33963 = (inp[7]) ? node33975 : node33964;
												assign node33964 = (inp[1]) ? node33968 : node33965;
													assign node33965 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node33968 = (inp[10]) ? node33970 : 4'b0011;
														assign node33970 = (inp[4]) ? 4'b0011 : node33971;
															assign node33971 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node33975 = (inp[1]) ? node33985 : node33976;
													assign node33976 = (inp[10]) ? 4'b0111 : node33977;
														assign node33977 = (inp[4]) ? node33981 : node33978;
															assign node33978 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node33981 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node33985 = (inp[12]) ? 4'b0110 : node33986;
														assign node33986 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node33990 = (inp[7]) ? node33998 : node33991;
												assign node33991 = (inp[1]) ? node33993 : 4'b0110;
													assign node33993 = (inp[4]) ? 4'b0110 : node33994;
														assign node33994 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node33998 = (inp[1]) ? 4'b0010 : node33999;
													assign node33999 = (inp[4]) ? node34001 : 4'b0010;
														assign node34001 = (inp[12]) ? 4'b0010 : 4'b0011;
										assign node34005 = (inp[12]) ? node34037 : node34006;
											assign node34006 = (inp[5]) ? node34026 : node34007;
												assign node34007 = (inp[7]) ? node34015 : node34008;
													assign node34008 = (inp[4]) ? node34012 : node34009;
														assign node34009 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node34012 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node34015 = (inp[10]) ? node34021 : node34016;
														assign node34016 = (inp[0]) ? 4'b0110 : node34017;
															assign node34017 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node34021 = (inp[1]) ? 4'b0111 : node34022;
															assign node34022 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node34026 = (inp[7]) ? node34032 : node34027;
													assign node34027 = (inp[4]) ? 4'b0111 : node34028;
														assign node34028 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node34032 = (inp[4]) ? node34034 : 4'b0011;
														assign node34034 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node34037 = (inp[5]) ? node34049 : node34038;
												assign node34038 = (inp[7]) ? node34044 : node34039;
													assign node34039 = (inp[4]) ? node34041 : 4'b0011;
														assign node34041 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node34044 = (inp[1]) ? 4'b0111 : node34045;
														assign node34045 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node34049 = (inp[7]) ? 4'b0011 : 4'b0111;
									assign node34052 = (inp[11]) ? node34098 : node34053;
										assign node34053 = (inp[12]) ? node34085 : node34054;
											assign node34054 = (inp[7]) ? node34072 : node34055;
												assign node34055 = (inp[5]) ? node34065 : node34056;
													assign node34056 = (inp[10]) ? 4'b0011 : node34057;
														assign node34057 = (inp[0]) ? node34059 : 4'b0011;
															assign node34059 = (inp[1]) ? 4'b0010 : node34060;
																assign node34060 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node34065 = (inp[10]) ? node34067 : 4'b0111;
														assign node34067 = (inp[4]) ? 4'b0111 : node34068;
															assign node34068 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node34072 = (inp[5]) ? node34080 : node34073;
													assign node34073 = (inp[4]) ? node34077 : node34074;
														assign node34074 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node34077 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node34080 = (inp[4]) ? node34082 : 4'b0011;
														assign node34082 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node34085 = (inp[5]) ? node34095 : node34086;
												assign node34086 = (inp[7]) ? node34092 : node34087;
													assign node34087 = (inp[4]) ? node34089 : 4'b0011;
														assign node34089 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node34092 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node34095 = (inp[7]) ? 4'b0011 : 4'b0111;
										assign node34098 = (inp[12]) ? node34124 : node34099;
											assign node34099 = (inp[4]) ? node34113 : node34100;
												assign node34100 = (inp[1]) ? node34108 : node34101;
													assign node34101 = (inp[7]) ? node34105 : node34102;
														assign node34102 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node34105 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node34108 = (inp[7]) ? 4'b0010 : node34109;
														assign node34109 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node34113 = (inp[1]) ? node34121 : node34114;
													assign node34114 = (inp[5]) ? node34118 : node34115;
														assign node34115 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node34118 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node34121 = (inp[7]) ? 4'b0110 : 4'b0010;
											assign node34124 = (inp[5]) ? node34136 : node34125;
												assign node34125 = (inp[7]) ? node34131 : node34126;
													assign node34126 = (inp[4]) ? node34128 : 4'b0010;
														assign node34128 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node34131 = (inp[1]) ? 4'b0110 : node34132;
														assign node34132 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node34136 = (inp[7]) ? 4'b0010 : 4'b0110;
						assign node34139 = (inp[7]) ? node34339 : node34140;
							assign node34140 = (inp[12]) ? node34254 : node34141;
								assign node34141 = (inp[4]) ? node34189 : node34142;
									assign node34142 = (inp[0]) ? node34166 : node34143;
										assign node34143 = (inp[13]) ? node34155 : node34144;
											assign node34144 = (inp[2]) ? node34150 : node34145;
												assign node34145 = (inp[5]) ? node34147 : 4'b0000;
													assign node34147 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node34150 = (inp[5]) ? node34152 : 4'b0001;
													assign node34152 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node34155 = (inp[2]) ? node34161 : node34156;
												assign node34156 = (inp[1]) ? node34158 : 4'b0001;
													assign node34158 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node34161 = (inp[1]) ? node34163 : 4'b0000;
													assign node34163 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node34166 = (inp[2]) ? node34178 : node34167;
											assign node34167 = (inp[13]) ? node34173 : node34168;
												assign node34168 = (inp[1]) ? node34170 : 4'b0000;
													assign node34170 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node34173 = (inp[5]) ? node34175 : 4'b0001;
													assign node34175 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node34178 = (inp[13]) ? node34184 : node34179;
												assign node34179 = (inp[5]) ? node34181 : 4'b0001;
													assign node34181 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node34184 = (inp[1]) ? node34186 : 4'b0000;
													assign node34186 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node34189 = (inp[0]) ? node34247 : node34190;
										assign node34190 = (inp[11]) ? node34220 : node34191;
											assign node34191 = (inp[9]) ? node34205 : node34192;
												assign node34192 = (inp[10]) ? node34200 : node34193;
													assign node34193 = (inp[13]) ? node34197 : node34194;
														assign node34194 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node34197 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node34200 = (inp[13]) ? node34202 : 4'b0101;
														assign node34202 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node34205 = (inp[10]) ? node34215 : node34206;
													assign node34206 = (inp[2]) ? 4'b0101 : node34207;
														assign node34207 = (inp[13]) ? node34211 : node34208;
															assign node34208 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node34211 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node34215 = (inp[5]) ? node34217 : 4'b0100;
														assign node34217 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node34220 = (inp[2]) ? node34242 : node34221;
												assign node34221 = (inp[1]) ? node34231 : node34222;
													assign node34222 = (inp[9]) ? node34224 : 4'b0100;
														assign node34224 = (inp[5]) ? node34228 : node34225;
															assign node34225 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node34228 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node34231 = (inp[9]) ? node34237 : node34232;
														assign node34232 = (inp[5]) ? 4'b0101 : node34233;
															assign node34233 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node34237 = (inp[13]) ? 4'b0100 : node34238;
															assign node34238 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node34242 = (inp[1]) ? 4'b0100 : node34243;
													assign node34243 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node34247 = (inp[13]) ? node34251 : node34248;
											assign node34248 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node34251 = (inp[5]) ? 4'b0100 : 4'b0101;
								assign node34254 = (inp[10]) ? node34304 : node34255;
									assign node34255 = (inp[5]) ? node34293 : node34256;
										assign node34256 = (inp[13]) ? node34278 : node34257;
											assign node34257 = (inp[4]) ? 4'b0100 : node34258;
												assign node34258 = (inp[0]) ? node34264 : node34259;
													assign node34259 = (inp[2]) ? 4'b0101 : node34260;
														assign node34260 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node34264 = (inp[9]) ? node34270 : node34265;
														assign node34265 = (inp[2]) ? node34267 : 4'b0100;
															assign node34267 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node34270 = (inp[1]) ? node34274 : node34271;
															assign node34271 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node34274 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node34278 = (inp[4]) ? 4'b0101 : node34279;
												assign node34279 = (inp[9]) ? node34281 : 4'b0100;
													assign node34281 = (inp[11]) ? node34287 : node34282;
														assign node34282 = (inp[2]) ? node34284 : 4'b0101;
															assign node34284 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node34287 = (inp[1]) ? node34289 : 4'b0100;
															assign node34289 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node34293 = (inp[13]) ? node34299 : node34294;
											assign node34294 = (inp[4]) ? 4'b0101 : node34295;
												assign node34295 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node34299 = (inp[2]) ? 4'b0100 : node34300;
												assign node34300 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node34304 = (inp[2]) ? node34324 : node34305;
										assign node34305 = (inp[13]) ? node34315 : node34306;
											assign node34306 = (inp[5]) ? node34312 : node34307;
												assign node34307 = (inp[1]) ? node34309 : 4'b0100;
													assign node34309 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node34312 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node34315 = (inp[4]) ? node34321 : node34316;
												assign node34316 = (inp[5]) ? 4'b0101 : node34317;
													assign node34317 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node34321 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node34324 = (inp[13]) ? node34332 : node34325;
											assign node34325 = (inp[5]) ? 4'b0101 : node34326;
												assign node34326 = (inp[1]) ? 4'b0100 : node34327;
													assign node34327 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node34332 = (inp[5]) ? 4'b0100 : node34333;
												assign node34333 = (inp[1]) ? 4'b0101 : node34334;
													assign node34334 = (inp[4]) ? 4'b0101 : 4'b0100;
							assign node34339 = (inp[12]) ? node34433 : node34340;
								assign node34340 = (inp[4]) ? node34364 : node34341;
									assign node34341 = (inp[13]) ? node34353 : node34342;
										assign node34342 = (inp[2]) ? node34348 : node34343;
											assign node34343 = (inp[1]) ? 4'b0100 : node34344;
												assign node34344 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node34348 = (inp[1]) ? 4'b0101 : node34349;
												assign node34349 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node34353 = (inp[2]) ? node34359 : node34354;
											assign node34354 = (inp[1]) ? 4'b0101 : node34355;
												assign node34355 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node34359 = (inp[5]) ? node34361 : 4'b0100;
												assign node34361 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node34364 = (inp[0]) ? node34418 : node34365;
										assign node34365 = (inp[9]) ? node34391 : node34366;
											assign node34366 = (inp[11]) ? node34380 : node34367;
												assign node34367 = (inp[2]) ? node34373 : node34368;
													assign node34368 = (inp[1]) ? node34370 : 4'b0000;
														assign node34370 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node34373 = (inp[1]) ? node34377 : node34374;
														assign node34374 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node34377 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node34380 = (inp[10]) ? node34386 : node34381;
													assign node34381 = (inp[13]) ? 4'b0000 : node34382;
														assign node34382 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node34386 = (inp[13]) ? 4'b0001 : node34387;
														assign node34387 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node34391 = (inp[2]) ? node34405 : node34392;
												assign node34392 = (inp[10]) ? node34400 : node34393;
													assign node34393 = (inp[13]) ? node34397 : node34394;
														assign node34394 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node34397 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node34400 = (inp[5]) ? node34402 : 4'b0000;
														assign node34402 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node34405 = (inp[5]) ? node34411 : node34406;
													assign node34406 = (inp[13]) ? 4'b0001 : node34407;
														assign node34407 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node34411 = (inp[1]) ? node34415 : node34412;
														assign node34412 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node34415 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node34418 = (inp[5]) ? node34426 : node34419;
											assign node34419 = (inp[1]) ? node34423 : node34420;
												assign node34420 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node34423 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node34426 = (inp[13]) ? node34430 : node34427;
												assign node34427 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node34430 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node34433 = (inp[13]) ? node34447 : node34434;
									assign node34434 = (inp[4]) ? 4'b0001 : node34435;
										assign node34435 = (inp[2]) ? node34441 : node34436;
											assign node34436 = (inp[5]) ? 4'b0000 : node34437;
												assign node34437 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node34441 = (inp[5]) ? 4'b0001 : node34442;
												assign node34442 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node34447 = (inp[4]) ? 4'b0000 : node34448;
										assign node34448 = (inp[2]) ? node34454 : node34449;
											assign node34449 = (inp[5]) ? 4'b0001 : node34450;
												assign node34450 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node34454 = (inp[1]) ? 4'b0000 : node34455;
												assign node34455 = (inp[5]) ? 4'b0000 : 4'b0001;
					assign node34460 = (inp[5]) ? node34972 : node34461;
						assign node34461 = (inp[14]) ? node34853 : node34462;
							assign node34462 = (inp[4]) ? node34732 : node34463;
								assign node34463 = (inp[12]) ? node34613 : node34464;
									assign node34464 = (inp[0]) ? node34548 : node34465;
										assign node34465 = (inp[2]) ? node34499 : node34466;
											assign node34466 = (inp[7]) ? node34488 : node34467;
												assign node34467 = (inp[13]) ? node34481 : node34468;
													assign node34468 = (inp[9]) ? node34470 : 4'b0000;
														assign node34470 = (inp[10]) ? node34476 : node34471;
															assign node34471 = (inp[11]) ? 4'b0000 : node34472;
																assign node34472 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node34476 = (inp[11]) ? node34478 : 4'b0000;
																assign node34478 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node34481 = (inp[11]) ? node34485 : node34482;
														assign node34482 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node34485 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node34488 = (inp[13]) ? node34494 : node34489;
													assign node34489 = (inp[1]) ? 4'b0000 : node34490;
														assign node34490 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node34494 = (inp[1]) ? node34496 : 4'b0000;
														assign node34496 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node34499 = (inp[10]) ? node34533 : node34500;
												assign node34500 = (inp[9]) ? node34518 : node34501;
													assign node34501 = (inp[7]) ? node34511 : node34502;
														assign node34502 = (inp[13]) ? node34504 : 4'b0001;
															assign node34504 = (inp[11]) ? node34508 : node34505;
																assign node34505 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node34508 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node34511 = (inp[13]) ? 4'b0001 : node34512;
															assign node34512 = (inp[1]) ? node34514 : 4'b0000;
																assign node34514 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node34518 = (inp[7]) ? node34526 : node34519;
														assign node34519 = (inp[1]) ? node34523 : node34520;
															assign node34520 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node34523 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node34526 = (inp[1]) ? node34530 : node34527;
															assign node34527 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node34530 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node34533 = (inp[1]) ? node34541 : node34534;
													assign node34534 = (inp[13]) ? 4'b0000 : node34535;
														assign node34535 = (inp[7]) ? node34537 : 4'b0000;
															assign node34537 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node34541 = (inp[11]) ? node34545 : node34542;
														assign node34542 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node34545 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node34548 = (inp[2]) ? node34574 : node34549;
											assign node34549 = (inp[10]) ? node34567 : node34550;
												assign node34550 = (inp[7]) ? 4'b0001 : node34551;
													assign node34551 = (inp[9]) ? node34561 : node34552;
														assign node34552 = (inp[13]) ? node34554 : 4'b0000;
															assign node34554 = (inp[1]) ? node34558 : node34555;
																assign node34555 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node34558 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node34561 = (inp[1]) ? node34563 : 4'b0001;
															assign node34563 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node34567 = (inp[1]) ? node34571 : node34568;
													assign node34568 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node34571 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node34574 = (inp[10]) ? node34600 : node34575;
												assign node34575 = (inp[13]) ? node34589 : node34576;
													assign node34576 = (inp[1]) ? node34584 : node34577;
														assign node34577 = (inp[11]) ? node34581 : node34578;
															assign node34578 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node34581 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node34584 = (inp[11]) ? 4'b0000 : node34585;
															assign node34585 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node34589 = (inp[9]) ? node34591 : 4'b0000;
														assign node34591 = (inp[7]) ? node34593 : 4'b0000;
															assign node34593 = (inp[1]) ? node34597 : node34594;
																assign node34594 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node34597 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node34600 = (inp[1]) ? node34608 : node34601;
													assign node34601 = (inp[11]) ? node34605 : node34602;
														assign node34602 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node34605 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node34608 = (inp[13]) ? 4'b0001 : node34609;
														assign node34609 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node34613 = (inp[10]) ? node34661 : node34614;
										assign node34614 = (inp[1]) ? node34638 : node34615;
											assign node34615 = (inp[13]) ? node34623 : node34616;
												assign node34616 = (inp[7]) ? node34620 : node34617;
													assign node34617 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node34620 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node34623 = (inp[2]) ? node34625 : 4'b0101;
													assign node34625 = (inp[9]) ? node34633 : node34626;
														assign node34626 = (inp[11]) ? node34630 : node34627;
															assign node34627 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node34630 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node34633 = (inp[11]) ? 4'b0101 : node34634;
															assign node34634 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node34638 = (inp[2]) ? node34654 : node34639;
												assign node34639 = (inp[0]) ? node34647 : node34640;
													assign node34640 = (inp[7]) ? node34644 : node34641;
														assign node34641 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node34644 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node34647 = (inp[11]) ? node34651 : node34648;
														assign node34648 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node34651 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node34654 = (inp[11]) ? node34658 : node34655;
													assign node34655 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node34658 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node34661 = (inp[1]) ? node34703 : node34662;
											assign node34662 = (inp[9]) ? node34690 : node34663;
												assign node34663 = (inp[13]) ? node34675 : node34664;
													assign node34664 = (inp[2]) ? node34666 : 4'b0101;
														assign node34666 = (inp[0]) ? node34672 : node34667;
															assign node34667 = (inp[11]) ? node34669 : 4'b0101;
																assign node34669 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node34672 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node34675 = (inp[0]) ? node34681 : node34676;
														assign node34676 = (inp[11]) ? 4'b0100 : node34677;
															assign node34677 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node34681 = (inp[2]) ? node34683 : 4'b0101;
															assign node34683 = (inp[7]) ? node34687 : node34684;
																assign node34684 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node34687 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node34690 = (inp[0]) ? node34696 : node34691;
													assign node34691 = (inp[11]) ? 4'b0100 : node34692;
														assign node34692 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node34696 = (inp[11]) ? node34700 : node34697;
														assign node34697 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node34700 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node34703 = (inp[9]) ? node34711 : node34704;
												assign node34704 = (inp[7]) ? node34708 : node34705;
													assign node34705 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node34708 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node34711 = (inp[2]) ? node34719 : node34712;
													assign node34712 = (inp[13]) ? node34714 : 4'b0100;
														assign node34714 = (inp[7]) ? node34716 : 4'b0101;
															assign node34716 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node34719 = (inp[0]) ? node34721 : 4'b0101;
														assign node34721 = (inp[13]) ? node34727 : node34722;
															assign node34722 = (inp[7]) ? 4'b0101 : node34723;
																assign node34723 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node34727 = (inp[7]) ? node34729 : 4'b0101;
																assign node34729 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node34732 = (inp[9]) ? node34800 : node34733;
									assign node34733 = (inp[11]) ? node34765 : node34734;
										assign node34734 = (inp[7]) ? node34760 : node34735;
											assign node34735 = (inp[12]) ? 4'b0100 : node34736;
												assign node34736 = (inp[13]) ? node34744 : node34737;
													assign node34737 = (inp[2]) ? node34741 : node34738;
														assign node34738 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node34741 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node34744 = (inp[10]) ? node34750 : node34745;
														assign node34745 = (inp[2]) ? 4'b0100 : node34746;
															assign node34746 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node34750 = (inp[0]) ? 4'b0101 : node34751;
															assign node34751 = (inp[1]) ? node34755 : node34752;
																assign node34752 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node34755 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node34760 = (inp[12]) ? 4'b0101 : node34761;
												assign node34761 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node34765 = (inp[7]) ? node34795 : node34766;
											assign node34766 = (inp[12]) ? 4'b0101 : node34767;
												assign node34767 = (inp[10]) ? node34775 : node34768;
													assign node34768 = (inp[2]) ? node34772 : node34769;
														assign node34769 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node34772 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node34775 = (inp[0]) ? node34787 : node34776;
														assign node34776 = (inp[13]) ? node34782 : node34777;
															assign node34777 = (inp[1]) ? 4'b0101 : node34778;
																assign node34778 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node34782 = (inp[1]) ? node34784 : 4'b0101;
																assign node34784 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node34787 = (inp[1]) ? node34791 : node34788;
															assign node34788 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node34791 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node34795 = (inp[1]) ? 4'b0100 : node34796;
												assign node34796 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node34800 = (inp[1]) ? node34838 : node34801;
										assign node34801 = (inp[12]) ? node34813 : node34802;
											assign node34802 = (inp[11]) ? node34808 : node34803;
												assign node34803 = (inp[7]) ? 4'b0100 : node34804;
													assign node34804 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node34808 = (inp[7]) ? 4'b0101 : node34809;
													assign node34809 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node34813 = (inp[13]) ? node34823 : node34814;
												assign node34814 = (inp[2]) ? 4'b0101 : node34815;
													assign node34815 = (inp[11]) ? node34819 : node34816;
														assign node34816 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node34819 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node34823 = (inp[2]) ? node34831 : node34824;
													assign node34824 = (inp[11]) ? node34828 : node34825;
														assign node34825 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node34828 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node34831 = (inp[7]) ? node34835 : node34832;
														assign node34832 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node34835 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node34838 = (inp[11]) ? node34846 : node34839;
											assign node34839 = (inp[7]) ? 4'b0101 : node34840;
												assign node34840 = (inp[2]) ? 4'b0100 : node34841;
													assign node34841 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node34846 = (inp[7]) ? 4'b0100 : node34847;
												assign node34847 = (inp[2]) ? 4'b0101 : node34848;
													assign node34848 = (inp[12]) ? 4'b0101 : 4'b0100;
							assign node34853 = (inp[4]) ? node34961 : node34854;
								assign node34854 = (inp[12]) ? node34870 : node34855;
									assign node34855 = (inp[0]) ? node34863 : node34856;
										assign node34856 = (inp[2]) ? node34860 : node34857;
											assign node34857 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node34860 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node34863 = (inp[2]) ? node34867 : node34864;
											assign node34864 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node34867 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node34870 = (inp[1]) ? node34932 : node34871;
										assign node34871 = (inp[10]) ? node34899 : node34872;
											assign node34872 = (inp[0]) ? node34886 : node34873;
												assign node34873 = (inp[13]) ? node34879 : node34874;
													assign node34874 = (inp[7]) ? 4'b0001 : node34875;
														assign node34875 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node34879 = (inp[2]) ? node34883 : node34880;
														assign node34880 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node34883 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node34886 = (inp[13]) ? 4'b0001 : node34887;
													assign node34887 = (inp[11]) ? node34893 : node34888;
														assign node34888 = (inp[7]) ? node34890 : 4'b0000;
															assign node34890 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node34893 = (inp[7]) ? node34895 : 4'b0001;
															assign node34895 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node34899 = (inp[0]) ? node34915 : node34900;
												assign node34900 = (inp[11]) ? node34908 : node34901;
													assign node34901 = (inp[7]) ? node34905 : node34902;
														assign node34902 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node34905 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node34908 = (inp[13]) ? node34910 : 4'b0001;
														assign node34910 = (inp[7]) ? node34912 : 4'b0001;
															assign node34912 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node34915 = (inp[11]) ? node34927 : node34916;
													assign node34916 = (inp[9]) ? node34922 : node34917;
														assign node34917 = (inp[2]) ? 4'b0001 : node34918;
															assign node34918 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node34922 = (inp[7]) ? node34924 : 4'b0001;
															assign node34924 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node34927 = (inp[7]) ? node34929 : 4'b0000;
														assign node34929 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node34932 = (inp[11]) ? node34954 : node34933;
											assign node34933 = (inp[10]) ? node34941 : node34934;
												assign node34934 = (inp[2]) ? node34938 : node34935;
													assign node34935 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node34938 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node34941 = (inp[0]) ? node34947 : node34942;
													assign node34942 = (inp[13]) ? node34944 : 4'b0001;
														assign node34944 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node34947 = (inp[2]) ? node34951 : node34948;
														assign node34948 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node34951 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node34954 = (inp[7]) ? node34958 : node34955;
												assign node34955 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node34958 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node34961 = (inp[7]) ? node34967 : node34962;
									assign node34962 = (inp[1]) ? 4'b0001 : node34963;
										assign node34963 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node34967 = (inp[1]) ? 4'b0000 : node34968;
										assign node34968 = (inp[12]) ? 4'b0000 : 4'b0001;
						assign node34972 = (inp[12]) ? node35146 : node34973;
							assign node34973 = (inp[4]) ? node35119 : node34974;
								assign node34974 = (inp[14]) ? node35076 : node34975;
									assign node34975 = (inp[9]) ? node34999 : node34976;
										assign node34976 = (inp[1]) ? node34988 : node34977;
											assign node34977 = (inp[11]) ? node34983 : node34978;
												assign node34978 = (inp[2]) ? 4'b0100 : node34979;
													assign node34979 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node34983 = (inp[7]) ? node34985 : 4'b0101;
													assign node34985 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node34988 = (inp[11]) ? node34994 : node34989;
												assign node34989 = (inp[2]) ? 4'b0101 : node34990;
													assign node34990 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node34994 = (inp[2]) ? 4'b0100 : node34995;
													assign node34995 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node34999 = (inp[7]) ? node35035 : node35000;
											assign node35000 = (inp[13]) ? node35014 : node35001;
												assign node35001 = (inp[2]) ? node35009 : node35002;
													assign node35002 = (inp[1]) ? node35006 : node35003;
														assign node35003 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node35006 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node35009 = (inp[1]) ? node35011 : 4'b0101;
														assign node35011 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node35014 = (inp[0]) ? node35028 : node35015;
													assign node35015 = (inp[2]) ? node35021 : node35016;
														assign node35016 = (inp[11]) ? node35018 : 4'b0101;
															assign node35018 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node35021 = (inp[11]) ? node35025 : node35022;
															assign node35022 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node35025 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node35028 = (inp[11]) ? node35032 : node35029;
														assign node35029 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node35032 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node35035 = (inp[0]) ? node35061 : node35036;
												assign node35036 = (inp[10]) ? node35050 : node35037;
													assign node35037 = (inp[11]) ? 4'b0100 : node35038;
														assign node35038 = (inp[13]) ? node35044 : node35039;
															assign node35039 = (inp[2]) ? 4'b0100 : node35040;
																assign node35040 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node35044 = (inp[1]) ? node35046 : 4'b0100;
																assign node35046 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node35050 = (inp[2]) ? node35052 : 4'b0101;
														assign node35052 = (inp[13]) ? 4'b0100 : node35053;
															assign node35053 = (inp[1]) ? node35057 : node35054;
																assign node35054 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node35057 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node35061 = (inp[10]) ? node35071 : node35062;
													assign node35062 = (inp[2]) ? 4'b0101 : node35063;
														assign node35063 = (inp[1]) ? node35067 : node35064;
															assign node35064 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node35067 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node35071 = (inp[11]) ? node35073 : 4'b0100;
														assign node35073 = (inp[1]) ? 4'b0101 : 4'b0100;
									assign node35076 = (inp[11]) ? node35104 : node35077;
										assign node35077 = (inp[7]) ? node35097 : node35078;
											assign node35078 = (inp[9]) ? node35086 : node35079;
												assign node35079 = (inp[1]) ? node35083 : node35080;
													assign node35080 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node35083 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node35086 = (inp[13]) ? node35092 : node35087;
													assign node35087 = (inp[1]) ? node35089 : 4'b0101;
														assign node35089 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node35092 = (inp[1]) ? 4'b0101 : node35093;
														assign node35093 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node35097 = (inp[1]) ? node35101 : node35098;
												assign node35098 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node35101 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node35104 = (inp[9]) ? node35112 : node35105;
											assign node35105 = (inp[1]) ? node35109 : node35106;
												assign node35106 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node35109 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node35112 = (inp[1]) ? node35116 : node35113;
												assign node35113 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node35116 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node35119 = (inp[1]) ? node35133 : node35120;
									assign node35120 = (inp[14]) ? 4'b0001 : node35121;
										assign node35121 = (inp[11]) ? node35127 : node35122;
											assign node35122 = (inp[2]) ? 4'b0000 : node35123;
												assign node35123 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node35127 = (inp[7]) ? 4'b0001 : node35128;
												assign node35128 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node35133 = (inp[14]) ? 4'b0000 : node35134;
										assign node35134 = (inp[11]) ? node35140 : node35135;
											assign node35135 = (inp[7]) ? 4'b0001 : node35136;
												assign node35136 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node35140 = (inp[2]) ? 4'b0000 : node35141;
												assign node35141 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node35146 = (inp[14]) ? node35158 : node35147;
								assign node35147 = (inp[11]) ? node35153 : node35148;
									assign node35148 = (inp[4]) ? 4'b0001 : node35149;
										assign node35149 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node35153 = (inp[4]) ? 4'b0000 : node35154;
										assign node35154 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node35158 = (inp[2]) ? 4'b0000 : node35159;
									assign node35159 = (inp[4]) ? 4'b0000 : 4'b0001;

endmodule