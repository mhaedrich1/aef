module dtc_split875_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node17;
	wire [8-1:0] node20;
	wire [8-1:0] node22;
	wire [8-1:0] node23;
	wire [8-1:0] node26;
	wire [8-1:0] node29;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node33;
	wire [8-1:0] node36;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node42;
	wire [8-1:0] node45;
	wire [8-1:0] node46;
	wire [8-1:0] node49;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node52;
	wire [8-1:0] node56;
	wire [8-1:0] node58;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node63;
	wire [8-1:0] node67;
	wire [8-1:0] node68;
	wire [8-1:0] node72;
	wire [8-1:0] node73;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node77;
	wire [8-1:0] node80;
	wire [8-1:0] node81;
	wire [8-1:0] node83;
	wire [8-1:0] node86;
	wire [8-1:0] node88;
	wire [8-1:0] node91;
	wire [8-1:0] node92;
	wire [8-1:0] node93;
	wire [8-1:0] node95;
	wire [8-1:0] node98;
	wire [8-1:0] node99;
	wire [8-1:0] node101;
	wire [8-1:0] node104;
	wire [8-1:0] node106;
	wire [8-1:0] node109;
	wire [8-1:0] node110;
	wire [8-1:0] node112;
	wire [8-1:0] node115;
	wire [8-1:0] node116;
	wire [8-1:0] node118;
	wire [8-1:0] node121;
	wire [8-1:0] node123;
	wire [8-1:0] node127;
	wire [8-1:0] node128;
	wire [8-1:0] node129;
	wire [8-1:0] node130;
	wire [8-1:0] node133;
	wire [8-1:0] node134;
	wire [8-1:0] node135;
	wire [8-1:0] node137;
	wire [8-1:0] node140;
	wire [8-1:0] node141;
	wire [8-1:0] node145;
	wire [8-1:0] node146;
	wire [8-1:0] node148;
	wire [8-1:0] node151;
	wire [8-1:0] node152;
	wire [8-1:0] node156;
	wire [8-1:0] node157;
	wire [8-1:0] node158;
	wire [8-1:0] node159;
	wire [8-1:0] node161;
	wire [8-1:0] node164;
	wire [8-1:0] node166;
	wire [8-1:0] node169;
	wire [8-1:0] node170;
	wire [8-1:0] node172;
	wire [8-1:0] node173;
	wire [8-1:0] node176;
	wire [8-1:0] node179;
	wire [8-1:0] node180;
	wire [8-1:0] node181;
	wire [8-1:0] node184;
	wire [8-1:0] node188;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node191;
	wire [8-1:0] node195;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node206;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node212;
	wire [8-1:0] node215;
	wire [8-1:0] node219;
	wire [8-1:0] node220;
	wire [8-1:0] node221;
	wire [8-1:0] node222;
	wire [8-1:0] node223;
	wire [8-1:0] node225;
	wire [8-1:0] node228;
	wire [8-1:0] node230;
	wire [8-1:0] node231;
	wire [8-1:0] node234;
	wire [8-1:0] node237;
	wire [8-1:0] node238;
	wire [8-1:0] node239;
	wire [8-1:0] node243;
	wire [8-1:0] node244;
	wire [8-1:0] node245;
	wire [8-1:0] node248;
	wire [8-1:0] node252;
	wire [8-1:0] node253;
	wire [8-1:0] node254;
	wire [8-1:0] node256;
	wire [8-1:0] node257;
	wire [8-1:0] node260;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node268;
	wire [8-1:0] node272;
	wire [8-1:0] node273;
	wire [8-1:0] node275;
	wire [8-1:0] node276;
	wire [8-1:0] node277;
	wire [8-1:0] node280;
	wire [8-1:0] node283;
	wire [8-1:0] node284;
	wire [8-1:0] node287;
	wire [8-1:0] node290;
	wire [8-1:0] node291;
	wire [8-1:0] node292;
	wire [8-1:0] node293;
	wire [8-1:0] node296;
	wire [8-1:0] node299;
	wire [8-1:0] node300;
	wire [8-1:0] node303;
	wire [8-1:0] node307;
	wire [8-1:0] node308;
	wire [8-1:0] node309;
	wire [8-1:0] node310;
	wire [8-1:0] node313;
	wire [8-1:0] node314;
	wire [8-1:0] node316;
	wire [8-1:0] node319;
	wire [8-1:0] node320;
	wire [8-1:0] node323;
	wire [8-1:0] node326;
	wire [8-1:0] node327;
	wire [8-1:0] node328;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node337;
	wire [8-1:0] node341;
	wire [8-1:0] node342;
	wire [8-1:0] node343;
	wire [8-1:0] node346;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node351;
	wire [8-1:0] node352;
	wire [8-1:0] node355;
	wire [8-1:0] node358;
	wire [8-1:0] node359;
	wire [8-1:0] node361;
	wire [8-1:0] node364;
	wire [8-1:0] node366;
	wire [8-1:0] node369;
	wire [8-1:0] node370;
	wire [8-1:0] node371;
	wire [8-1:0] node372;
	wire [8-1:0] node374;
	wire [8-1:0] node377;
	wire [8-1:0] node378;
	wire [8-1:0] node381;
	wire [8-1:0] node384;
	wire [8-1:0] node385;
	wire [8-1:0] node388;
	wire [8-1:0] node389;
	wire [8-1:0] node392;
	wire [8-1:0] node395;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node400;
	wire [8-1:0] node401;
	wire [8-1:0] node402;
	wire [8-1:0] node403;
	wire [8-1:0] node404;
	wire [8-1:0] node405;
	wire [8-1:0] node406;
	wire [8-1:0] node410;
	wire [8-1:0] node411;
	wire [8-1:0] node415;
	wire [8-1:0] node416;
	wire [8-1:0] node417;
	wire [8-1:0] node418;
	wire [8-1:0] node421;
	wire [8-1:0] node422;
	wire [8-1:0] node426;
	wire [8-1:0] node427;
	wire [8-1:0] node431;
	wire [8-1:0] node432;
	wire [8-1:0] node433;
	wire [8-1:0] node436;
	wire [8-1:0] node438;
	wire [8-1:0] node441;
	wire [8-1:0] node443;
	wire [8-1:0] node446;
	wire [8-1:0] node447;
	wire [8-1:0] node448;
	wire [8-1:0] node450;
	wire [8-1:0] node453;
	wire [8-1:0] node454;
	wire [8-1:0] node458;
	wire [8-1:0] node459;
	wire [8-1:0] node460;
	wire [8-1:0] node463;
	wire [8-1:0] node466;
	wire [8-1:0] node467;
	wire [8-1:0] node468;
	wire [8-1:0] node471;
	wire [8-1:0] node472;
	wire [8-1:0] node476;
	wire [8-1:0] node477;
	wire [8-1:0] node478;
	wire [8-1:0] node483;
	wire [8-1:0] node484;
	wire [8-1:0] node485;
	wire [8-1:0] node486;
	wire [8-1:0] node487;
	wire [8-1:0] node490;
	wire [8-1:0] node491;
	wire [8-1:0] node494;
	wire [8-1:0] node495;
	wire [8-1:0] node499;
	wire [8-1:0] node500;
	wire [8-1:0] node502;
	wire [8-1:0] node505;
	wire [8-1:0] node508;
	wire [8-1:0] node509;
	wire [8-1:0] node510;
	wire [8-1:0] node511;
	wire [8-1:0] node515;
	wire [8-1:0] node518;
	wire [8-1:0] node519;
	wire [8-1:0] node520;
	wire [8-1:0] node524;
	wire [8-1:0] node525;
	wire [8-1:0] node529;
	wire [8-1:0] node530;
	wire [8-1:0] node531;
	wire [8-1:0] node532;
	wire [8-1:0] node534;
	wire [8-1:0] node537;
	wire [8-1:0] node539;
	wire [8-1:0] node541;
	wire [8-1:0] node544;
	wire [8-1:0] node545;
	wire [8-1:0] node546;
	wire [8-1:0] node550;
	wire [8-1:0] node551;
	wire [8-1:0] node554;
	wire [8-1:0] node556;
	wire [8-1:0] node559;
	wire [8-1:0] node560;
	wire [8-1:0] node561;
	wire [8-1:0] node562;
	wire [8-1:0] node565;
	wire [8-1:0] node567;
	wire [8-1:0] node570;
	wire [8-1:0] node571;
	wire [8-1:0] node573;
	wire [8-1:0] node576;
	wire [8-1:0] node578;
	wire [8-1:0] node581;
	wire [8-1:0] node582;
	wire [8-1:0] node583;
	wire [8-1:0] node584;
	wire [8-1:0] node587;
	wire [8-1:0] node590;
	wire [8-1:0] node591;
	wire [8-1:0] node594;
	wire [8-1:0] node597;
	wire [8-1:0] node600;
	wire [8-1:0] node601;
	wire [8-1:0] node602;
	wire [8-1:0] node603;
	wire [8-1:0] node605;
	wire [8-1:0] node606;
	wire [8-1:0] node610;
	wire [8-1:0] node611;
	wire [8-1:0] node612;
	wire [8-1:0] node613;
	wire [8-1:0] node614;
	wire [8-1:0] node618;
	wire [8-1:0] node620;
	wire [8-1:0] node623;
	wire [8-1:0] node624;
	wire [8-1:0] node628;
	wire [8-1:0] node629;
	wire [8-1:0] node630;
	wire [8-1:0] node631;
	wire [8-1:0] node634;
	wire [8-1:0] node637;
	wire [8-1:0] node638;
	wire [8-1:0] node641;
	wire [8-1:0] node644;
	wire [8-1:0] node645;
	wire [8-1:0] node649;
	wire [8-1:0] node650;
	wire [8-1:0] node651;
	wire [8-1:0] node652;
	wire [8-1:0] node655;
	wire [8-1:0] node657;
	wire [8-1:0] node660;
	wire [8-1:0] node662;
	wire [8-1:0] node663;
	wire [8-1:0] node666;
	wire [8-1:0] node669;
	wire [8-1:0] node670;
	wire [8-1:0] node672;
	wire [8-1:0] node676;
	wire [8-1:0] node677;
	wire [8-1:0] node678;
	wire [8-1:0] node679;
	wire [8-1:0] node680;
	wire [8-1:0] node683;
	wire [8-1:0] node686;
	wire [8-1:0] node687;
	wire [8-1:0] node688;
	wire [8-1:0] node690;
	wire [8-1:0] node693;
	wire [8-1:0] node694;
	wire [8-1:0] node698;
	wire [8-1:0] node699;
	wire [8-1:0] node701;
	wire [8-1:0] node704;
	wire [8-1:0] node705;
	wire [8-1:0] node709;
	wire [8-1:0] node710;
	wire [8-1:0] node711;
	wire [8-1:0] node713;
	wire [8-1:0] node716;
	wire [8-1:0] node718;
	wire [8-1:0] node721;
	wire [8-1:0] node722;
	wire [8-1:0] node724;
	wire [8-1:0] node727;
	wire [8-1:0] node730;
	wire [8-1:0] node731;
	wire [8-1:0] node732;
	wire [8-1:0] node733;
	wire [8-1:0] node735;
	wire [8-1:0] node736;
	wire [8-1:0] node739;
	wire [8-1:0] node742;
	wire [8-1:0] node743;
	wire [8-1:0] node745;
	wire [8-1:0] node748;
	wire [8-1:0] node751;
	wire [8-1:0] node752;
	wire [8-1:0] node754;
	wire [8-1:0] node757;
	wire [8-1:0] node758;
	wire [8-1:0] node759;
	wire [8-1:0] node762;
	wire [8-1:0] node765;
	wire [8-1:0] node766;
	wire [8-1:0] node769;
	wire [8-1:0] node772;
	wire [8-1:0] node773;
	wire [8-1:0] node774;
	wire [8-1:0] node775;
	wire [8-1:0] node777;
	wire [8-1:0] node780;
	wire [8-1:0] node781;
	wire [8-1:0] node784;
	wire [8-1:0] node787;
	wire [8-1:0] node788;
	wire [8-1:0] node791;
	wire [8-1:0] node794;
	wire [8-1:0] node795;
	wire [8-1:0] node796;
	wire [8-1:0] node797;
	wire [8-1:0] node801;
	wire [8-1:0] node802;
	wire [8-1:0] node805;
	wire [8-1:0] node808;
	wire [8-1:0] node811;
	wire [8-1:0] node812;
	wire [8-1:0] node813;
	wire [8-1:0] node814;
	wire [8-1:0] node815;
	wire [8-1:0] node816;
	wire [8-1:0] node817;
	wire [8-1:0] node819;
	wire [8-1:0] node822;
	wire [8-1:0] node824;
	wire [8-1:0] node827;
	wire [8-1:0] node828;
	wire [8-1:0] node832;
	wire [8-1:0] node833;
	wire [8-1:0] node834;
	wire [8-1:0] node838;
	wire [8-1:0] node839;
	wire [8-1:0] node841;
	wire [8-1:0] node844;
	wire [8-1:0] node845;
	wire [8-1:0] node849;
	wire [8-1:0] node850;
	wire [8-1:0] node851;
	wire [8-1:0] node853;
	wire [8-1:0] node856;
	wire [8-1:0] node857;
	wire [8-1:0] node861;
	wire [8-1:0] node863;
	wire [8-1:0] node866;
	wire [8-1:0] node867;
	wire [8-1:0] node868;
	wire [8-1:0] node869;
	wire [8-1:0] node870;
	wire [8-1:0] node871;
	wire [8-1:0] node875;
	wire [8-1:0] node876;
	wire [8-1:0] node878;
	wire [8-1:0] node881;
	wire [8-1:0] node884;
	wire [8-1:0] node885;
	wire [8-1:0] node886;
	wire [8-1:0] node890;
	wire [8-1:0] node892;
	wire [8-1:0] node893;
	wire [8-1:0] node896;
	wire [8-1:0] node899;
	wire [8-1:0] node900;
	wire [8-1:0] node901;
	wire [8-1:0] node902;
	wire [8-1:0] node903;
	wire [8-1:0] node907;
	wire [8-1:0] node909;
	wire [8-1:0] node912;
	wire [8-1:0] node913;
	wire [8-1:0] node914;
	wire [8-1:0] node918;
	wire [8-1:0] node919;
	wire [8-1:0] node922;
	wire [8-1:0] node925;
	wire [8-1:0] node926;
	wire [8-1:0] node928;
	wire [8-1:0] node931;
	wire [8-1:0] node932;
	wire [8-1:0] node933;
	wire [8-1:0] node937;
	wire [8-1:0] node939;
	wire [8-1:0] node942;
	wire [8-1:0] node943;
	wire [8-1:0] node944;
	wire [8-1:0] node946;
	wire [8-1:0] node949;
	wire [8-1:0] node950;
	wire [8-1:0] node953;
	wire [8-1:0] node955;
	wire [8-1:0] node958;
	wire [8-1:0] node959;
	wire [8-1:0] node960;
	wire [8-1:0] node961;
	wire [8-1:0] node964;
	wire [8-1:0] node965;
	wire [8-1:0] node969;
	wire [8-1:0] node970;
	wire [8-1:0] node971;
	wire [8-1:0] node975;
	wire [8-1:0] node976;
	wire [8-1:0] node979;
	wire [8-1:0] node982;
	wire [8-1:0] node983;
	wire [8-1:0] node984;
	wire [8-1:0] node985;
	wire [8-1:0] node988;
	wire [8-1:0] node991;
	wire [8-1:0] node993;
	wire [8-1:0] node996;
	wire [8-1:0] node997;
	wire [8-1:0] node998;
	wire [8-1:0] node1001;
	wire [8-1:0] node1004;
	wire [8-1:0] node1005;
	wire [8-1:0] node1008;
	wire [8-1:0] node1011;
	wire [8-1:0] node1012;
	wire [8-1:0] node1013;
	wire [8-1:0] node1014;
	wire [8-1:0] node1015;
	wire [8-1:0] node1016;
	wire [8-1:0] node1017;
	wire [8-1:0] node1020;
	wire [8-1:0] node1023;
	wire [8-1:0] node1024;
	wire [8-1:0] node1025;
	wire [8-1:0] node1029;
	wire [8-1:0] node1030;
	wire [8-1:0] node1033;
	wire [8-1:0] node1036;
	wire [8-1:0] node1037;
	wire [8-1:0] node1040;
	wire [8-1:0] node1041;
	wire [8-1:0] node1044;
	wire [8-1:0] node1047;
	wire [8-1:0] node1048;
	wire [8-1:0] node1049;
	wire [8-1:0] node1050;
	wire [8-1:0] node1054;
	wire [8-1:0] node1055;
	wire [8-1:0] node1056;
	wire [8-1:0] node1059;
	wire [8-1:0] node1062;
	wire [8-1:0] node1064;
	wire [8-1:0] node1067;
	wire [8-1:0] node1068;
	wire [8-1:0] node1069;
	wire [8-1:0] node1072;
	wire [8-1:0] node1075;
	wire [8-1:0] node1076;
	wire [8-1:0] node1077;
	wire [8-1:0] node1081;
	wire [8-1:0] node1083;
	wire [8-1:0] node1086;
	wire [8-1:0] node1087;
	wire [8-1:0] node1088;
	wire [8-1:0] node1089;
	wire [8-1:0] node1093;
	wire [8-1:0] node1094;
	wire [8-1:0] node1097;
	wire [8-1:0] node1100;
	wire [8-1:0] node1101;
	wire [8-1:0] node1102;
	wire [8-1:0] node1106;
	wire [8-1:0] node1107;
	wire [8-1:0] node1110;
	wire [8-1:0] node1113;
	wire [8-1:0] node1114;
	wire [8-1:0] node1115;
	wire [8-1:0] node1116;
	wire [8-1:0] node1117;
	wire [8-1:0] node1118;
	wire [8-1:0] node1119;
	wire [8-1:0] node1123;
	wire [8-1:0] node1125;
	wire [8-1:0] node1128;
	wire [8-1:0] node1130;
	wire [8-1:0] node1133;
	wire [8-1:0] node1134;
	wire [8-1:0] node1135;
	wire [8-1:0] node1136;
	wire [8-1:0] node1139;
	wire [8-1:0] node1142;
	wire [8-1:0] node1143;
	wire [8-1:0] node1146;
	wire [8-1:0] node1149;
	wire [8-1:0] node1152;
	wire [8-1:0] node1153;
	wire [8-1:0] node1154;
	wire [8-1:0] node1155;
	wire [8-1:0] node1156;
	wire [8-1:0] node1159;
	wire [8-1:0] node1162;
	wire [8-1:0] node1164;
	wire [8-1:0] node1167;
	wire [8-1:0] node1168;
	wire [8-1:0] node1169;
	wire [8-1:0] node1172;
	wire [8-1:0] node1175;
	wire [8-1:0] node1176;
	wire [8-1:0] node1180;
	wire [8-1:0] node1181;
	wire [8-1:0] node1182;
	wire [8-1:0] node1185;
	wire [8-1:0] node1188;
	wire [8-1:0] node1191;
	wire [8-1:0] node1192;
	wire [8-1:0] node1193;
	wire [8-1:0] node1194;
	wire [8-1:0] node1195;
	wire [8-1:0] node1196;
	wire [8-1:0] node1199;
	wire [8-1:0] node1203;
	wire [8-1:0] node1204;
	wire [8-1:0] node1206;
	wire [8-1:0] node1209;
	wire [8-1:0] node1211;
	wire [8-1:0] node1214;
	wire [8-1:0] node1215;
	wire [8-1:0] node1216;
	wire [8-1:0] node1217;
	wire [8-1:0] node1222;
	wire [8-1:0] node1223;
	wire [8-1:0] node1224;
	wire [8-1:0] node1227;
	wire [8-1:0] node1231;
	wire [8-1:0] node1232;
	wire [8-1:0] node1233;
	wire [8-1:0] node1234;
	wire [8-1:0] node1235;
	wire [8-1:0] node1238;
	wire [8-1:0] node1241;
	wire [8-1:0] node1242;
	wire [8-1:0] node1245;
	wire [8-1:0] node1248;
	wire [8-1:0] node1249;
	wire [8-1:0] node1250;
	wire [8-1:0] node1253;
	wire [8-1:0] node1256;
	wire [8-1:0] node1257;
	wire [8-1:0] node1260;
	wire [8-1:0] node1263;
	wire [8-1:0] node1266;
	wire [8-1:0] node1267;
	wire [8-1:0] node1268;
	wire [8-1:0] node1269;
	wire [8-1:0] node1270;
	wire [8-1:0] node1272;
	wire [8-1:0] node1273;
	wire [8-1:0] node1277;
	wire [8-1:0] node1278;
	wire [8-1:0] node1279;
	wire [8-1:0] node1283;
	wire [8-1:0] node1284;
	wire [8-1:0] node1285;
	wire [8-1:0] node1288;
	wire [8-1:0] node1292;
	wire [8-1:0] node1293;
	wire [8-1:0] node1294;
	wire [8-1:0] node1295;
	wire [8-1:0] node1296;
	wire [8-1:0] node1299;
	wire [8-1:0] node1301;
	wire [8-1:0] node1304;
	wire [8-1:0] node1305;
	wire [8-1:0] node1308;
	wire [8-1:0] node1309;
	wire [8-1:0] node1313;
	wire [8-1:0] node1314;
	wire [8-1:0] node1315;
	wire [8-1:0] node1316;
	wire [8-1:0] node1319;
	wire [8-1:0] node1322;
	wire [8-1:0] node1324;
	wire [8-1:0] node1327;
	wire [8-1:0] node1328;
	wire [8-1:0] node1332;
	wire [8-1:0] node1333;
	wire [8-1:0] node1334;
	wire [8-1:0] node1335;
	wire [8-1:0] node1336;
	wire [8-1:0] node1339;
	wire [8-1:0] node1342;
	wire [8-1:0] node1343;
	wire [8-1:0] node1344;
	wire [8-1:0] node1348;
	wire [8-1:0] node1349;
	wire [8-1:0] node1352;
	wire [8-1:0] node1355;
	wire [8-1:0] node1356;
	wire [8-1:0] node1357;
	wire [8-1:0] node1358;
	wire [8-1:0] node1361;
	wire [8-1:0] node1365;
	wire [8-1:0] node1366;
	wire [8-1:0] node1367;
	wire [8-1:0] node1370;
	wire [8-1:0] node1373;
	wire [8-1:0] node1374;
	wire [8-1:0] node1377;
	wire [8-1:0] node1380;
	wire [8-1:0] node1381;
	wire [8-1:0] node1382;
	wire [8-1:0] node1383;
	wire [8-1:0] node1387;
	wire [8-1:0] node1388;
	wire [8-1:0] node1392;
	wire [8-1:0] node1393;
	wire [8-1:0] node1397;
	wire [8-1:0] node1398;
	wire [8-1:0] node1399;
	wire [8-1:0] node1400;
	wire [8-1:0] node1401;
	wire [8-1:0] node1402;
	wire [8-1:0] node1403;
	wire [8-1:0] node1407;
	wire [8-1:0] node1409;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1417;
	wire [8-1:0] node1418;
	wire [8-1:0] node1419;
	wire [8-1:0] node1420;
	wire [8-1:0] node1421;
	wire [8-1:0] node1424;
	wire [8-1:0] node1427;
	wire [8-1:0] node1428;
	wire [8-1:0] node1431;
	wire [8-1:0] node1434;
	wire [8-1:0] node1435;
	wire [8-1:0] node1436;
	wire [8-1:0] node1440;
	wire [8-1:0] node1442;
	wire [8-1:0] node1445;
	wire [8-1:0] node1446;
	wire [8-1:0] node1447;
	wire [8-1:0] node1448;
	wire [8-1:0] node1451;
	wire [8-1:0] node1454;
	wire [8-1:0] node1456;
	wire [8-1:0] node1459;
	wire [8-1:0] node1460;
	wire [8-1:0] node1462;
	wire [8-1:0] node1465;
	wire [8-1:0] node1466;
	wire [8-1:0] node1469;
	wire [8-1:0] node1472;
	wire [8-1:0] node1473;
	wire [8-1:0] node1474;
	wire [8-1:0] node1476;
	wire [8-1:0] node1479;
	wire [8-1:0] node1480;
	wire [8-1:0] node1481;
	wire [8-1:0] node1485;
	wire [8-1:0] node1486;
	wire [8-1:0] node1490;
	wire [8-1:0] node1491;
	wire [8-1:0] node1492;
	wire [8-1:0] node1493;
	wire [8-1:0] node1496;
	wire [8-1:0] node1499;
	wire [8-1:0] node1500;
	wire [8-1:0] node1501;
	wire [8-1:0] node1504;
	wire [8-1:0] node1507;
	wire [8-1:0] node1509;
	wire [8-1:0] node1512;
	wire [8-1:0] node1513;
	wire [8-1:0] node1514;
	wire [8-1:0] node1517;
	wire [8-1:0] node1520;
	wire [8-1:0] node1521;
	wire [8-1:0] node1522;
	wire [8-1:0] node1525;
	wire [8-1:0] node1528;
	wire [8-1:0] node1529;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1536;
	wire [8-1:0] node1537;
	wire [8-1:0] node1539;
	wire [8-1:0] node1540;
	wire [8-1:0] node1543;
	wire [8-1:0] node1546;
	wire [8-1:0] node1548;
	wire [8-1:0] node1551;
	wire [8-1:0] node1552;
	wire [8-1:0] node1554;
	wire [8-1:0] node1558;
	wire [8-1:0] node1559;
	wire [8-1:0] node1560;
	wire [8-1:0] node1561;
	wire [8-1:0] node1562;
	wire [8-1:0] node1563;
	wire [8-1:0] node1564;
	wire [8-1:0] node1567;
	wire [8-1:0] node1570;
	wire [8-1:0] node1571;
	wire [8-1:0] node1572;
	wire [8-1:0] node1574;
	wire [8-1:0] node1577;
	wire [8-1:0] node1579;
	wire [8-1:0] node1582;
	wire [8-1:0] node1583;
	wire [8-1:0] node1585;
	wire [8-1:0] node1588;
	wire [8-1:0] node1590;
	wire [8-1:0] node1593;
	wire [8-1:0] node1594;
	wire [8-1:0] node1595;
	wire [8-1:0] node1598;
	wire [8-1:0] node1601;
	wire [8-1:0] node1602;
	wire [8-1:0] node1604;
	wire [8-1:0] node1607;
	wire [8-1:0] node1608;
	wire [8-1:0] node1611;
	wire [8-1:0] node1612;
	wire [8-1:0] node1616;
	wire [8-1:0] node1617;
	wire [8-1:0] node1618;
	wire [8-1:0] node1619;
	wire [8-1:0] node1621;
	wire [8-1:0] node1624;
	wire [8-1:0] node1625;
	wire [8-1:0] node1626;
	wire [8-1:0] node1630;
	wire [8-1:0] node1632;
	wire [8-1:0] node1635;
	wire [8-1:0] node1636;
	wire [8-1:0] node1637;
	wire [8-1:0] node1639;
	wire [8-1:0] node1642;
	wire [8-1:0] node1644;
	wire [8-1:0] node1647;
	wire [8-1:0] node1648;
	wire [8-1:0] node1650;
	wire [8-1:0] node1653;
	wire [8-1:0] node1654;
	wire [8-1:0] node1658;
	wire [8-1:0] node1659;
	wire [8-1:0] node1660;
	wire [8-1:0] node1661;
	wire [8-1:0] node1665;
	wire [8-1:0] node1666;
	wire [8-1:0] node1667;
	wire [8-1:0] node1670;
	wire [8-1:0] node1673;
	wire [8-1:0] node1675;
	wire [8-1:0] node1678;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1683;
	wire [8-1:0] node1686;
	wire [8-1:0] node1687;
	wire [8-1:0] node1688;
	wire [8-1:0] node1692;
	wire [8-1:0] node1693;
	wire [8-1:0] node1697;
	wire [8-1:0] node1698;
	wire [8-1:0] node1699;
	wire [8-1:0] node1700;
	wire [8-1:0] node1701;
	wire [8-1:0] node1704;
	wire [8-1:0] node1707;
	wire [8-1:0] node1708;
	wire [8-1:0] node1709;
	wire [8-1:0] node1711;
	wire [8-1:0] node1715;
	wire [8-1:0] node1716;
	wire [8-1:0] node1718;
	wire [8-1:0] node1721;
	wire [8-1:0] node1723;
	wire [8-1:0] node1726;
	wire [8-1:0] node1727;
	wire [8-1:0] node1728;
	wire [8-1:0] node1731;
	wire [8-1:0] node1734;
	wire [8-1:0] node1735;
	wire [8-1:0] node1736;
	wire [8-1:0] node1738;
	wire [8-1:0] node1741;
	wire [8-1:0] node1742;
	wire [8-1:0] node1746;
	wire [8-1:0] node1747;
	wire [8-1:0] node1749;
	wire [8-1:0] node1752;
	wire [8-1:0] node1754;
	wire [8-1:0] node1757;
	wire [8-1:0] node1758;
	wire [8-1:0] node1759;
	wire [8-1:0] node1760;
	wire [8-1:0] node1762;
	wire [8-1:0] node1765;
	wire [8-1:0] node1766;
	wire [8-1:0] node1769;
	wire [8-1:0] node1771;
	wire [8-1:0] node1774;
	wire [8-1:0] node1775;
	wire [8-1:0] node1776;
	wire [8-1:0] node1778;
	wire [8-1:0] node1781;
	wire [8-1:0] node1782;
	wire [8-1:0] node1786;
	wire [8-1:0] node1787;
	wire [8-1:0] node1788;
	wire [8-1:0] node1793;
	wire [8-1:0] node1794;
	wire [8-1:0] node1795;
	wire [8-1:0] node1796;
	wire [8-1:0] node1800;
	wire [8-1:0] node1801;
	wire [8-1:0] node1804;
	wire [8-1:0] node1805;
	wire [8-1:0] node1808;
	wire [8-1:0] node1811;
	wire [8-1:0] node1812;
	wire [8-1:0] node1814;
	wire [8-1:0] node1815;
	wire [8-1:0] node1819;
	wire [8-1:0] node1820;
	wire [8-1:0] node1821;
	wire [8-1:0] node1824;
	wire [8-1:0] node1828;
	wire [8-1:0] node1829;
	wire [8-1:0] node1830;
	wire [8-1:0] node1831;
	wire [8-1:0] node1832;
	wire [8-1:0] node1834;
	wire [8-1:0] node1837;
	wire [8-1:0] node1838;
	wire [8-1:0] node1840;
	wire [8-1:0] node1843;
	wire [8-1:0] node1845;
	wire [8-1:0] node1848;
	wire [8-1:0] node1849;
	wire [8-1:0] node1850;
	wire [8-1:0] node1851;
	wire [8-1:0] node1855;
	wire [8-1:0] node1856;
	wire [8-1:0] node1859;
	wire [8-1:0] node1860;
	wire [8-1:0] node1863;
	wire [8-1:0] node1866;
	wire [8-1:0] node1867;
	wire [8-1:0] node1868;
	wire [8-1:0] node1872;
	wire [8-1:0] node1873;
	wire [8-1:0] node1876;
	wire [8-1:0] node1879;
	wire [8-1:0] node1880;
	wire [8-1:0] node1881;
	wire [8-1:0] node1882;
	wire [8-1:0] node1886;
	wire [8-1:0] node1887;
	wire [8-1:0] node1888;
	wire [8-1:0] node1892;
	wire [8-1:0] node1893;
	wire [8-1:0] node1897;
	wire [8-1:0] node1898;
	wire [8-1:0] node1899;
	wire [8-1:0] node1901;
	wire [8-1:0] node1904;
	wire [8-1:0] node1906;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1911;
	wire [8-1:0] node1912;
	wire [8-1:0] node1915;
	wire [8-1:0] node1918;
	wire [8-1:0] node1919;
	wire [8-1:0] node1922;
	wire [8-1:0] node1925;
	wire [8-1:0] node1926;
	wire [8-1:0] node1929;
	wire [8-1:0] node1932;
	wire [8-1:0] node1933;
	wire [8-1:0] node1934;
	wire [8-1:0] node1935;
	wire [8-1:0] node1936;
	wire [8-1:0] node1937;
	wire [8-1:0] node1940;
	wire [8-1:0] node1943;
	wire [8-1:0] node1944;
	wire [8-1:0] node1946;
	wire [8-1:0] node1949;
	wire [8-1:0] node1950;
	wire [8-1:0] node1954;
	wire [8-1:0] node1955;
	wire [8-1:0] node1956;
	wire [8-1:0] node1959;
	wire [8-1:0] node1962;
	wire [8-1:0] node1963;
	wire [8-1:0] node1965;
	wire [8-1:0] node1968;
	wire [8-1:0] node1970;
	wire [8-1:0] node1973;
	wire [8-1:0] node1974;
	wire [8-1:0] node1975;
	wire [8-1:0] node1976;
	wire [8-1:0] node1977;
	wire [8-1:0] node1980;
	wire [8-1:0] node1983;
	wire [8-1:0] node1984;
	wire [8-1:0] node1987;
	wire [8-1:0] node1990;
	wire [8-1:0] node1991;
	wire [8-1:0] node1992;
	wire [8-1:0] node1995;
	wire [8-1:0] node1998;
	wire [8-1:0] node1999;
	wire [8-1:0] node2003;
	wire [8-1:0] node2004;
	wire [8-1:0] node2005;
	wire [8-1:0] node2006;
	wire [8-1:0] node2009;
	wire [8-1:0] node2012;
	wire [8-1:0] node2015;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2021;
	wire [8-1:0] node2024;
	wire [8-1:0] node2025;
	wire [8-1:0] node2026;
	wire [8-1:0] node2027;
	wire [8-1:0] node2028;
	wire [8-1:0] node2029;
	wire [8-1:0] node2032;
	wire [8-1:0] node2035;
	wire [8-1:0] node2036;
	wire [8-1:0] node2039;
	wire [8-1:0] node2042;
	wire [8-1:0] node2044;
	wire [8-1:0] node2045;
	wire [8-1:0] node2048;
	wire [8-1:0] node2051;
	wire [8-1:0] node2052;
	wire [8-1:0] node2053;
	wire [8-1:0] node2054;
	wire [8-1:0] node2057;
	wire [8-1:0] node2060;
	wire [8-1:0] node2062;
	wire [8-1:0] node2065;
	wire [8-1:0] node2066;
	wire [8-1:0] node2067;
	wire [8-1:0] node2070;
	wire [8-1:0] node2073;
	wire [8-1:0] node2074;
	wire [8-1:0] node2077;
	wire [8-1:0] node2080;
	wire [8-1:0] node2081;
	wire [8-1:0] node2082;
	wire [8-1:0] node2085;
	wire [8-1:0] node2088;
	wire [8-1:0] node2091;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2094;
	wire [8-1:0] node2095;
	wire [8-1:0] node2096;
	wire [8-1:0] node2097;
	wire [8-1:0] node2098;
	wire [8-1:0] node2102;
	wire [8-1:0] node2104;
	wire [8-1:0] node2107;
	wire [8-1:0] node2108;
	wire [8-1:0] node2109;
	wire [8-1:0] node2113;
	wire [8-1:0] node2115;
	wire [8-1:0] node2118;
	wire [8-1:0] node2119;
	wire [8-1:0] node2120;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2124;
	wire [8-1:0] node2125;
	wire [8-1:0] node2129;
	wire [8-1:0] node2131;
	wire [8-1:0] node2134;
	wire [8-1:0] node2135;
	wire [8-1:0] node2136;
	wire [8-1:0] node2140;
	wire [8-1:0] node2141;
	wire [8-1:0] node2143;
	wire [8-1:0] node2146;
	wire [8-1:0] node2147;
	wire [8-1:0] node2151;
	wire [8-1:0] node2152;
	wire [8-1:0] node2153;
	wire [8-1:0] node2157;
	wire [8-1:0] node2158;
	wire [8-1:0] node2159;
	wire [8-1:0] node2163;
	wire [8-1:0] node2164;
	wire [8-1:0] node2168;
	wire [8-1:0] node2169;
	wire [8-1:0] node2170;
	wire [8-1:0] node2171;
	wire [8-1:0] node2172;
	wire [8-1:0] node2176;
	wire [8-1:0] node2177;
	wire [8-1:0] node2179;
	wire [8-1:0] node2182;
	wire [8-1:0] node2185;
	wire [8-1:0] node2186;
	wire [8-1:0] node2187;
	wire [8-1:0] node2188;
	wire [8-1:0] node2192;
	wire [8-1:0] node2194;
	wire [8-1:0] node2197;
	wire [8-1:0] node2199;
	wire [8-1:0] node2202;
	wire [8-1:0] node2203;
	wire [8-1:0] node2204;
	wire [8-1:0] node2206;
	wire [8-1:0] node2209;
	wire [8-1:0] node2211;
	wire [8-1:0] node2214;
	wire [8-1:0] node2216;
	wire [8-1:0] node2219;
	wire [8-1:0] node2220;
	wire [8-1:0] node2221;
	wire [8-1:0] node2222;
	wire [8-1:0] node2223;
	wire [8-1:0] node2227;
	wire [8-1:0] node2228;
	wire [8-1:0] node2232;
	wire [8-1:0] node2233;
	wire [8-1:0] node2234;
	wire [8-1:0] node2235;
	wire [8-1:0] node2237;
	wire [8-1:0] node2240;
	wire [8-1:0] node2242;
	wire [8-1:0] node2245;
	wire [8-1:0] node2246;
	wire [8-1:0] node2250;
	wire [8-1:0] node2251;
	wire [8-1:0] node2253;
	wire [8-1:0] node2256;
	wire [8-1:0] node2257;
	wire [8-1:0] node2259;
	wire [8-1:0] node2262;
	wire [8-1:0] node2264;
	wire [8-1:0] node2267;
	wire [8-1:0] node2268;
	wire [8-1:0] node2269;
	wire [8-1:0] node2270;
	wire [8-1:0] node2274;
	wire [8-1:0] node2275;
	wire [8-1:0] node2276;
	wire [8-1:0] node2280;
	wire [8-1:0] node2281;
	wire [8-1:0] node2285;
	wire [8-1:0] node2286;
	wire [8-1:0] node2290;
	wire [8-1:0] node2291;
	wire [8-1:0] node2292;
	wire [8-1:0] node2293;
	wire [8-1:0] node2294;
	wire [8-1:0] node2295;
	wire [8-1:0] node2296;
	wire [8-1:0] node2297;
	wire [8-1:0] node2301;
	wire [8-1:0] node2303;
	wire [8-1:0] node2306;
	wire [8-1:0] node2308;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2313;
	wire [8-1:0] node2316;
	wire [8-1:0] node2317;
	wire [8-1:0] node2320;
	wire [8-1:0] node2323;
	wire [8-1:0] node2324;
	wire [8-1:0] node2325;
	wire [8-1:0] node2328;
	wire [8-1:0] node2329;
	wire [8-1:0] node2332;
	wire [8-1:0] node2335;
	wire [8-1:0] node2336;
	wire [8-1:0] node2339;
	wire [8-1:0] node2340;
	wire [8-1:0] node2343;
	wire [8-1:0] node2346;
	wire [8-1:0] node2347;
	wire [8-1:0] node2348;
	wire [8-1:0] node2349;
	wire [8-1:0] node2350;
	wire [8-1:0] node2353;
	wire [8-1:0] node2356;
	wire [8-1:0] node2357;
	wire [8-1:0] node2360;
	wire [8-1:0] node2362;
	wire [8-1:0] node2365;
	wire [8-1:0] node2366;
	wire [8-1:0] node2367;
	wire [8-1:0] node2368;
	wire [8-1:0] node2371;
	wire [8-1:0] node2373;
	wire [8-1:0] node2376;
	wire [8-1:0] node2377;
	wire [8-1:0] node2378;
	wire [8-1:0] node2381;
	wire [8-1:0] node2384;
	wire [8-1:0] node2386;
	wire [8-1:0] node2389;
	wire [8-1:0] node2390;
	wire [8-1:0] node2391;
	wire [8-1:0] node2393;
	wire [8-1:0] node2396;
	wire [8-1:0] node2397;
	wire [8-1:0] node2400;
	wire [8-1:0] node2403;
	wire [8-1:0] node2404;
	wire [8-1:0] node2405;
	wire [8-1:0] node2408;
	wire [8-1:0] node2411;
	wire [8-1:0] node2412;
	wire [8-1:0] node2415;
	wire [8-1:0] node2418;
	wire [8-1:0] node2419;
	wire [8-1:0] node2420;
	wire [8-1:0] node2423;
	wire [8-1:0] node2426;
	wire [8-1:0] node2427;
	wire [8-1:0] node2428;
	wire [8-1:0] node2429;
	wire [8-1:0] node2430;
	wire [8-1:0] node2433;
	wire [8-1:0] node2436;
	wire [8-1:0] node2437;
	wire [8-1:0] node2441;
	wire [8-1:0] node2442;
	wire [8-1:0] node2444;
	wire [8-1:0] node2447;
	wire [8-1:0] node2449;
	wire [8-1:0] node2452;
	wire [8-1:0] node2453;
	wire [8-1:0] node2454;
	wire [8-1:0] node2456;
	wire [8-1:0] node2459;
	wire [8-1:0] node2461;
	wire [8-1:0] node2464;
	wire [8-1:0] node2465;
	wire [8-1:0] node2467;
	wire [8-1:0] node2470;
	wire [8-1:0] node2472;
	wire [8-1:0] node2475;
	wire [8-1:0] node2476;
	wire [8-1:0] node2477;
	wire [8-1:0] node2478;
	wire [8-1:0] node2479;
	wire [8-1:0] node2480;
	wire [8-1:0] node2484;
	wire [8-1:0] node2485;
	wire [8-1:0] node2488;
	wire [8-1:0] node2489;
	wire [8-1:0] node2492;
	wire [8-1:0] node2495;
	wire [8-1:0] node2496;
	wire [8-1:0] node2497;
	wire [8-1:0] node2498;
	wire [8-1:0] node2502;
	wire [8-1:0] node2503;
	wire [8-1:0] node2505;
	wire [8-1:0] node2508;
	wire [8-1:0] node2511;
	wire [8-1:0] node2512;
	wire [8-1:0] node2515;
	wire [8-1:0] node2516;
	wire [8-1:0] node2518;
	wire [8-1:0] node2521;
	wire [8-1:0] node2523;
	wire [8-1:0] node2526;
	wire [8-1:0] node2527;
	wire [8-1:0] node2528;
	wire [8-1:0] node2529;
	wire [8-1:0] node2530;
	wire [8-1:0] node2531;
	wire [8-1:0] node2535;
	wire [8-1:0] node2536;
	wire [8-1:0] node2540;
	wire [8-1:0] node2542;
	wire [8-1:0] node2545;
	wire [8-1:0] node2546;
	wire [8-1:0] node2547;
	wire [8-1:0] node2551;
	wire [8-1:0] node2552;
	wire [8-1:0] node2555;
	wire [8-1:0] node2558;
	wire [8-1:0] node2559;
	wire [8-1:0] node2560;
	wire [8-1:0] node2561;
	wire [8-1:0] node2565;
	wire [8-1:0] node2568;
	wire [8-1:0] node2569;
	wire [8-1:0] node2570;
	wire [8-1:0] node2572;
	wire [8-1:0] node2575;
	wire [8-1:0] node2576;
	wire [8-1:0] node2580;
	wire [8-1:0] node2581;
	wire [8-1:0] node2584;
	wire [8-1:0] node2587;
	wire [8-1:0] node2588;
	wire [8-1:0] node2589;
	wire [8-1:0] node2590;
	wire [8-1:0] node2591;
	wire [8-1:0] node2592;
	wire [8-1:0] node2597;
	wire [8-1:0] node2598;
	wire [8-1:0] node2599;
	wire [8-1:0] node2603;
	wire [8-1:0] node2604;
	wire [8-1:0] node2608;
	wire [8-1:0] node2609;
	wire [8-1:0] node2610;
	wire [8-1:0] node2611;
	wire [8-1:0] node2615;
	wire [8-1:0] node2616;
	wire [8-1:0] node2620;
	wire [8-1:0] node2622;
	wire [8-1:0] node2625;
	wire [8-1:0] node2626;
	wire [8-1:0] node2627;
	wire [8-1:0] node2628;
	wire [8-1:0] node2631;
	wire [8-1:0] node2632;
	wire [8-1:0] node2635;
	wire [8-1:0] node2638;
	wire [8-1:0] node2639;
	wire [8-1:0] node2640;
	wire [8-1:0] node2641;
	wire [8-1:0] node2644;
	wire [8-1:0] node2647;
	wire [8-1:0] node2648;
	wire [8-1:0] node2652;
	wire [8-1:0] node2653;
	wire [8-1:0] node2655;
	wire [8-1:0] node2658;
	wire [8-1:0] node2661;
	wire [8-1:0] node2662;
	wire [8-1:0] node2663;
	wire [8-1:0] node2664;
	wire [8-1:0] node2667;
	wire [8-1:0] node2669;
	wire [8-1:0] node2672;
	wire [8-1:0] node2673;
	wire [8-1:0] node2674;
	wire [8-1:0] node2677;
	wire [8-1:0] node2680;
	wire [8-1:0] node2683;
	wire [8-1:0] node2684;
	wire [8-1:0] node2685;
	wire [8-1:0] node2688;
	wire [8-1:0] node2691;
	wire [8-1:0] node2692;
	wire [8-1:0] node2695;
	wire [8-1:0] node2698;
	wire [8-1:0] node2699;
	wire [8-1:0] node2700;
	wire [8-1:0] node2701;
	wire [8-1:0] node2702;
	wire [8-1:0] node2703;
	wire [8-1:0] node2704;
	wire [8-1:0] node2706;
	wire [8-1:0] node2709;
	wire [8-1:0] node2711;
	wire [8-1:0] node2714;
	wire [8-1:0] node2715;
	wire [8-1:0] node2717;
	wire [8-1:0] node2720;
	wire [8-1:0] node2722;
	wire [8-1:0] node2725;
	wire [8-1:0] node2727;
	wire [8-1:0] node2730;
	wire [8-1:0] node2731;
	wire [8-1:0] node2732;
	wire [8-1:0] node2733;
	wire [8-1:0] node2736;
	wire [8-1:0] node2738;
	wire [8-1:0] node2741;
	wire [8-1:0] node2744;
	wire [8-1:0] node2745;
	wire [8-1:0] node2747;
	wire [8-1:0] node2749;
	wire [8-1:0] node2752;
	wire [8-1:0] node2754;
	wire [8-1:0] node2757;
	wire [8-1:0] node2758;
	wire [8-1:0] node2759;
	wire [8-1:0] node2760;
	wire [8-1:0] node2761;
	wire [8-1:0] node2765;
	wire [8-1:0] node2767;
	wire [8-1:0] node2768;
	wire [8-1:0] node2771;
	wire [8-1:0] node2774;
	wire [8-1:0] node2775;
	wire [8-1:0] node2778;
	wire [8-1:0] node2780;
	wire [8-1:0] node2783;
	wire [8-1:0] node2784;
	wire [8-1:0] node2785;
	wire [8-1:0] node2787;
	wire [8-1:0] node2789;
	wire [8-1:0] node2792;
	wire [8-1:0] node2794;
	wire [8-1:0] node2797;
	wire [8-1:0] node2799;
	wire [8-1:0] node2801;
	wire [8-1:0] node2804;
	wire [8-1:0] node2805;
	wire [8-1:0] node2806;
	wire [8-1:0] node2807;
	wire [8-1:0] node2808;
	wire [8-1:0] node2811;
	wire [8-1:0] node2812;
	wire [8-1:0] node2815;
	wire [8-1:0] node2818;
	wire [8-1:0] node2819;
	wire [8-1:0] node2820;
	wire [8-1:0] node2823;
	wire [8-1:0] node2824;
	wire [8-1:0] node2827;
	wire [8-1:0] node2830;
	wire [8-1:0] node2831;
	wire [8-1:0] node2834;
	wire [8-1:0] node2835;
	wire [8-1:0] node2838;
	wire [8-1:0] node2841;
	wire [8-1:0] node2842;
	wire [8-1:0] node2843;
	wire [8-1:0] node2844;
	wire [8-1:0] node2845;
	wire [8-1:0] node2846;
	wire [8-1:0] node2849;
	wire [8-1:0] node2852;
	wire [8-1:0] node2853;
	wire [8-1:0] node2856;
	wire [8-1:0] node2859;
	wire [8-1:0] node2860;
	wire [8-1:0] node2861;
	wire [8-1:0] node2865;
	wire [8-1:0] node2866;
	wire [8-1:0] node2870;
	wire [8-1:0] node2871;
	wire [8-1:0] node2872;
	wire [8-1:0] node2873;
	wire [8-1:0] node2876;
	wire [8-1:0] node2879;
	wire [8-1:0] node2880;
	wire [8-1:0] node2884;
	wire [8-1:0] node2885;
	wire [8-1:0] node2886;
	wire [8-1:0] node2890;
	wire [8-1:0] node2891;
	wire [8-1:0] node2894;
	wire [8-1:0] node2897;
	wire [8-1:0] node2898;
	wire [8-1:0] node2899;
	wire [8-1:0] node2900;
	wire [8-1:0] node2901;
	wire [8-1:0] node2904;
	wire [8-1:0] node2907;
	wire [8-1:0] node2908;
	wire [8-1:0] node2911;
	wire [8-1:0] node2914;
	wire [8-1:0] node2915;
	wire [8-1:0] node2916;
	wire [8-1:0] node2919;
	wire [8-1:0] node2922;
	wire [8-1:0] node2923;
	wire [8-1:0] node2926;
	wire [8-1:0] node2929;
	wire [8-1:0] node2930;
	wire [8-1:0] node2931;
	wire [8-1:0] node2932;
	wire [8-1:0] node2935;
	wire [8-1:0] node2938;
	wire [8-1:0] node2941;
	wire [8-1:0] node2942;
	wire [8-1:0] node2944;
	wire [8-1:0] node2947;
	wire [8-1:0] node2949;
	wire [8-1:0] node2952;
	wire [8-1:0] node2953;
	wire [8-1:0] node2954;
	wire [8-1:0] node2955;
	wire [8-1:0] node2956;
	wire [8-1:0] node2959;
	wire [8-1:0] node2960;
	wire [8-1:0] node2963;
	wire [8-1:0] node2966;
	wire [8-1:0] node2967;
	wire [8-1:0] node2968;
	wire [8-1:0] node2969;
	wire [8-1:0] node2972;
	wire [8-1:0] node2975;
	wire [8-1:0] node2976;
	wire [8-1:0] node2979;
	wire [8-1:0] node2982;
	wire [8-1:0] node2983;
	wire [8-1:0] node2985;
	wire [8-1:0] node2988;
	wire [8-1:0] node2991;
	wire [8-1:0] node2992;
	wire [8-1:0] node2993;
	wire [8-1:0] node2994;
	wire [8-1:0] node2996;
	wire [8-1:0] node2999;
	wire [8-1:0] node3001;
	wire [8-1:0] node3004;
	wire [8-1:0] node3005;
	wire [8-1:0] node3008;
	wire [8-1:0] node3011;
	wire [8-1:0] node3012;
	wire [8-1:0] node3013;
	wire [8-1:0] node3014;
	wire [8-1:0] node3017;
	wire [8-1:0] node3020;
	wire [8-1:0] node3023;
	wire [8-1:0] node3024;
	wire [8-1:0] node3027;
	wire [8-1:0] node3030;
	wire [8-1:0] node3031;
	wire [8-1:0] node3032;
	wire [8-1:0] node3033;
	wire [8-1:0] node3036;
	wire [8-1:0] node3037;
	wire [8-1:0] node3039;
	wire [8-1:0] node3042;
	wire [8-1:0] node3043;
	wire [8-1:0] node3047;
	wire [8-1:0] node3048;
	wire [8-1:0] node3049;
	wire [8-1:0] node3052;
	wire [8-1:0] node3055;
	wire [8-1:0] node3056;
	wire [8-1:0] node3058;
	wire [8-1:0] node3061;
	wire [8-1:0] node3062;
	wire [8-1:0] node3066;
	wire [8-1:0] node3067;
	wire [8-1:0] node3068;
	wire [8-1:0] node3069;
	wire [8-1:0] node3071;
	wire [8-1:0] node3074;
	wire [8-1:0] node3077;
	wire [8-1:0] node3078;
	wire [8-1:0] node3080;
	wire [8-1:0] node3083;
	wire [8-1:0] node3084;
	wire [8-1:0] node3088;
	wire [8-1:0] node3089;
	wire [8-1:0] node3090;
	wire [8-1:0] node3093;
	wire [8-1:0] node3096;
	wire [8-1:0] node3097;
	wire [8-1:0] node3100;
	wire [8-1:0] node3103;
	wire [8-1:0] node3104;
	wire [8-1:0] node3105;
	wire [8-1:0] node3106;
	wire [8-1:0] node3107;
	wire [8-1:0] node3108;
	wire [8-1:0] node3109;
	wire [8-1:0] node3111;
	wire [8-1:0] node3114;
	wire [8-1:0] node3115;
	wire [8-1:0] node3117;
	wire [8-1:0] node3120;
	wire [8-1:0] node3122;
	wire [8-1:0] node3125;
	wire [8-1:0] node3126;
	wire [8-1:0] node3127;
	wire [8-1:0] node3129;
	wire [8-1:0] node3132;
	wire [8-1:0] node3133;
	wire [8-1:0] node3135;
	wire [8-1:0] node3138;
	wire [8-1:0] node3140;
	wire [8-1:0] node3143;
	wire [8-1:0] node3144;
	wire [8-1:0] node3146;
	wire [8-1:0] node3149;
	wire [8-1:0] node3150;
	wire [8-1:0] node3153;
	wire [8-1:0] node3154;
	wire [8-1:0] node3157;
	wire [8-1:0] node3160;
	wire [8-1:0] node3161;
	wire [8-1:0] node3162;
	wire [8-1:0] node3163;
	wire [8-1:0] node3164;
	wire [8-1:0] node3165;
	wire [8-1:0] node3168;
	wire [8-1:0] node3171;
	wire [8-1:0] node3172;
	wire [8-1:0] node3175;
	wire [8-1:0] node3178;
	wire [8-1:0] node3179;
	wire [8-1:0] node3180;
	wire [8-1:0] node3184;
	wire [8-1:0] node3185;
	wire [8-1:0] node3188;
	wire [8-1:0] node3191;
	wire [8-1:0] node3192;
	wire [8-1:0] node3193;
	wire [8-1:0] node3194;
	wire [8-1:0] node3197;
	wire [8-1:0] node3200;
	wire [8-1:0] node3201;
	wire [8-1:0] node3202;
	wire [8-1:0] node3205;
	wire [8-1:0] node3208;
	wire [8-1:0] node3209;
	wire [8-1:0] node3212;
	wire [8-1:0] node3215;
	wire [8-1:0] node3216;
	wire [8-1:0] node3217;
	wire [8-1:0] node3220;
	wire [8-1:0] node3223;
	wire [8-1:0] node3224;
	wire [8-1:0] node3227;
	wire [8-1:0] node3230;
	wire [8-1:0] node3231;
	wire [8-1:0] node3232;
	wire [8-1:0] node3233;
	wire [8-1:0] node3234;
	wire [8-1:0] node3238;
	wire [8-1:0] node3239;
	wire [8-1:0] node3242;
	wire [8-1:0] node3245;
	wire [8-1:0] node3246;
	wire [8-1:0] node3247;
	wire [8-1:0] node3248;
	wire [8-1:0] node3251;
	wire [8-1:0] node3254;
	wire [8-1:0] node3255;
	wire [8-1:0] node3258;
	wire [8-1:0] node3261;
	wire [8-1:0] node3262;
	wire [8-1:0] node3265;
	wire [8-1:0] node3268;
	wire [8-1:0] node3269;
	wire [8-1:0] node3270;
	wire [8-1:0] node3271;
	wire [8-1:0] node3274;
	wire [8-1:0] node3277;
	wire [8-1:0] node3278;
	wire [8-1:0] node3281;
	wire [8-1:0] node3284;
	wire [8-1:0] node3285;
	wire [8-1:0] node3286;
	wire [8-1:0] node3289;
	wire [8-1:0] node3292;
	wire [8-1:0] node3293;
	wire [8-1:0] node3296;
	wire [8-1:0] node3299;
	wire [8-1:0] node3300;
	wire [8-1:0] node3301;
	wire [8-1:0] node3302;
	wire [8-1:0] node3304;
	wire [8-1:0] node3307;
	wire [8-1:0] node3308;
	wire [8-1:0] node3310;
	wire [8-1:0] node3313;
	wire [8-1:0] node3315;
	wire [8-1:0] node3318;
	wire [8-1:0] node3319;
	wire [8-1:0] node3320;
	wire [8-1:0] node3321;
	wire [8-1:0] node3322;
	wire [8-1:0] node3324;
	wire [8-1:0] node3327;
	wire [8-1:0] node3328;
	wire [8-1:0] node3332;
	wire [8-1:0] node3333;
	wire [8-1:0] node3336;
	wire [8-1:0] node3339;
	wire [8-1:0] node3340;
	wire [8-1:0] node3341;
	wire [8-1:0] node3344;
	wire [8-1:0] node3347;
	wire [8-1:0] node3348;
	wire [8-1:0] node3349;
	wire [8-1:0] node3353;
	wire [8-1:0] node3356;
	wire [8-1:0] node3357;
	wire [8-1:0] node3358;
	wire [8-1:0] node3359;
	wire [8-1:0] node3361;
	wire [8-1:0] node3364;
	wire [8-1:0] node3365;
	wire [8-1:0] node3368;
	wire [8-1:0] node3371;
	wire [8-1:0] node3372;
	wire [8-1:0] node3373;
	wire [8-1:0] node3376;
	wire [8-1:0] node3379;
	wire [8-1:0] node3380;
	wire [8-1:0] node3383;
	wire [8-1:0] node3386;
	wire [8-1:0] node3387;
	wire [8-1:0] node3388;
	wire [8-1:0] node3391;
	wire [8-1:0] node3394;
	wire [8-1:0] node3395;
	wire [8-1:0] node3398;
	wire [8-1:0] node3401;
	wire [8-1:0] node3402;
	wire [8-1:0] node3403;
	wire [8-1:0] node3404;
	wire [8-1:0] node3406;
	wire [8-1:0] node3409;
	wire [8-1:0] node3410;
	wire [8-1:0] node3411;
	wire [8-1:0] node3414;
	wire [8-1:0] node3417;
	wire [8-1:0] node3418;
	wire [8-1:0] node3421;
	wire [8-1:0] node3424;
	wire [8-1:0] node3425;
	wire [8-1:0] node3426;
	wire [8-1:0] node3427;
	wire [8-1:0] node3431;
	wire [8-1:0] node3434;
	wire [8-1:0] node3435;
	wire [8-1:0] node3436;
	wire [8-1:0] node3440;
	wire [8-1:0] node3443;
	wire [8-1:0] node3444;
	wire [8-1:0] node3445;
	wire [8-1:0] node3447;
	wire [8-1:0] node3450;
	wire [8-1:0] node3451;
	wire [8-1:0] node3452;
	wire [8-1:0] node3453;
	wire [8-1:0] node3457;
	wire [8-1:0] node3459;
	wire [8-1:0] node3462;
	wire [8-1:0] node3463;
	wire [8-1:0] node3464;
	wire [8-1:0] node3467;
	wire [8-1:0] node3470;
	wire [8-1:0] node3471;
	wire [8-1:0] node3474;
	wire [8-1:0] node3477;
	wire [8-1:0] node3478;
	wire [8-1:0] node3479;
	wire [8-1:0] node3480;
	wire [8-1:0] node3484;
	wire [8-1:0] node3487;
	wire [8-1:0] node3488;
	wire [8-1:0] node3489;
	wire [8-1:0] node3491;
	wire [8-1:0] node3495;
	wire [8-1:0] node3497;
	wire [8-1:0] node3500;
	wire [8-1:0] node3501;
	wire [8-1:0] node3503;
	wire [8-1:0] node3505;
	wire [8-1:0] node3508;
	wire [8-1:0] node3509;
	wire [8-1:0] node3510;
	wire [8-1:0] node3511;
	wire [8-1:0] node3512;
	wire [8-1:0] node3513;
	wire [8-1:0] node3516;
	wire [8-1:0] node3519;
	wire [8-1:0] node3520;
	wire [8-1:0] node3524;
	wire [8-1:0] node3525;
	wire [8-1:0] node3529;
	wire [8-1:0] node3530;
	wire [8-1:0] node3531;
	wire [8-1:0] node3532;
	wire [8-1:0] node3536;
	wire [8-1:0] node3537;
	wire [8-1:0] node3540;
	wire [8-1:0] node3543;
	wire [8-1:0] node3544;
	wire [8-1:0] node3545;
	wire [8-1:0] node3549;
	wire [8-1:0] node3550;
	wire [8-1:0] node3554;
	wire [8-1:0] node3555;
	wire [8-1:0] node3556;
	wire [8-1:0] node3557;
	wire [8-1:0] node3558;
	wire [8-1:0] node3562;
	wire [8-1:0] node3563;
	wire [8-1:0] node3567;
	wire [8-1:0] node3568;
	wire [8-1:0] node3569;
	wire [8-1:0] node3573;
	wire [8-1:0] node3576;
	wire [8-1:0] node3577;
	wire [8-1:0] node3578;
	wire [8-1:0] node3580;
	wire [8-1:0] node3584;
	wire [8-1:0] node3586;
	wire [8-1:0] node3589;
	wire [8-1:0] node3590;
	wire [8-1:0] node3591;
	wire [8-1:0] node3592;
	wire [8-1:0] node3593;
	wire [8-1:0] node3594;
	wire [8-1:0] node3595;
	wire [8-1:0] node3598;
	wire [8-1:0] node3599;
	wire [8-1:0] node3602;
	wire [8-1:0] node3605;
	wire [8-1:0] node3606;
	wire [8-1:0] node3607;
	wire [8-1:0] node3610;
	wire [8-1:0] node3611;
	wire [8-1:0] node3614;
	wire [8-1:0] node3617;
	wire [8-1:0] node3618;
	wire [8-1:0] node3621;
	wire [8-1:0] node3622;
	wire [8-1:0] node3625;
	wire [8-1:0] node3628;
	wire [8-1:0] node3629;
	wire [8-1:0] node3630;
	wire [8-1:0] node3631;
	wire [8-1:0] node3632;
	wire [8-1:0] node3633;
	wire [8-1:0] node3636;
	wire [8-1:0] node3639;
	wire [8-1:0] node3640;
	wire [8-1:0] node3643;
	wire [8-1:0] node3646;
	wire [8-1:0] node3647;
	wire [8-1:0] node3648;
	wire [8-1:0] node3652;
	wire [8-1:0] node3653;
	wire [8-1:0] node3656;
	wire [8-1:0] node3659;
	wire [8-1:0] node3660;
	wire [8-1:0] node3661;
	wire [8-1:0] node3662;
	wire [8-1:0] node3665;
	wire [8-1:0] node3668;
	wire [8-1:0] node3669;
	wire [8-1:0] node3672;
	wire [8-1:0] node3675;
	wire [8-1:0] node3676;
	wire [8-1:0] node3677;
	wire [8-1:0] node3681;
	wire [8-1:0] node3683;
	wire [8-1:0] node3686;
	wire [8-1:0] node3687;
	wire [8-1:0] node3688;
	wire [8-1:0] node3689;
	wire [8-1:0] node3691;
	wire [8-1:0] node3694;
	wire [8-1:0] node3695;
	wire [8-1:0] node3698;
	wire [8-1:0] node3701;
	wire [8-1:0] node3702;
	wire [8-1:0] node3704;
	wire [8-1:0] node3707;
	wire [8-1:0] node3709;
	wire [8-1:0] node3712;
	wire [8-1:0] node3713;
	wire [8-1:0] node3714;
	wire [8-1:0] node3715;
	wire [8-1:0] node3718;
	wire [8-1:0] node3721;
	wire [8-1:0] node3722;
	wire [8-1:0] node3726;
	wire [8-1:0] node3727;
	wire [8-1:0] node3728;
	wire [8-1:0] node3731;
	wire [8-1:0] node3734;
	wire [8-1:0] node3735;
	wire [8-1:0] node3739;
	wire [8-1:0] node3740;
	wire [8-1:0] node3741;
	wire [8-1:0] node3742;
	wire [8-1:0] node3745;
	wire [8-1:0] node3746;
	wire [8-1:0] node3749;
	wire [8-1:0] node3752;
	wire [8-1:0] node3753;
	wire [8-1:0] node3754;
	wire [8-1:0] node3757;
	wire [8-1:0] node3758;
	wire [8-1:0] node3761;
	wire [8-1:0] node3764;
	wire [8-1:0] node3765;
	wire [8-1:0] node3768;
	wire [8-1:0] node3769;
	wire [8-1:0] node3772;
	wire [8-1:0] node3775;
	wire [8-1:0] node3776;
	wire [8-1:0] node3777;
	wire [8-1:0] node3778;
	wire [8-1:0] node3779;
	wire [8-1:0] node3782;
	wire [8-1:0] node3783;
	wire [8-1:0] node3786;
	wire [8-1:0] node3789;
	wire [8-1:0] node3790;
	wire [8-1:0] node3791;
	wire [8-1:0] node3794;
	wire [8-1:0] node3797;
	wire [8-1:0] node3798;
	wire [8-1:0] node3801;
	wire [8-1:0] node3804;
	wire [8-1:0] node3805;
	wire [8-1:0] node3806;
	wire [8-1:0] node3807;
	wire [8-1:0] node3810;
	wire [8-1:0] node3813;
	wire [8-1:0] node3814;
	wire [8-1:0] node3817;
	wire [8-1:0] node3820;
	wire [8-1:0] node3821;
	wire [8-1:0] node3823;
	wire [8-1:0] node3826;
	wire [8-1:0] node3827;
	wire [8-1:0] node3830;
	wire [8-1:0] node3833;
	wire [8-1:0] node3834;
	wire [8-1:0] node3835;
	wire [8-1:0] node3836;
	wire [8-1:0] node3837;
	wire [8-1:0] node3840;
	wire [8-1:0] node3843;
	wire [8-1:0] node3844;
	wire [8-1:0] node3847;
	wire [8-1:0] node3850;
	wire [8-1:0] node3852;
	wire [8-1:0] node3853;
	wire [8-1:0] node3856;
	wire [8-1:0] node3859;
	wire [8-1:0] node3860;
	wire [8-1:0] node3861;
	wire [8-1:0] node3862;
	wire [8-1:0] node3865;
	wire [8-1:0] node3868;
	wire [8-1:0] node3869;
	wire [8-1:0] node3872;
	wire [8-1:0] node3875;
	wire [8-1:0] node3876;
	wire [8-1:0] node3877;
	wire [8-1:0] node3880;
	wire [8-1:0] node3883;
	wire [8-1:0] node3884;
	wire [8-1:0] node3887;
	wire [8-1:0] node3890;
	wire [8-1:0] node3891;
	wire [8-1:0] node3892;
	wire [8-1:0] node3893;
	wire [8-1:0] node3896;
	wire [8-1:0] node3897;
	wire [8-1:0] node3898;
	wire [8-1:0] node3899;
	wire [8-1:0] node3903;
	wire [8-1:0] node3904;
	wire [8-1:0] node3907;
	wire [8-1:0] node3910;
	wire [8-1:0] node3911;
	wire [8-1:0] node3912;
	wire [8-1:0] node3915;
	wire [8-1:0] node3918;
	wire [8-1:0] node3921;
	wire [8-1:0] node3922;
	wire [8-1:0] node3924;
	wire [8-1:0] node3925;
	wire [8-1:0] node3928;
	wire [8-1:0] node3931;
	wire [8-1:0] node3933;
	wire [8-1:0] node3936;
	wire [8-1:0] node3937;
	wire [8-1:0] node3938;
	wire [8-1:0] node3940;
	wire [8-1:0] node3941;
	wire [8-1:0] node3942;
	wire [8-1:0] node3945;
	wire [8-1:0] node3948;
	wire [8-1:0] node3949;
	wire [8-1:0] node3952;
	wire [8-1:0] node3955;
	wire [8-1:0] node3957;
	wire [8-1:0] node3958;
	wire [8-1:0] node3961;
	wire [8-1:0] node3964;
	wire [8-1:0] node3965;
	wire [8-1:0] node3968;
	wire [8-1:0] node3969;
	wire [8-1:0] node3970;
	wire [8-1:0] node3973;
	wire [8-1:0] node3976;
	wire [8-1:0] node3977;
	wire [8-1:0] node3980;
	wire [8-1:0] node3983;
	wire [8-1:0] node3984;
	wire [8-1:0] node3985;
	wire [8-1:0] node3986;
	wire [8-1:0] node3987;
	wire [8-1:0] node3988;
	wire [8-1:0] node3989;
	wire [8-1:0] node3992;
	wire [8-1:0] node3993;
	wire [8-1:0] node3996;
	wire [8-1:0] node3999;
	wire [8-1:0] node4000;
	wire [8-1:0] node4001;
	wire [8-1:0] node4002;
	wire [8-1:0] node4005;
	wire [8-1:0] node4008;
	wire [8-1:0] node4011;
	wire [8-1:0] node4012;
	wire [8-1:0] node4013;
	wire [8-1:0] node4017;
	wire [8-1:0] node4018;
	wire [8-1:0] node4022;
	wire [8-1:0] node4023;
	wire [8-1:0] node4024;
	wire [8-1:0] node4026;
	wire [8-1:0] node4028;
	wire [8-1:0] node4031;
	wire [8-1:0] node4033;
	wire [8-1:0] node4034;
	wire [8-1:0] node4037;
	wire [8-1:0] node4040;
	wire [8-1:0] node4041;
	wire [8-1:0] node4042;
	wire [8-1:0] node4043;
	wire [8-1:0] node4047;
	wire [8-1:0] node4049;
	wire [8-1:0] node4052;
	wire [8-1:0] node4053;
	wire [8-1:0] node4056;
	wire [8-1:0] node4059;
	wire [8-1:0] node4060;
	wire [8-1:0] node4061;
	wire [8-1:0] node4062;
	wire [8-1:0] node4065;
	wire [8-1:0] node4066;
	wire [8-1:0] node4069;
	wire [8-1:0] node4072;
	wire [8-1:0] node4073;
	wire [8-1:0] node4074;
	wire [8-1:0] node4075;
	wire [8-1:0] node4078;
	wire [8-1:0] node4081;
	wire [8-1:0] node4082;
	wire [8-1:0] node4086;
	wire [8-1:0] node4087;
	wire [8-1:0] node4088;
	wire [8-1:0] node4091;
	wire [8-1:0] node4094;
	wire [8-1:0] node4096;
	wire [8-1:0] node4099;
	wire [8-1:0] node4100;
	wire [8-1:0] node4101;
	wire [8-1:0] node4104;
	wire [8-1:0] node4105;
	wire [8-1:0] node4108;
	wire [8-1:0] node4111;
	wire [8-1:0] node4112;
	wire [8-1:0] node4113;
	wire [8-1:0] node4114;
	wire [8-1:0] node4117;
	wire [8-1:0] node4120;
	wire [8-1:0] node4121;
	wire [8-1:0] node4124;
	wire [8-1:0] node4127;
	wire [8-1:0] node4129;
	wire [8-1:0] node4130;
	wire [8-1:0] node4134;
	wire [8-1:0] node4135;
	wire [8-1:0] node4136;
	wire [8-1:0] node4138;
	wire [8-1:0] node4139;
	wire [8-1:0] node4142;
	wire [8-1:0] node4145;
	wire [8-1:0] node4146;
	wire [8-1:0] node4150;
	wire [8-1:0] node4151;
	wire [8-1:0] node4153;
	wire [8-1:0] node4154;
	wire [8-1:0] node4157;
	wire [8-1:0] node4160;
	wire [8-1:0] node4161;
	wire [8-1:0] node4165;
	wire [8-1:0] node4166;
	wire [8-1:0] node4167;
	wire [8-1:0] node4168;
	wire [8-1:0] node4169;
	wire [8-1:0] node4170;
	wire [8-1:0] node4171;
	wire [8-1:0] node4172;
	wire [8-1:0] node4177;
	wire [8-1:0] node4178;
	wire [8-1:0] node4180;
	wire [8-1:0] node4183;
	wire [8-1:0] node4184;
	wire [8-1:0] node4188;
	wire [8-1:0] node4189;
	wire [8-1:0] node4190;
	wire [8-1:0] node4191;
	wire [8-1:0] node4194;
	wire [8-1:0] node4197;
	wire [8-1:0] node4200;
	wire [8-1:0] node4201;
	wire [8-1:0] node4204;
	wire [8-1:0] node4205;
	wire [8-1:0] node4209;
	wire [8-1:0] node4210;
	wire [8-1:0] node4211;
	wire [8-1:0] node4212;
	wire [8-1:0] node4215;
	wire [8-1:0] node4216;
	wire [8-1:0] node4220;
	wire [8-1:0] node4221;
	wire [8-1:0] node4223;
	wire [8-1:0] node4227;
	wire [8-1:0] node4228;
	wire [8-1:0] node4229;
	wire [8-1:0] node4232;
	wire [8-1:0] node4235;
	wire [8-1:0] node4236;
	wire [8-1:0] node4238;
	wire [8-1:0] node4241;
	wire [8-1:0] node4244;
	wire [8-1:0] node4245;
	wire [8-1:0] node4246;
	wire [8-1:0] node4249;
	wire [8-1:0] node4252;
	wire [8-1:0] node4255;
	wire [8-1:0] node4256;
	wire [8-1:0] node4257;
	wire [8-1:0] node4258;
	wire [8-1:0] node4259;
	wire [8-1:0] node4260;
	wire [8-1:0] node4263;
	wire [8-1:0] node4266;
	wire [8-1:0] node4267;
	wire [8-1:0] node4270;
	wire [8-1:0] node4273;
	wire [8-1:0] node4274;
	wire [8-1:0] node4275;
	wire [8-1:0] node4278;
	wire [8-1:0] node4281;
	wire [8-1:0] node4282;
	wire [8-1:0] node4285;
	wire [8-1:0] node4288;
	wire [8-1:0] node4289;
	wire [8-1:0] node4290;
	wire [8-1:0] node4291;
	wire [8-1:0] node4294;
	wire [8-1:0] node4297;
	wire [8-1:0] node4298;
	wire [8-1:0] node4301;
	wire [8-1:0] node4304;
	wire [8-1:0] node4305;
	wire [8-1:0] node4306;
	wire [8-1:0] node4309;
	wire [8-1:0] node4312;
	wire [8-1:0] node4313;
	wire [8-1:0] node4316;
	wire [8-1:0] node4319;
	wire [8-1:0] node4322;
	wire [8-1:0] node4323;
	wire [8-1:0] node4324;
	wire [8-1:0] node4325;
	wire [8-1:0] node4326;
	wire [8-1:0] node4327;
	wire [8-1:0] node4328;
	wire [8-1:0] node4329;
	wire [8-1:0] node4330;
	wire [8-1:0] node4331;
	wire [8-1:0] node4332;
	wire [8-1:0] node4333;
	wire [8-1:0] node4337;
	wire [8-1:0] node4338;
	wire [8-1:0] node4342;
	wire [8-1:0] node4343;
	wire [8-1:0] node4347;
	wire [8-1:0] node4348;
	wire [8-1:0] node4349;
	wire [8-1:0] node4350;
	wire [8-1:0] node4352;
	wire [8-1:0] node4355;
	wire [8-1:0] node4356;
	wire [8-1:0] node4359;
	wire [8-1:0] node4362;
	wire [8-1:0] node4363;
	wire [8-1:0] node4364;
	wire [8-1:0] node4367;
	wire [8-1:0] node4370;
	wire [8-1:0] node4371;
	wire [8-1:0] node4374;
	wire [8-1:0] node4377;
	wire [8-1:0] node4378;
	wire [8-1:0] node4379;
	wire [8-1:0] node4380;
	wire [8-1:0] node4383;
	wire [8-1:0] node4386;
	wire [8-1:0] node4387;
	wire [8-1:0] node4390;
	wire [8-1:0] node4393;
	wire [8-1:0] node4394;
	wire [8-1:0] node4395;
	wire [8-1:0] node4398;
	wire [8-1:0] node4402;
	wire [8-1:0] node4403;
	wire [8-1:0] node4404;
	wire [8-1:0] node4405;
	wire [8-1:0] node4406;
	wire [8-1:0] node4410;
	wire [8-1:0] node4411;
	wire [8-1:0] node4415;
	wire [8-1:0] node4416;
	wire [8-1:0] node4420;
	wire [8-1:0] node4421;
	wire [8-1:0] node4422;
	wire [8-1:0] node4423;
	wire [8-1:0] node4426;
	wire [8-1:0] node4429;
	wire [8-1:0] node4430;
	wire [8-1:0] node4431;
	wire [8-1:0] node4434;
	wire [8-1:0] node4437;
	wire [8-1:0] node4438;
	wire [8-1:0] node4441;
	wire [8-1:0] node4444;
	wire [8-1:0] node4445;
	wire [8-1:0] node4446;
	wire [8-1:0] node4449;
	wire [8-1:0] node4452;
	wire [8-1:0] node4453;
	wire [8-1:0] node4456;
	wire [8-1:0] node4459;
	wire [8-1:0] node4460;
	wire [8-1:0] node4462;
	wire [8-1:0] node4464;
	wire [8-1:0] node4467;
	wire [8-1:0] node4468;
	wire [8-1:0] node4470;
	wire [8-1:0] node4473;
	wire [8-1:0] node4475;
	wire [8-1:0] node4476;
	wire [8-1:0] node4479;
	wire [8-1:0] node4482;
	wire [8-1:0] node4483;
	wire [8-1:0] node4484;
	wire [8-1:0] node4485;
	wire [8-1:0] node4486;
	wire [8-1:0] node4487;
	wire [8-1:0] node4490;
	wire [8-1:0] node4494;
	wire [8-1:0] node4496;
	wire [8-1:0] node4499;
	wire [8-1:0] node4500;
	wire [8-1:0] node4502;
	wire [8-1:0] node4506;
	wire [8-1:0] node4507;
	wire [8-1:0] node4508;
	wire [8-1:0] node4509;
	wire [8-1:0] node4510;
	wire [8-1:0] node4511;
	wire [8-1:0] node4512;
	wire [8-1:0] node4515;
	wire [8-1:0] node4518;
	wire [8-1:0] node4519;
	wire [8-1:0] node4522;
	wire [8-1:0] node4525;
	wire [8-1:0] node4526;
	wire [8-1:0] node4529;
	wire [8-1:0] node4532;
	wire [8-1:0] node4533;
	wire [8-1:0] node4534;
	wire [8-1:0] node4535;
	wire [8-1:0] node4538;
	wire [8-1:0] node4541;
	wire [8-1:0] node4542;
	wire [8-1:0] node4546;
	wire [8-1:0] node4547;
	wire [8-1:0] node4550;
	wire [8-1:0] node4553;
	wire [8-1:0] node4554;
	wire [8-1:0] node4555;
	wire [8-1:0] node4557;
	wire [8-1:0] node4560;
	wire [8-1:0] node4562;
	wire [8-1:0] node4565;
	wire [8-1:0] node4566;
	wire [8-1:0] node4570;
	wire [8-1:0] node4571;
	wire [8-1:0] node4572;
	wire [8-1:0] node4573;
	wire [8-1:0] node4574;
	wire [8-1:0] node4577;
	wire [8-1:0] node4580;
	wire [8-1:0] node4583;
	wire [8-1:0] node4584;
	wire [8-1:0] node4585;
	wire [8-1:0] node4588;
	wire [8-1:0] node4591;
	wire [8-1:0] node4592;
	wire [8-1:0] node4594;
	wire [8-1:0] node4597;
	wire [8-1:0] node4598;
	wire [8-1:0] node4601;
	wire [8-1:0] node4604;
	wire [8-1:0] node4605;
	wire [8-1:0] node4607;
	wire [8-1:0] node4608;
	wire [8-1:0] node4612;
	wire [8-1:0] node4614;
	wire [8-1:0] node4617;
	wire [8-1:0] node4618;
	wire [8-1:0] node4619;
	wire [8-1:0] node4620;
	wire [8-1:0] node4621;
	wire [8-1:0] node4622;
	wire [8-1:0] node4623;
	wire [8-1:0] node4626;
	wire [8-1:0] node4629;
	wire [8-1:0] node4630;
	wire [8-1:0] node4631;
	wire [8-1:0] node4632;
	wire [8-1:0] node4636;
	wire [8-1:0] node4637;
	wire [8-1:0] node4641;
	wire [8-1:0] node4643;
	wire [8-1:0] node4644;
	wire [8-1:0] node4648;
	wire [8-1:0] node4649;
	wire [8-1:0] node4650;
	wire [8-1:0] node4652;
	wire [8-1:0] node4655;
	wire [8-1:0] node4657;
	wire [8-1:0] node4660;
	wire [8-1:0] node4661;
	wire [8-1:0] node4664;
	wire [8-1:0] node4665;
	wire [8-1:0] node4667;
	wire [8-1:0] node4670;
	wire [8-1:0] node4671;
	wire [8-1:0] node4675;
	wire [8-1:0] node4676;
	wire [8-1:0] node4677;
	wire [8-1:0] node4678;
	wire [8-1:0] node4679;
	wire [8-1:0] node4683;
	wire [8-1:0] node4684;
	wire [8-1:0] node4685;
	wire [8-1:0] node4688;
	wire [8-1:0] node4691;
	wire [8-1:0] node4693;
	wire [8-1:0] node4696;
	wire [8-1:0] node4697;
	wire [8-1:0] node4698;
	wire [8-1:0] node4702;
	wire [8-1:0] node4703;
	wire [8-1:0] node4704;
	wire [8-1:0] node4707;
	wire [8-1:0] node4710;
	wire [8-1:0] node4711;
	wire [8-1:0] node4714;
	wire [8-1:0] node4717;
	wire [8-1:0] node4718;
	wire [8-1:0] node4719;
	wire [8-1:0] node4720;
	wire [8-1:0] node4723;
	wire [8-1:0] node4724;
	wire [8-1:0] node4728;
	wire [8-1:0] node4731;
	wire [8-1:0] node4732;
	wire [8-1:0] node4733;
	wire [8-1:0] node4734;
	wire [8-1:0] node4738;
	wire [8-1:0] node4740;
	wire [8-1:0] node4743;
	wire [8-1:0] node4745;
	wire [8-1:0] node4746;
	wire [8-1:0] node4750;
	wire [8-1:0] node4751;
	wire [8-1:0] node4752;
	wire [8-1:0] node4753;
	wire [8-1:0] node4754;
	wire [8-1:0] node4756;
	wire [8-1:0] node4759;
	wire [8-1:0] node4761;
	wire [8-1:0] node4764;
	wire [8-1:0] node4765;
	wire [8-1:0] node4767;
	wire [8-1:0] node4770;
	wire [8-1:0] node4772;
	wire [8-1:0] node4775;
	wire [8-1:0] node4776;
	wire [8-1:0] node4777;
	wire [8-1:0] node4779;
	wire [8-1:0] node4782;
	wire [8-1:0] node4784;
	wire [8-1:0] node4787;
	wire [8-1:0] node4788;
	wire [8-1:0] node4791;
	wire [8-1:0] node4792;
	wire [8-1:0] node4794;
	wire [8-1:0] node4797;
	wire [8-1:0] node4798;
	wire [8-1:0] node4802;
	wire [8-1:0] node4803;
	wire [8-1:0] node4804;
	wire [8-1:0] node4805;
	wire [8-1:0] node4806;
	wire [8-1:0] node4808;
	wire [8-1:0] node4812;
	wire [8-1:0] node4813;
	wire [8-1:0] node4815;
	wire [8-1:0] node4818;
	wire [8-1:0] node4821;
	wire [8-1:0] node4822;
	wire [8-1:0] node4823;
	wire [8-1:0] node4827;
	wire [8-1:0] node4828;
	wire [8-1:0] node4829;
	wire [8-1:0] node4832;
	wire [8-1:0] node4835;
	wire [8-1:0] node4836;
	wire [8-1:0] node4839;
	wire [8-1:0] node4842;
	wire [8-1:0] node4843;
	wire [8-1:0] node4844;
	wire [8-1:0] node4845;
	wire [8-1:0] node4848;
	wire [8-1:0] node4851;
	wire [8-1:0] node4852;
	wire [8-1:0] node4853;
	wire [8-1:0] node4856;
	wire [8-1:0] node4859;
	wire [8-1:0] node4861;
	wire [8-1:0] node4864;
	wire [8-1:0] node4865;
	wire [8-1:0] node4866;
	wire [8-1:0] node4867;
	wire [8-1:0] node4870;
	wire [8-1:0] node4873;
	wire [8-1:0] node4874;
	wire [8-1:0] node4878;
	wire [8-1:0] node4881;
	wire [8-1:0] node4882;
	wire [8-1:0] node4883;
	wire [8-1:0] node4884;
	wire [8-1:0] node4885;
	wire [8-1:0] node4886;
	wire [8-1:0] node4887;
	wire [8-1:0] node4891;
	wire [8-1:0] node4892;
	wire [8-1:0] node4894;
	wire [8-1:0] node4897;
	wire [8-1:0] node4900;
	wire [8-1:0] node4901;
	wire [8-1:0] node4902;
	wire [8-1:0] node4905;
	wire [8-1:0] node4906;
	wire [8-1:0] node4909;
	wire [8-1:0] node4912;
	wire [8-1:0] node4914;
	wire [8-1:0] node4917;
	wire [8-1:0] node4918;
	wire [8-1:0] node4919;
	wire [8-1:0] node4921;
	wire [8-1:0] node4924;
	wire [8-1:0] node4926;
	wire [8-1:0] node4929;
	wire [8-1:0] node4931;
	wire [8-1:0] node4934;
	wire [8-1:0] node4935;
	wire [8-1:0] node4936;
	wire [8-1:0] node4937;
	wire [8-1:0] node4938;
	wire [8-1:0] node4942;
	wire [8-1:0] node4945;
	wire [8-1:0] node4946;
	wire [8-1:0] node4950;
	wire [8-1:0] node4951;
	wire [8-1:0] node4952;
	wire [8-1:0] node4953;
	wire [8-1:0] node4954;
	wire [8-1:0] node4957;
	wire [8-1:0] node4960;
	wire [8-1:0] node4961;
	wire [8-1:0] node4965;
	wire [8-1:0] node4966;
	wire [8-1:0] node4967;
	wire [8-1:0] node4971;
	wire [8-1:0] node4972;
	wire [8-1:0] node4976;
	wire [8-1:0] node4977;
	wire [8-1:0] node4978;
	wire [8-1:0] node4981;
	wire [8-1:0] node4984;
	wire [8-1:0] node4987;
	wire [8-1:0] node4988;
	wire [8-1:0] node4989;
	wire [8-1:0] node4990;
	wire [8-1:0] node4991;
	wire [8-1:0] node4992;
	wire [8-1:0] node4994;
	wire [8-1:0] node4997;
	wire [8-1:0] node4998;
	wire [8-1:0] node5001;
	wire [8-1:0] node5004;
	wire [8-1:0] node5005;
	wire [8-1:0] node5006;
	wire [8-1:0] node5009;
	wire [8-1:0] node5012;
	wire [8-1:0] node5013;
	wire [8-1:0] node5016;
	wire [8-1:0] node5019;
	wire [8-1:0] node5020;
	wire [8-1:0] node5021;
	wire [8-1:0] node5022;
	wire [8-1:0] node5026;
	wire [8-1:0] node5027;
	wire [8-1:0] node5031;
	wire [8-1:0] node5032;
	wire [8-1:0] node5033;
	wire [8-1:0] node5036;
	wire [8-1:0] node5040;
	wire [8-1:0] node5041;
	wire [8-1:0] node5042;
	wire [8-1:0] node5043;
	wire [8-1:0] node5046;
	wire [8-1:0] node5049;
	wire [8-1:0] node5050;
	wire [8-1:0] node5051;
	wire [8-1:0] node5055;
	wire [8-1:0] node5056;
	wire [8-1:0] node5060;
	wire [8-1:0] node5061;
	wire [8-1:0] node5062;
	wire [8-1:0] node5065;
	wire [8-1:0] node5068;
	wire [8-1:0] node5070;
	wire [8-1:0] node5071;
	wire [8-1:0] node5075;
	wire [8-1:0] node5076;
	wire [8-1:0] node5077;
	wire [8-1:0] node5078;
	wire [8-1:0] node5079;
	wire [8-1:0] node5081;
	wire [8-1:0] node5084;
	wire [8-1:0] node5085;
	wire [8-1:0] node5088;
	wire [8-1:0] node5091;
	wire [8-1:0] node5092;
	wire [8-1:0] node5093;
	wire [8-1:0] node5096;
	wire [8-1:0] node5099;
	wire [8-1:0] node5100;
	wire [8-1:0] node5103;
	wire [8-1:0] node5106;
	wire [8-1:0] node5107;
	wire [8-1:0] node5108;
	wire [8-1:0] node5110;
	wire [8-1:0] node5113;
	wire [8-1:0] node5115;
	wire [8-1:0] node5118;
	wire [8-1:0] node5119;
	wire [8-1:0] node5120;
	wire [8-1:0] node5123;
	wire [8-1:0] node5126;
	wire [8-1:0] node5127;
	wire [8-1:0] node5130;
	wire [8-1:0] node5133;
	wire [8-1:0] node5134;
	wire [8-1:0] node5135;
	wire [8-1:0] node5138;
	wire [8-1:0] node5141;
	wire [8-1:0] node5144;
	wire [8-1:0] node5145;
	wire [8-1:0] node5146;
	wire [8-1:0] node5147;
	wire [8-1:0] node5148;
	wire [8-1:0] node5149;
	wire [8-1:0] node5150;
	wire [8-1:0] node5151;
	wire [8-1:0] node5152;
	wire [8-1:0] node5156;
	wire [8-1:0] node5157;
	wire [8-1:0] node5160;
	wire [8-1:0] node5163;
	wire [8-1:0] node5164;
	wire [8-1:0] node5165;
	wire [8-1:0] node5169;
	wire [8-1:0] node5171;
	wire [8-1:0] node5172;
	wire [8-1:0] node5176;
	wire [8-1:0] node5178;
	wire [8-1:0] node5180;
	wire [8-1:0] node5183;
	wire [8-1:0] node5184;
	wire [8-1:0] node5185;
	wire [8-1:0] node5186;
	wire [8-1:0] node5188;
	wire [8-1:0] node5191;
	wire [8-1:0] node5193;
	wire [8-1:0] node5196;
	wire [8-1:0] node5198;
	wire [8-1:0] node5201;
	wire [8-1:0] node5203;
	wire [8-1:0] node5204;
	wire [8-1:0] node5207;
	wire [8-1:0] node5210;
	wire [8-1:0] node5211;
	wire [8-1:0] node5212;
	wire [8-1:0] node5213;
	wire [8-1:0] node5214;
	wire [8-1:0] node5217;
	wire [8-1:0] node5220;
	wire [8-1:0] node5221;
	wire [8-1:0] node5222;
	wire [8-1:0] node5224;
	wire [8-1:0] node5227;
	wire [8-1:0] node5229;
	wire [8-1:0] node5232;
	wire [8-1:0] node5233;
	wire [8-1:0] node5234;
	wire [8-1:0] node5238;
	wire [8-1:0] node5239;
	wire [8-1:0] node5243;
	wire [8-1:0] node5244;
	wire [8-1:0] node5245;
	wire [8-1:0] node5248;
	wire [8-1:0] node5251;
	wire [8-1:0] node5252;
	wire [8-1:0] node5254;
	wire [8-1:0] node5255;
	wire [8-1:0] node5259;
	wire [8-1:0] node5260;
	wire [8-1:0] node5261;
	wire [8-1:0] node5265;
	wire [8-1:0] node5266;
	wire [8-1:0] node5270;
	wire [8-1:0] node5271;
	wire [8-1:0] node5272;
	wire [8-1:0] node5273;
	wire [8-1:0] node5274;
	wire [8-1:0] node5276;
	wire [8-1:0] node5280;
	wire [8-1:0] node5281;
	wire [8-1:0] node5283;
	wire [8-1:0] node5286;
	wire [8-1:0] node5288;
	wire [8-1:0] node5291;
	wire [8-1:0] node5292;
	wire [8-1:0] node5293;
	wire [8-1:0] node5294;
	wire [8-1:0] node5297;
	wire [8-1:0] node5300;
	wire [8-1:0] node5301;
	wire [8-1:0] node5305;
	wire [8-1:0] node5307;
	wire [8-1:0] node5310;
	wire [8-1:0] node5311;
	wire [8-1:0] node5312;
	wire [8-1:0] node5313;
	wire [8-1:0] node5315;
	wire [8-1:0] node5318;
	wire [8-1:0] node5320;
	wire [8-1:0] node5323;
	wire [8-1:0] node5325;
	wire [8-1:0] node5326;
	wire [8-1:0] node5329;
	wire [8-1:0] node5332;
	wire [8-1:0] node5333;
	wire [8-1:0] node5334;
	wire [8-1:0] node5335;
	wire [8-1:0] node5340;
	wire [8-1:0] node5341;
	wire [8-1:0] node5342;
	wire [8-1:0] node5347;
	wire [8-1:0] node5348;
	wire [8-1:0] node5349;
	wire [8-1:0] node5350;
	wire [8-1:0] node5351;
	wire [8-1:0] node5353;
	wire [8-1:0] node5356;
	wire [8-1:0] node5358;
	wire [8-1:0] node5361;
	wire [8-1:0] node5362;
	wire [8-1:0] node5363;
	wire [8-1:0] node5365;
	wire [8-1:0] node5368;
	wire [8-1:0] node5370;
	wire [8-1:0] node5373;
	wire [8-1:0] node5374;
	wire [8-1:0] node5376;
	wire [8-1:0] node5379;
	wire [8-1:0] node5381;
	wire [8-1:0] node5384;
	wire [8-1:0] node5385;
	wire [8-1:0] node5386;
	wire [8-1:0] node5388;
	wire [8-1:0] node5391;
	wire [8-1:0] node5392;
	wire [8-1:0] node5393;
	wire [8-1:0] node5396;
	wire [8-1:0] node5397;
	wire [8-1:0] node5401;
	wire [8-1:0] node5403;
	wire [8-1:0] node5404;
	wire [8-1:0] node5408;
	wire [8-1:0] node5409;
	wire [8-1:0] node5410;
	wire [8-1:0] node5413;
	wire [8-1:0] node5416;
	wire [8-1:0] node5417;
	wire [8-1:0] node5418;
	wire [8-1:0] node5420;
	wire [8-1:0] node5423;
	wire [8-1:0] node5424;
	wire [8-1:0] node5428;
	wire [8-1:0] node5429;
	wire [8-1:0] node5431;
	wire [8-1:0] node5435;
	wire [8-1:0] node5436;
	wire [8-1:0] node5437;
	wire [8-1:0] node5438;
	wire [8-1:0] node5439;
	wire [8-1:0] node5440;
	wire [8-1:0] node5444;
	wire [8-1:0] node5445;
	wire [8-1:0] node5448;
	wire [8-1:0] node5451;
	wire [8-1:0] node5452;
	wire [8-1:0] node5455;
	wire [8-1:0] node5458;
	wire [8-1:0] node5459;
	wire [8-1:0] node5460;
	wire [8-1:0] node5461;
	wire [8-1:0] node5463;
	wire [8-1:0] node5466;
	wire [8-1:0] node5469;
	wire [8-1:0] node5470;
	wire [8-1:0] node5473;
	wire [8-1:0] node5476;
	wire [8-1:0] node5477;
	wire [8-1:0] node5481;
	wire [8-1:0] node5482;
	wire [8-1:0] node5483;
	wire [8-1:0] node5484;
	wire [8-1:0] node5485;
	wire [8-1:0] node5487;
	wire [8-1:0] node5490;
	wire [8-1:0] node5492;
	wire [8-1:0] node5495;
	wire [8-1:0] node5496;
	wire [8-1:0] node5500;
	wire [8-1:0] node5501;
	wire [8-1:0] node5502;
	wire [8-1:0] node5506;
	wire [8-1:0] node5507;
	wire [8-1:0] node5509;
	wire [8-1:0] node5512;
	wire [8-1:0] node5515;
	wire [8-1:0] node5516;
	wire [8-1:0] node5517;
	wire [8-1:0] node5519;
	wire [8-1:0] node5520;
	wire [8-1:0] node5524;
	wire [8-1:0] node5525;
	wire [8-1:0] node5526;
	wire [8-1:0] node5531;
	wire [8-1:0] node5532;
	wire [8-1:0] node5533;
	wire [8-1:0] node5535;
	wire [8-1:0] node5539;
	wire [8-1:0] node5540;
	wire [8-1:0] node5542;
	wire [8-1:0] node5545;
	wire [8-1:0] node5546;
	wire [8-1:0] node5550;
	wire [8-1:0] node5551;
	wire [8-1:0] node5552;
	wire [8-1:0] node5553;
	wire [8-1:0] node5554;
	wire [8-1:0] node5555;
	wire [8-1:0] node5556;
	wire [8-1:0] node5557;
	wire [8-1:0] node5561;
	wire [8-1:0] node5562;
	wire [8-1:0] node5566;
	wire [8-1:0] node5567;
	wire [8-1:0] node5571;
	wire [8-1:0] node5572;
	wire [8-1:0] node5573;
	wire [8-1:0] node5574;
	wire [8-1:0] node5578;
	wire [8-1:0] node5579;
	wire [8-1:0] node5583;
	wire [8-1:0] node5584;
	wire [8-1:0] node5588;
	wire [8-1:0] node5589;
	wire [8-1:0] node5590;
	wire [8-1:0] node5591;
	wire [8-1:0] node5595;
	wire [8-1:0] node5596;
	wire [8-1:0] node5600;
	wire [8-1:0] node5601;
	wire [8-1:0] node5605;
	wire [8-1:0] node5606;
	wire [8-1:0] node5607;
	wire [8-1:0] node5608;
	wire [8-1:0] node5609;
	wire [8-1:0] node5611;
	wire [8-1:0] node5614;
	wire [8-1:0] node5617;
	wire [8-1:0] node5618;
	wire [8-1:0] node5622;
	wire [8-1:0] node5623;
	wire [8-1:0] node5624;
	wire [8-1:0] node5625;
	wire [8-1:0] node5628;
	wire [8-1:0] node5631;
	wire [8-1:0] node5632;
	wire [8-1:0] node5633;
	wire [8-1:0] node5637;
	wire [8-1:0] node5638;
	wire [8-1:0] node5642;
	wire [8-1:0] node5643;
	wire [8-1:0] node5644;
	wire [8-1:0] node5645;
	wire [8-1:0] node5648;
	wire [8-1:0] node5651;
	wire [8-1:0] node5653;
	wire [8-1:0] node5656;
	wire [8-1:0] node5657;
	wire [8-1:0] node5660;
	wire [8-1:0] node5663;
	wire [8-1:0] node5664;
	wire [8-1:0] node5665;
	wire [8-1:0] node5666;
	wire [8-1:0] node5668;
	wire [8-1:0] node5669;
	wire [8-1:0] node5672;
	wire [8-1:0] node5675;
	wire [8-1:0] node5676;
	wire [8-1:0] node5680;
	wire [8-1:0] node5681;
	wire [8-1:0] node5682;
	wire [8-1:0] node5683;
	wire [8-1:0] node5687;
	wire [8-1:0] node5688;
	wire [8-1:0] node5692;
	wire [8-1:0] node5693;
	wire [8-1:0] node5695;
	wire [8-1:0] node5698;
	wire [8-1:0] node5699;
	wire [8-1:0] node5702;
	wire [8-1:0] node5705;
	wire [8-1:0] node5706;
	wire [8-1:0] node5707;
	wire [8-1:0] node5708;
	wire [8-1:0] node5712;
	wire [8-1:0] node5713;
	wire [8-1:0] node5716;
	wire [8-1:0] node5717;
	wire [8-1:0] node5720;
	wire [8-1:0] node5723;
	wire [8-1:0] node5724;
	wire [8-1:0] node5725;
	wire [8-1:0] node5726;
	wire [8-1:0] node5730;
	wire [8-1:0] node5733;
	wire [8-1:0] node5734;
	wire [8-1:0] node5736;
	wire [8-1:0] node5739;
	wire [8-1:0] node5740;
	wire [8-1:0] node5744;
	wire [8-1:0] node5745;
	wire [8-1:0] node5746;
	wire [8-1:0] node5747;
	wire [8-1:0] node5748;
	wire [8-1:0] node5749;
	wire [8-1:0] node5750;
	wire [8-1:0] node5752;
	wire [8-1:0] node5755;
	wire [8-1:0] node5756;
	wire [8-1:0] node5759;
	wire [8-1:0] node5762;
	wire [8-1:0] node5763;
	wire [8-1:0] node5765;
	wire [8-1:0] node5768;
	wire [8-1:0] node5771;
	wire [8-1:0] node5772;
	wire [8-1:0] node5773;
	wire [8-1:0] node5775;
	wire [8-1:0] node5778;
	wire [8-1:0] node5781;
	wire [8-1:0] node5782;
	wire [8-1:0] node5785;
	wire [8-1:0] node5788;
	wire [8-1:0] node5789;
	wire [8-1:0] node5790;
	wire [8-1:0] node5791;
	wire [8-1:0] node5794;
	wire [8-1:0] node5797;
	wire [8-1:0] node5798;
	wire [8-1:0] node5801;
	wire [8-1:0] node5804;
	wire [8-1:0] node5805;
	wire [8-1:0] node5806;
	wire [8-1:0] node5809;
	wire [8-1:0] node5812;
	wire [8-1:0] node5813;
	wire [8-1:0] node5815;
	wire [8-1:0] node5818;
	wire [8-1:0] node5820;
	wire [8-1:0] node5823;
	wire [8-1:0] node5824;
	wire [8-1:0] node5825;
	wire [8-1:0] node5827;
	wire [8-1:0] node5830;
	wire [8-1:0] node5831;
	wire [8-1:0] node5834;
	wire [8-1:0] node5837;
	wire [8-1:0] node5838;
	wire [8-1:0] node5839;
	wire [8-1:0] node5842;
	wire [8-1:0] node5845;
	wire [8-1:0] node5846;
	wire [8-1:0] node5849;
	wire [8-1:0] node5852;
	wire [8-1:0] node5853;
	wire [8-1:0] node5854;
	wire [8-1:0] node5855;
	wire [8-1:0] node5856;
	wire [8-1:0] node5857;
	wire [8-1:0] node5860;
	wire [8-1:0] node5861;
	wire [8-1:0] node5864;
	wire [8-1:0] node5867;
	wire [8-1:0] node5868;
	wire [8-1:0] node5870;
	wire [8-1:0] node5873;
	wire [8-1:0] node5874;
	wire [8-1:0] node5877;
	wire [8-1:0] node5880;
	wire [8-1:0] node5881;
	wire [8-1:0] node5882;
	wire [8-1:0] node5885;
	wire [8-1:0] node5888;
	wire [8-1:0] node5891;
	wire [8-1:0] node5892;
	wire [8-1:0] node5893;
	wire [8-1:0] node5894;
	wire [8-1:0] node5895;
	wire [8-1:0] node5898;
	wire [8-1:0] node5901;
	wire [8-1:0] node5904;
	wire [8-1:0] node5906;
	wire [8-1:0] node5907;
	wire [8-1:0] node5911;
	wire [8-1:0] node5912;
	wire [8-1:0] node5913;
	wire [8-1:0] node5916;
	wire [8-1:0] node5918;
	wire [8-1:0] node5921;
	wire [8-1:0] node5924;
	wire [8-1:0] node5925;
	wire [8-1:0] node5926;
	wire [8-1:0] node5927;
	wire [8-1:0] node5928;
	wire [8-1:0] node5929;
	wire [8-1:0] node5932;
	wire [8-1:0] node5936;
	wire [8-1:0] node5937;
	wire [8-1:0] node5939;
	wire [8-1:0] node5943;
	wire [8-1:0] node5944;
	wire [8-1:0] node5945;
	wire [8-1:0] node5947;
	wire [8-1:0] node5951;
	wire [8-1:0] node5952;
	wire [8-1:0] node5954;
	wire [8-1:0] node5958;
	wire [8-1:0] node5959;
	wire [8-1:0] node5960;
	wire [8-1:0] node5961;
	wire [8-1:0] node5963;
	wire [8-1:0] node5966;
	wire [8-1:0] node5967;
	wire [8-1:0] node5971;
	wire [8-1:0] node5972;
	wire [8-1:0] node5973;
	wire [8-1:0] node5976;
	wire [8-1:0] node5979;
	wire [8-1:0] node5980;
	wire [8-1:0] node5983;
	wire [8-1:0] node5986;
	wire [8-1:0] node5989;
	wire [8-1:0] node5990;
	wire [8-1:0] node5991;
	wire [8-1:0] node5992;
	wire [8-1:0] node5993;
	wire [8-1:0] node5994;
	wire [8-1:0] node5995;
	wire [8-1:0] node5996;
	wire [8-1:0] node5997;
	wire [8-1:0] node5998;
	wire [8-1:0] node6002;
	wire [8-1:0] node6003;
	wire [8-1:0] node6007;
	wire [8-1:0] node6008;
	wire [8-1:0] node6012;
	wire [8-1:0] node6013;
	wire [8-1:0] node6014;
	wire [8-1:0] node6015;
	wire [8-1:0] node6019;
	wire [8-1:0] node6020;
	wire [8-1:0] node6024;
	wire [8-1:0] node6025;
	wire [8-1:0] node6029;
	wire [8-1:0] node6030;
	wire [8-1:0] node6031;
	wire [8-1:0] node6032;
	wire [8-1:0] node6036;
	wire [8-1:0] node6037;
	wire [8-1:0] node6041;
	wire [8-1:0] node6042;
	wire [8-1:0] node6046;
	wire [8-1:0] node6047;
	wire [8-1:0] node6048;
	wire [8-1:0] node6049;
	wire [8-1:0] node6050;
	wire [8-1:0] node6051;
	wire [8-1:0] node6055;
	wire [8-1:0] node6056;
	wire [8-1:0] node6060;
	wire [8-1:0] node6061;
	wire [8-1:0] node6065;
	wire [8-1:0] node6066;
	wire [8-1:0] node6067;
	wire [8-1:0] node6068;
	wire [8-1:0] node6072;
	wire [8-1:0] node6073;
	wire [8-1:0] node6077;
	wire [8-1:0] node6078;
	wire [8-1:0] node6082;
	wire [8-1:0] node6083;
	wire [8-1:0] node6084;
	wire [8-1:0] node6085;
	wire [8-1:0] node6089;
	wire [8-1:0] node6090;
	wire [8-1:0] node6094;
	wire [8-1:0] node6095;
	wire [8-1:0] node6099;
	wire [8-1:0] node6100;
	wire [8-1:0] node6101;
	wire [8-1:0] node6102;
	wire [8-1:0] node6103;
	wire [8-1:0] node6104;
	wire [8-1:0] node6108;
	wire [8-1:0] node6109;
	wire [8-1:0] node6113;
	wire [8-1:0] node6114;
	wire [8-1:0] node6118;
	wire [8-1:0] node6119;
	wire [8-1:0] node6120;
	wire [8-1:0] node6121;
	wire [8-1:0] node6125;
	wire [8-1:0] node6126;
	wire [8-1:0] node6130;
	wire [8-1:0] node6131;
	wire [8-1:0] node6135;
	wire [8-1:0] node6136;
	wire [8-1:0] node6137;
	wire [8-1:0] node6138;
	wire [8-1:0] node6142;
	wire [8-1:0] node6143;
	wire [8-1:0] node6147;
	wire [8-1:0] node6148;
	wire [8-1:0] node6152;
	wire [8-1:0] node6153;
	wire [8-1:0] node6154;
	wire [8-1:0] node6155;
	wire [8-1:0] node6156;
	wire [8-1:0] node6157;
	wire [8-1:0] node6159;
	wire [8-1:0] node6161;
	wire [8-1:0] node6164;
	wire [8-1:0] node6166;
	wire [8-1:0] node6169;
	wire [8-1:0] node6170;
	wire [8-1:0] node6172;
	wire [8-1:0] node6175;
	wire [8-1:0] node6178;
	wire [8-1:0] node6179;
	wire [8-1:0] node6180;
	wire [8-1:0] node6181;
	wire [8-1:0] node6182;
	wire [8-1:0] node6184;
	wire [8-1:0] node6187;
	wire [8-1:0] node6188;
	wire [8-1:0] node6191;
	wire [8-1:0] node6194;
	wire [8-1:0] node6195;
	wire [8-1:0] node6196;
	wire [8-1:0] node6199;
	wire [8-1:0] node6202;
	wire [8-1:0] node6203;
	wire [8-1:0] node6206;
	wire [8-1:0] node6209;
	wire [8-1:0] node6210;
	wire [8-1:0] node6211;
	wire [8-1:0] node6215;
	wire [8-1:0] node6216;
	wire [8-1:0] node6220;
	wire [8-1:0] node6221;
	wire [8-1:0] node6222;
	wire [8-1:0] node6223;
	wire [8-1:0] node6224;
	wire [8-1:0] node6228;
	wire [8-1:0] node6229;
	wire [8-1:0] node6232;
	wire [8-1:0] node6235;
	wire [8-1:0] node6236;
	wire [8-1:0] node6238;
	wire [8-1:0] node6241;
	wire [8-1:0] node6242;
	wire [8-1:0] node6245;
	wire [8-1:0] node6248;
	wire [8-1:0] node6249;
	wire [8-1:0] node6250;
	wire [8-1:0] node6253;
	wire [8-1:0] node6256;
	wire [8-1:0] node6257;
	wire [8-1:0] node6260;
	wire [8-1:0] node6263;
	wire [8-1:0] node6264;
	wire [8-1:0] node6265;
	wire [8-1:0] node6266;
	wire [8-1:0] node6268;
	wire [8-1:0] node6271;
	wire [8-1:0] node6274;
	wire [8-1:0] node6275;
	wire [8-1:0] node6279;
	wire [8-1:0] node6280;
	wire [8-1:0] node6281;
	wire [8-1:0] node6282;
	wire [8-1:0] node6283;
	wire [8-1:0] node6286;
	wire [8-1:0] node6289;
	wire [8-1:0] node6292;
	wire [8-1:0] node6293;
	wire [8-1:0] node6296;
	wire [8-1:0] node6297;
	wire [8-1:0] node6301;
	wire [8-1:0] node6302;
	wire [8-1:0] node6303;
	wire [8-1:0] node6304;
	wire [8-1:0] node6307;
	wire [8-1:0] node6310;
	wire [8-1:0] node6311;
	wire [8-1:0] node6314;
	wire [8-1:0] node6317;
	wire [8-1:0] node6318;
	wire [8-1:0] node6321;
	wire [8-1:0] node6324;
	wire [8-1:0] node6325;
	wire [8-1:0] node6326;
	wire [8-1:0] node6327;
	wire [8-1:0] node6328;
	wire [8-1:0] node6331;
	wire [8-1:0] node6332;
	wire [8-1:0] node6333;
	wire [8-1:0] node6334;
	wire [8-1:0] node6337;
	wire [8-1:0] node6340;
	wire [8-1:0] node6341;
	wire [8-1:0] node6345;
	wire [8-1:0] node6346;
	wire [8-1:0] node6347;
	wire [8-1:0] node6350;
	wire [8-1:0] node6353;
	wire [8-1:0] node6354;
	wire [8-1:0] node6357;
	wire [8-1:0] node6360;
	wire [8-1:0] node6361;
	wire [8-1:0] node6364;
	wire [8-1:0] node6365;
	wire [8-1:0] node6366;
	wire [8-1:0] node6370;
	wire [8-1:0] node6371;
	wire [8-1:0] node6375;
	wire [8-1:0] node6376;
	wire [8-1:0] node6377;
	wire [8-1:0] node6378;
	wire [8-1:0] node6379;
	wire [8-1:0] node6383;
	wire [8-1:0] node6386;
	wire [8-1:0] node6387;
	wire [8-1:0] node6390;
	wire [8-1:0] node6393;
	wire [8-1:0] node6394;
	wire [8-1:0] node6395;
	wire [8-1:0] node6396;
	wire [8-1:0] node6398;
	wire [8-1:0] node6401;
	wire [8-1:0] node6402;
	wire [8-1:0] node6406;
	wire [8-1:0] node6407;
	wire [8-1:0] node6410;
	wire [8-1:0] node6413;
	wire [8-1:0] node6414;
	wire [8-1:0] node6415;
	wire [8-1:0] node6416;
	wire [8-1:0] node6419;
	wire [8-1:0] node6422;
	wire [8-1:0] node6423;
	wire [8-1:0] node6426;
	wire [8-1:0] node6429;
	wire [8-1:0] node6430;
	wire [8-1:0] node6431;
	wire [8-1:0] node6434;
	wire [8-1:0] node6437;
	wire [8-1:0] node6438;
	wire [8-1:0] node6441;
	wire [8-1:0] node6444;
	wire [8-1:0] node6445;
	wire [8-1:0] node6446;
	wire [8-1:0] node6447;
	wire [8-1:0] node6448;
	wire [8-1:0] node6451;
	wire [8-1:0] node6454;
	wire [8-1:0] node6455;
	wire [8-1:0] node6459;
	wire [8-1:0] node6460;
	wire [8-1:0] node6461;
	wire [8-1:0] node6462;
	wire [8-1:0] node6463;
	wire [8-1:0] node6466;
	wire [8-1:0] node6469;
	wire [8-1:0] node6471;
	wire [8-1:0] node6474;
	wire [8-1:0] node6475;
	wire [8-1:0] node6476;
	wire [8-1:0] node6479;
	wire [8-1:0] node6482;
	wire [8-1:0] node6483;
	wire [8-1:0] node6486;
	wire [8-1:0] node6489;
	wire [8-1:0] node6490;
	wire [8-1:0] node6491;
	wire [8-1:0] node6492;
	wire [8-1:0] node6495;
	wire [8-1:0] node6498;
	wire [8-1:0] node6499;
	wire [8-1:0] node6502;
	wire [8-1:0] node6505;
	wire [8-1:0] node6506;
	wire [8-1:0] node6507;
	wire [8-1:0] node6510;
	wire [8-1:0] node6513;
	wire [8-1:0] node6515;
	wire [8-1:0] node6518;
	wire [8-1:0] node6519;
	wire [8-1:0] node6520;
	wire [8-1:0] node6521;
	wire [8-1:0] node6524;
	wire [8-1:0] node6525;
	wire [8-1:0] node6526;
	wire [8-1:0] node6529;
	wire [8-1:0] node6532;
	wire [8-1:0] node6533;
	wire [8-1:0] node6536;
	wire [8-1:0] node6539;
	wire [8-1:0] node6540;
	wire [8-1:0] node6541;
	wire [8-1:0] node6544;
	wire [8-1:0] node6547;
	wire [8-1:0] node6548;
	wire [8-1:0] node6551;
	wire [8-1:0] node6554;
	wire [8-1:0] node6555;
	wire [8-1:0] node6556;
	wire [8-1:0] node6557;
	wire [8-1:0] node6561;
	wire [8-1:0] node6562;
	wire [8-1:0] node6563;
	wire [8-1:0] node6566;
	wire [8-1:0] node6569;
	wire [8-1:0] node6570;
	wire [8-1:0] node6573;
	wire [8-1:0] node6576;
	wire [8-1:0] node6577;
	wire [8-1:0] node6578;
	wire [8-1:0] node6579;
	wire [8-1:0] node6583;
	wire [8-1:0] node6584;
	wire [8-1:0] node6588;
	wire [8-1:0] node6589;
	wire [8-1:0] node6591;
	wire [8-1:0] node6594;
	wire [8-1:0] node6595;
	wire [8-1:0] node6598;
	wire [8-1:0] node6601;
	wire [8-1:0] node6602;
	wire [8-1:0] node6603;
	wire [8-1:0] node6604;
	wire [8-1:0] node6605;
	wire [8-1:0] node6606;
	wire [8-1:0] node6607;
	wire [8-1:0] node6608;
	wire [8-1:0] node6609;
	wire [8-1:0] node6612;
	wire [8-1:0] node6615;
	wire [8-1:0] node6618;
	wire [8-1:0] node6619;
	wire [8-1:0] node6620;
	wire [8-1:0] node6622;
	wire [8-1:0] node6625;
	wire [8-1:0] node6626;
	wire [8-1:0] node6629;
	wire [8-1:0] node6632;
	wire [8-1:0] node6634;
	wire [8-1:0] node6637;
	wire [8-1:0] node6638;
	wire [8-1:0] node6639;
	wire [8-1:0] node6640;
	wire [8-1:0] node6643;
	wire [8-1:0] node6646;
	wire [8-1:0] node6648;
	wire [8-1:0] node6649;
	wire [8-1:0] node6652;
	wire [8-1:0] node6655;
	wire [8-1:0] node6656;
	wire [8-1:0] node6657;
	wire [8-1:0] node6659;
	wire [8-1:0] node6662;
	wire [8-1:0] node6665;
	wire [8-1:0] node6666;
	wire [8-1:0] node6669;
	wire [8-1:0] node6672;
	wire [8-1:0] node6673;
	wire [8-1:0] node6674;
	wire [8-1:0] node6675;
	wire [8-1:0] node6676;
	wire [8-1:0] node6679;
	wire [8-1:0] node6682;
	wire [8-1:0] node6683;
	wire [8-1:0] node6685;
	wire [8-1:0] node6688;
	wire [8-1:0] node6689;
	wire [8-1:0] node6693;
	wire [8-1:0] node6694;
	wire [8-1:0] node6695;
	wire [8-1:0] node6697;
	wire [8-1:0] node6700;
	wire [8-1:0] node6703;
	wire [8-1:0] node6704;
	wire [8-1:0] node6707;
	wire [8-1:0] node6710;
	wire [8-1:0] node6711;
	wire [8-1:0] node6712;
	wire [8-1:0] node6713;
	wire [8-1:0] node6716;
	wire [8-1:0] node6719;
	wire [8-1:0] node6720;
	wire [8-1:0] node6723;
	wire [8-1:0] node6726;
	wire [8-1:0] node6727;
	wire [8-1:0] node6728;
	wire [8-1:0] node6731;
	wire [8-1:0] node6734;
	wire [8-1:0] node6735;
	wire [8-1:0] node6736;
	wire [8-1:0] node6739;
	wire [8-1:0] node6743;
	wire [8-1:0] node6744;
	wire [8-1:0] node6745;
	wire [8-1:0] node6746;
	wire [8-1:0] node6747;
	wire [8-1:0] node6749;
	wire [8-1:0] node6750;
	wire [8-1:0] node6753;
	wire [8-1:0] node6756;
	wire [8-1:0] node6757;
	wire [8-1:0] node6758;
	wire [8-1:0] node6761;
	wire [8-1:0] node6764;
	wire [8-1:0] node6765;
	wire [8-1:0] node6768;
	wire [8-1:0] node6771;
	wire [8-1:0] node6772;
	wire [8-1:0] node6773;
	wire [8-1:0] node6774;
	wire [8-1:0] node6778;
	wire [8-1:0] node6779;
	wire [8-1:0] node6782;
	wire [8-1:0] node6785;
	wire [8-1:0] node6786;
	wire [8-1:0] node6787;
	wire [8-1:0] node6790;
	wire [8-1:0] node6793;
	wire [8-1:0] node6794;
	wire [8-1:0] node6797;
	wire [8-1:0] node6800;
	wire [8-1:0] node6801;
	wire [8-1:0] node6802;
	wire [8-1:0] node6803;
	wire [8-1:0] node6806;
	wire [8-1:0] node6809;
	wire [8-1:0] node6810;
	wire [8-1:0] node6813;
	wire [8-1:0] node6816;
	wire [8-1:0] node6817;
	wire [8-1:0] node6818;
	wire [8-1:0] node6821;
	wire [8-1:0] node6824;
	wire [8-1:0] node6825;
	wire [8-1:0] node6828;
	wire [8-1:0] node6831;
	wire [8-1:0] node6832;
	wire [8-1:0] node6833;
	wire [8-1:0] node6834;
	wire [8-1:0] node6835;
	wire [8-1:0] node6838;
	wire [8-1:0] node6841;
	wire [8-1:0] node6842;
	wire [8-1:0] node6845;
	wire [8-1:0] node6848;
	wire [8-1:0] node6849;
	wire [8-1:0] node6851;
	wire [8-1:0] node6852;
	wire [8-1:0] node6855;
	wire [8-1:0] node6858;
	wire [8-1:0] node6859;
	wire [8-1:0] node6862;
	wire [8-1:0] node6865;
	wire [8-1:0] node6866;
	wire [8-1:0] node6867;
	wire [8-1:0] node6868;
	wire [8-1:0] node6869;
	wire [8-1:0] node6873;
	wire [8-1:0] node6874;
	wire [8-1:0] node6877;
	wire [8-1:0] node6880;
	wire [8-1:0] node6881;
	wire [8-1:0] node6884;
	wire [8-1:0] node6887;
	wire [8-1:0] node6888;
	wire [8-1:0] node6889;
	wire [8-1:0] node6892;
	wire [8-1:0] node6895;
	wire [8-1:0] node6896;
	wire [8-1:0] node6899;
	wire [8-1:0] node6902;
	wire [8-1:0] node6903;
	wire [8-1:0] node6904;
	wire [8-1:0] node6905;
	wire [8-1:0] node6906;
	wire [8-1:0] node6910;
	wire [8-1:0] node6911;
	wire [8-1:0] node6913;
	wire [8-1:0] node6916;
	wire [8-1:0] node6917;
	wire [8-1:0] node6921;
	wire [8-1:0] node6922;
	wire [8-1:0] node6924;
	wire [8-1:0] node6927;
	wire [8-1:0] node6928;
	wire [8-1:0] node6932;
	wire [8-1:0] node6933;
	wire [8-1:0] node6934;
	wire [8-1:0] node6935;
	wire [8-1:0] node6936;
	wire [8-1:0] node6940;
	wire [8-1:0] node6941;
	wire [8-1:0] node6945;
	wire [8-1:0] node6946;
	wire [8-1:0] node6950;
	wire [8-1:0] node6951;
	wire [8-1:0] node6952;
	wire [8-1:0] node6954;
	wire [8-1:0] node6957;
	wire [8-1:0] node6958;
	wire [8-1:0] node6961;
	wire [8-1:0] node6964;
	wire [8-1:0] node6965;
	wire [8-1:0] node6966;
	wire [8-1:0] node6970;
	wire [8-1:0] node6971;
	wire [8-1:0] node6975;
	wire [8-1:0] node6976;
	wire [8-1:0] node6977;
	wire [8-1:0] node6978;
	wire [8-1:0] node6979;
	wire [8-1:0] node6980;
	wire [8-1:0] node6981;
	wire [8-1:0] node6982;
	wire [8-1:0] node6985;
	wire [8-1:0] node6987;
	wire [8-1:0] node6990;
	wire [8-1:0] node6991;
	wire [8-1:0] node6992;
	wire [8-1:0] node6995;
	wire [8-1:0] node6998;
	wire [8-1:0] node6999;
	wire [8-1:0] node7002;
	wire [8-1:0] node7005;
	wire [8-1:0] node7006;
	wire [8-1:0] node7007;
	wire [8-1:0] node7009;
	wire [8-1:0] node7012;
	wire [8-1:0] node7014;
	wire [8-1:0] node7017;
	wire [8-1:0] node7018;
	wire [8-1:0] node7019;
	wire [8-1:0] node7022;
	wire [8-1:0] node7025;
	wire [8-1:0] node7026;
	wire [8-1:0] node7030;
	wire [8-1:0] node7031;
	wire [8-1:0] node7032;
	wire [8-1:0] node7033;
	wire [8-1:0] node7034;
	wire [8-1:0] node7037;
	wire [8-1:0] node7040;
	wire [8-1:0] node7042;
	wire [8-1:0] node7045;
	wire [8-1:0] node7046;
	wire [8-1:0] node7048;
	wire [8-1:0] node7051;
	wire [8-1:0] node7052;
	wire [8-1:0] node7056;
	wire [8-1:0] node7057;
	wire [8-1:0] node7058;
	wire [8-1:0] node7060;
	wire [8-1:0] node7063;
	wire [8-1:0] node7064;
	wire [8-1:0] node7067;
	wire [8-1:0] node7070;
	wire [8-1:0] node7071;
	wire [8-1:0] node7072;
	wire [8-1:0] node7076;
	wire [8-1:0] node7077;
	wire [8-1:0] node7081;
	wire [8-1:0] node7082;
	wire [8-1:0] node7083;
	wire [8-1:0] node7084;
	wire [8-1:0] node7085;
	wire [8-1:0] node7088;
	wire [8-1:0] node7091;
	wire [8-1:0] node7094;
	wire [8-1:0] node7095;
	wire [8-1:0] node7096;
	wire [8-1:0] node7099;
	wire [8-1:0] node7102;
	wire [8-1:0] node7105;
	wire [8-1:0] node7106;
	wire [8-1:0] node7107;
	wire [8-1:0] node7110;
	wire [8-1:0] node7113;
	wire [8-1:0] node7116;
	wire [8-1:0] node7117;
	wire [8-1:0] node7118;
	wire [8-1:0] node7119;
	wire [8-1:0] node7120;
	wire [8-1:0] node7122;
	wire [8-1:0] node7123;
	wire [8-1:0] node7126;
	wire [8-1:0] node7129;
	wire [8-1:0] node7130;
	wire [8-1:0] node7131;
	wire [8-1:0] node7134;
	wire [8-1:0] node7138;
	wire [8-1:0] node7139;
	wire [8-1:0] node7140;
	wire [8-1:0] node7143;
	wire [8-1:0] node7146;
	wire [8-1:0] node7147;
	wire [8-1:0] node7149;
	wire [8-1:0] node7152;
	wire [8-1:0] node7155;
	wire [8-1:0] node7156;
	wire [8-1:0] node7157;
	wire [8-1:0] node7158;
	wire [8-1:0] node7161;
	wire [8-1:0] node7164;
	wire [8-1:0] node7165;
	wire [8-1:0] node7166;
	wire [8-1:0] node7170;
	wire [8-1:0] node7171;
	wire [8-1:0] node7175;
	wire [8-1:0] node7176;
	wire [8-1:0] node7177;
	wire [8-1:0] node7178;
	wire [8-1:0] node7181;
	wire [8-1:0] node7184;
	wire [8-1:0] node7185;
	wire [8-1:0] node7189;
	wire [8-1:0] node7192;
	wire [8-1:0] node7193;
	wire [8-1:0] node7194;
	wire [8-1:0] node7195;
	wire [8-1:0] node7196;
	wire [8-1:0] node7197;
	wire [8-1:0] node7200;
	wire [8-1:0] node7204;
	wire [8-1:0] node7205;
	wire [8-1:0] node7207;
	wire [8-1:0] node7211;
	wire [8-1:0] node7212;
	wire [8-1:0] node7213;
	wire [8-1:0] node7214;
	wire [8-1:0] node7217;
	wire [8-1:0] node7221;
	wire [8-1:0] node7222;
	wire [8-1:0] node7223;
	wire [8-1:0] node7226;
	wire [8-1:0] node7230;
	wire [8-1:0] node7231;
	wire [8-1:0] node7232;
	wire [8-1:0] node7233;
	wire [8-1:0] node7235;
	wire [8-1:0] node7238;
	wire [8-1:0] node7239;
	wire [8-1:0] node7242;
	wire [8-1:0] node7245;
	wire [8-1:0] node7246;
	wire [8-1:0] node7247;
	wire [8-1:0] node7251;
	wire [8-1:0] node7253;
	wire [8-1:0] node7256;
	wire [8-1:0] node7259;
	wire [8-1:0] node7260;
	wire [8-1:0] node7261;
	wire [8-1:0] node7262;
	wire [8-1:0] node7263;
	wire [8-1:0] node7264;
	wire [8-1:0] node7265;
	wire [8-1:0] node7266;
	wire [8-1:0] node7269;
	wire [8-1:0] node7272;
	wire [8-1:0] node7274;
	wire [8-1:0] node7277;
	wire [8-1:0] node7278;
	wire [8-1:0] node7279;
	wire [8-1:0] node7282;
	wire [8-1:0] node7285;
	wire [8-1:0] node7286;
	wire [8-1:0] node7290;
	wire [8-1:0] node7291;
	wire [8-1:0] node7292;
	wire [8-1:0] node7293;
	wire [8-1:0] node7296;
	wire [8-1:0] node7299;
	wire [8-1:0] node7300;
	wire [8-1:0] node7303;
	wire [8-1:0] node7306;
	wire [8-1:0] node7307;
	wire [8-1:0] node7308;
	wire [8-1:0] node7311;
	wire [8-1:0] node7314;
	wire [8-1:0] node7315;
	wire [8-1:0] node7318;
	wire [8-1:0] node7321;
	wire [8-1:0] node7322;
	wire [8-1:0] node7323;
	wire [8-1:0] node7326;
	wire [8-1:0] node7329;
	wire [8-1:0] node7332;
	wire [8-1:0] node7333;
	wire [8-1:0] node7334;
	wire [8-1:0] node7335;
	wire [8-1:0] node7336;
	wire [8-1:0] node7337;
	wire [8-1:0] node7340;
	wire [8-1:0] node7344;
	wire [8-1:0] node7345;
	wire [8-1:0] node7347;
	wire [8-1:0] node7351;
	wire [8-1:0] node7352;
	wire [8-1:0] node7353;
	wire [8-1:0] node7357;
	wire [8-1:0] node7358;
	wire [8-1:0] node7360;
	wire [8-1:0] node7364;
	wire [8-1:0] node7365;
	wire [8-1:0] node7366;
	wire [8-1:0] node7367;
	wire [8-1:0] node7368;
	wire [8-1:0] node7371;
	wire [8-1:0] node7374;
	wire [8-1:0] node7375;
	wire [8-1:0] node7378;
	wire [8-1:0] node7381;
	wire [8-1:0] node7382;
	wire [8-1:0] node7383;
	wire [8-1:0] node7386;
	wire [8-1:0] node7389;
	wire [8-1:0] node7390;
	wire [8-1:0] node7393;
	wire [8-1:0] node7396;
	wire [8-1:0] node7399;
	wire [8-1:0] node7400;
	wire [8-1:0] node7401;
	wire [8-1:0] node7402;
	wire [8-1:0] node7403;
	wire [8-1:0] node7404;
	wire [8-1:0] node7405;
	wire [8-1:0] node7409;
	wire [8-1:0] node7410;
	wire [8-1:0] node7414;
	wire [8-1:0] node7415;
	wire [8-1:0] node7416;
	wire [8-1:0] node7420;
	wire [8-1:0] node7421;
	wire [8-1:0] node7424;
	wire [8-1:0] node7427;
	wire [8-1:0] node7428;
	wire [8-1:0] node7429;
	wire [8-1:0] node7430;
	wire [8-1:0] node7433;
	wire [8-1:0] node7436;
	wire [8-1:0] node7437;
	wire [8-1:0] node7441;
	wire [8-1:0] node7442;
	wire [8-1:0] node7443;
	wire [8-1:0] node7446;
	wire [8-1:0] node7449;
	wire [8-1:0] node7451;
	wire [8-1:0] node7454;
	wire [8-1:0] node7455;
	wire [8-1:0] node7456;
	wire [8-1:0] node7457;
	wire [8-1:0] node7458;
	wire [8-1:0] node7461;
	wire [8-1:0] node7464;
	wire [8-1:0] node7466;
	wire [8-1:0] node7469;
	wire [8-1:0] node7470;
	wire [8-1:0] node7471;
	wire [8-1:0] node7475;
	wire [8-1:0] node7476;
	wire [8-1:0] node7479;
	wire [8-1:0] node7482;
	wire [8-1:0] node7483;
	wire [8-1:0] node7484;
	wire [8-1:0] node7485;
	wire [8-1:0] node7488;
	wire [8-1:0] node7492;
	wire [8-1:0] node7493;
	wire [8-1:0] node7494;
	wire [8-1:0] node7497;
	wire [8-1:0] node7500;
	wire [8-1:0] node7501;
	wire [8-1:0] node7504;
	wire [8-1:0] node7507;
	wire [8-1:0] node7508;
	wire [8-1:0] node7509;
	wire [8-1:0] node7512;
	wire [8-1:0] node7515;
	wire [8-1:0] node7518;
	wire [8-1:0] node7519;
	wire [8-1:0] node7520;
	wire [8-1:0] node7521;
	wire [8-1:0] node7524;
	wire [8-1:0] node7525;
	wire [8-1:0] node7526;
	wire [8-1:0] node7527;
	wire [8-1:0] node7528;
	wire [8-1:0] node7530;
	wire [8-1:0] node7533;
	wire [8-1:0] node7535;
	wire [8-1:0] node7538;
	wire [8-1:0] node7539;
	wire [8-1:0] node7540;
	wire [8-1:0] node7542;
	wire [8-1:0] node7545;
	wire [8-1:0] node7547;
	wire [8-1:0] node7550;
	wire [8-1:0] node7552;
	wire [8-1:0] node7555;
	wire [8-1:0] node7556;
	wire [8-1:0] node7557;
	wire [8-1:0] node7558;
	wire [8-1:0] node7560;
	wire [8-1:0] node7563;
	wire [8-1:0] node7565;
	wire [8-1:0] node7568;
	wire [8-1:0] node7569;
	wire [8-1:0] node7570;
	wire [8-1:0] node7573;
	wire [8-1:0] node7574;
	wire [8-1:0] node7578;
	wire [8-1:0] node7580;
	wire [8-1:0] node7583;
	wire [8-1:0] node7584;
	wire [8-1:0] node7586;
	wire [8-1:0] node7589;
	wire [8-1:0] node7590;
	wire [8-1:0] node7592;
	wire [8-1:0] node7595;
	wire [8-1:0] node7597;
	wire [8-1:0] node7600;
	wire [8-1:0] node7601;
	wire [8-1:0] node7602;
	wire [8-1:0] node7603;
	wire [8-1:0] node7604;
	wire [8-1:0] node7606;
	wire [8-1:0] node7609;
	wire [8-1:0] node7611;
	wire [8-1:0] node7614;
	wire [8-1:0] node7615;
	wire [8-1:0] node7616;
	wire [8-1:0] node7619;
	wire [8-1:0] node7620;
	wire [8-1:0] node7624;
	wire [8-1:0] node7626;
	wire [8-1:0] node7629;
	wire [8-1:0] node7630;
	wire [8-1:0] node7631;
	wire [8-1:0] node7632;
	wire [8-1:0] node7634;
	wire [8-1:0] node7638;
	wire [8-1:0] node7639;
	wire [8-1:0] node7640;
	wire [8-1:0] node7643;
	wire [8-1:0] node7644;
	wire [8-1:0] node7648;
	wire [8-1:0] node7651;
	wire [8-1:0] node7652;
	wire [8-1:0] node7654;
	wire [8-1:0] node7657;
	wire [8-1:0] node7658;
	wire [8-1:0] node7660;
	wire [8-1:0] node7663;
	wire [8-1:0] node7665;
	wire [8-1:0] node7668;
	wire [8-1:0] node7669;
	wire [8-1:0] node7670;
	wire [8-1:0] node7672;
	wire [8-1:0] node7675;
	wire [8-1:0] node7676;
	wire [8-1:0] node7678;
	wire [8-1:0] node7681;
	wire [8-1:0] node7683;
	wire [8-1:0] node7686;
	wire [8-1:0] node7687;
	wire [8-1:0] node7688;
	wire [8-1:0] node7690;
	wire [8-1:0] node7693;
	wire [8-1:0] node7695;
	wire [8-1:0] node7697;
	wire [8-1:0] node7700;
	wire [8-1:0] node7701;
	wire [8-1:0] node7703;
	wire [8-1:0] node7706;
	wire [8-1:0] node7707;
	wire [8-1:0] node7709;
	wire [8-1:0] node7712;
	wire [8-1:0] node7714;
	wire [8-1:0] node7717;
	wire [8-1:0] node7718;
	wire [8-1:0] node7719;
	wire [8-1:0] node7720;
	wire [8-1:0] node7721;
	wire [8-1:0] node7724;
	wire [8-1:0] node7726;
	wire [8-1:0] node7727;
	wire [8-1:0] node7731;
	wire [8-1:0] node7732;
	wire [8-1:0] node7733;
	wire [8-1:0] node7735;
	wire [8-1:0] node7739;
	wire [8-1:0] node7740;
	wire [8-1:0] node7741;
	wire [8-1:0] node7744;
	wire [8-1:0] node7746;
	wire [8-1:0] node7750;
	wire [8-1:0] node7751;
	wire [8-1:0] node7752;
	wire [8-1:0] node7754;
	wire [8-1:0] node7755;
	wire [8-1:0] node7759;
	wire [8-1:0] node7760;
	wire [8-1:0] node7761;
	wire [8-1:0] node7764;
	wire [8-1:0] node7766;
	wire [8-1:0] node7770;
	wire [8-1:0] node7771;
	wire [8-1:0] node7772;
	wire [8-1:0] node7773;
	wire [8-1:0] node7775;
	wire [8-1:0] node7778;
	wire [8-1:0] node7780;
	wire [8-1:0] node7783;
	wire [8-1:0] node7784;
	wire [8-1:0] node7786;
	wire [8-1:0] node7789;
	wire [8-1:0] node7790;
	wire [8-1:0] node7793;
	wire [8-1:0] node7795;
	wire [8-1:0] node7798;
	wire [8-1:0] node7801;
	wire [8-1:0] node7802;
	wire [8-1:0] node7803;
	wire [8-1:0] node7804;
	wire [8-1:0] node7805;
	wire [8-1:0] node7807;
	wire [8-1:0] node7811;
	wire [8-1:0] node7812;
	wire [8-1:0] node7813;
	wire [8-1:0] node7816;
	wire [8-1:0] node7818;
	wire [8-1:0] node7822;
	wire [8-1:0] node7823;
	wire [8-1:0] node7824;
	wire [8-1:0] node7825;
	wire [8-1:0] node7826;
	wire [8-1:0] node7830;
	wire [8-1:0] node7832;
	wire [8-1:0] node7835;
	wire [8-1:0] node7836;
	wire [8-1:0] node7838;
	wire [8-1:0] node7841;
	wire [8-1:0] node7842;
	wire [8-1:0] node7843;
	wire [8-1:0] node7847;
	wire [8-1:0] node7850;
	wire [8-1:0] node7853;
	wire [8-1:0] node7854;
	wire [8-1:0] node7855;
	wire [8-1:0] node7856;
	wire [8-1:0] node7857;
	wire [8-1:0] node7858;
	wire [8-1:0] node7862;
	wire [8-1:0] node7863;
	wire [8-1:0] node7865;
	wire [8-1:0] node7868;
	wire [8-1:0] node7870;
	wire [8-1:0] node7873;
	wire [8-1:0] node7874;
	wire [8-1:0] node7875;
	wire [8-1:0] node7877;
	wire [8-1:0] node7880;
	wire [8-1:0] node7882;
	wire [8-1:0] node7885;
	wire [8-1:0] node7886;
	wire [8-1:0] node7890;
	wire [8-1:0] node7891;
	wire [8-1:0] node7892;
	wire [8-1:0] node7894;
	wire [8-1:0] node7897;
	wire [8-1:0] node7898;
	wire [8-1:0] node7900;
	wire [8-1:0] node7903;
	wire [8-1:0] node7906;
	wire [8-1:0] node7907;
	wire [8-1:0] node7908;
	wire [8-1:0] node7909;
	wire [8-1:0] node7913;
	wire [8-1:0] node7914;
	wire [8-1:0] node7918;
	wire [8-1:0] node7919;
	wire [8-1:0] node7920;
	wire [8-1:0] node7924;
	wire [8-1:0] node7925;
	wire [8-1:0] node7928;
	wire [8-1:0] node7931;
	wire [8-1:0] node7932;
	wire [8-1:0] node7935;
	wire [8-1:0] node7938;
	wire [8-1:0] node7939;
	wire [8-1:0] node7940;
	wire [8-1:0] node7942;
	wire [8-1:0] node7943;
	wire [8-1:0] node7944;
	wire [8-1:0] node7945;
	wire [8-1:0] node7946;
	wire [8-1:0] node7947;
	wire [8-1:0] node7951;
	wire [8-1:0] node7952;
	wire [8-1:0] node7956;
	wire [8-1:0] node7958;
	wire [8-1:0] node7961;
	wire [8-1:0] node7962;
	wire [8-1:0] node7963;
	wire [8-1:0] node7964;
	wire [8-1:0] node7968;
	wire [8-1:0] node7969;
	wire [8-1:0] node7971;
	wire [8-1:0] node7974;
	wire [8-1:0] node7976;
	wire [8-1:0] node7979;
	wire [8-1:0] node7980;
	wire [8-1:0] node7981;
	wire [8-1:0] node7982;
	wire [8-1:0] node7986;
	wire [8-1:0] node7988;
	wire [8-1:0] node7991;
	wire [8-1:0] node7992;
	wire [8-1:0] node7996;
	wire [8-1:0] node7997;
	wire [8-1:0] node7998;
	wire [8-1:0] node7999;
	wire [8-1:0] node8000;
	wire [8-1:0] node8002;
	wire [8-1:0] node8005;
	wire [8-1:0] node8006;
	wire [8-1:0] node8010;
	wire [8-1:0] node8011;
	wire [8-1:0] node8015;
	wire [8-1:0] node8016;
	wire [8-1:0] node8017;
	wire [8-1:0] node8019;
	wire [8-1:0] node8022;
	wire [8-1:0] node8023;
	wire [8-1:0] node8025;
	wire [8-1:0] node8028;
	wire [8-1:0] node8029;
	wire [8-1:0] node8033;
	wire [8-1:0] node8034;
	wire [8-1:0] node8035;
	wire [8-1:0] node8038;
	wire [8-1:0] node8040;
	wire [8-1:0] node8043;
	wire [8-1:0] node8045;
	wire [8-1:0] node8048;
	wire [8-1:0] node8049;
	wire [8-1:0] node8050;
	wire [8-1:0] node8051;
	wire [8-1:0] node8052;
	wire [8-1:0] node8056;
	wire [8-1:0] node8057;
	wire [8-1:0] node8059;
	wire [8-1:0] node8062;
	wire [8-1:0] node8064;
	wire [8-1:0] node8067;
	wire [8-1:0] node8068;
	wire [8-1:0] node8069;
	wire [8-1:0] node8071;
	wire [8-1:0] node8074;
	wire [8-1:0] node8075;
	wire [8-1:0] node8079;
	wire [8-1:0] node8081;
	wire [8-1:0] node8084;
	wire [8-1:0] node8085;
	wire [8-1:0] node8087;
	wire [8-1:0] node8090;
	wire [8-1:0] node8091;
	wire [8-1:0] node8093;
	wire [8-1:0] node8096;
	wire [8-1:0] node8098;
	wire [8-1:0] node8101;
	wire [8-1:0] node8102;
	wire [8-1:0] node8103;
	wire [8-1:0] node8104;
	wire [8-1:0] node8106;
	wire [8-1:0] node8107;
	wire [8-1:0] node8111;
	wire [8-1:0] node8112;
	wire [8-1:0] node8113;
	wire [8-1:0] node8115;
	wire [8-1:0] node8118;
	wire [8-1:0] node8121;
	wire [8-1:0] node8123;
	wire [8-1:0] node8124;
	wire [8-1:0] node8128;
	wire [8-1:0] node8129;
	wire [8-1:0] node8130;
	wire [8-1:0] node8131;
	wire [8-1:0] node8133;
	wire [8-1:0] node8136;
	wire [8-1:0] node8138;
	wire [8-1:0] node8141;
	wire [8-1:0] node8144;
	wire [8-1:0] node8145;
	wire [8-1:0] node8146;
	wire [8-1:0] node8147;
	wire [8-1:0] node8149;
	wire [8-1:0] node8153;
	wire [8-1:0] node8154;
	wire [8-1:0] node8156;
	wire [8-1:0] node8159;
	wire [8-1:0] node8161;
	wire [8-1:0] node8164;
	wire [8-1:0] node8167;
	wire [8-1:0] node8168;
	wire [8-1:0] node8169;
	wire [8-1:0] node8170;
	wire [8-1:0] node8171;
	wire [8-1:0] node8173;
	wire [8-1:0] node8176;
	wire [8-1:0] node8179;
	wire [8-1:0] node8181;
	wire [8-1:0] node8182;
	wire [8-1:0] node8186;
	wire [8-1:0] node8187;
	wire [8-1:0] node8188;
	wire [8-1:0] node8189;
	wire [8-1:0] node8191;
	wire [8-1:0] node8194;
	wire [8-1:0] node8196;
	wire [8-1:0] node8199;
	wire [8-1:0] node8200;
	wire [8-1:0] node8202;
	wire [8-1:0] node8205;
	wire [8-1:0] node8207;
	wire [8-1:0] node8210;
	wire [8-1:0] node8213;
	wire [8-1:0] node8214;
	wire [8-1:0] node8215;
	wire [8-1:0] node8216;
	wire [8-1:0] node8217;
	wire [8-1:0] node8219;
	wire [8-1:0] node8222;
	wire [8-1:0] node8224;
	wire [8-1:0] node8227;
	wire [8-1:0] node8228;
	wire [8-1:0] node8230;
	wire [8-1:0] node8233;
	wire [8-1:0] node8235;
	wire [8-1:0] node8238;
	wire [8-1:0] node8241;
	wire [8-1:0] node8242;
	wire [8-1:0] node8243;
	wire [8-1:0] node8244;
	wire [8-1:0] node8246;
	wire [8-1:0] node8249;
	wire [8-1:0] node8250;
	wire [8-1:0] node8252;
	wire [8-1:0] node8255;
	wire [8-1:0] node8257;
	wire [8-1:0] node8260;
	wire [8-1:0] node8261;
	wire [8-1:0] node8262;
	wire [8-1:0] node8266;
	wire [8-1:0] node8268;
	wire [8-1:0] node8270;
	wire [8-1:0] node8273;
	wire [8-1:0] node8276;
	wire [8-1:0] node8277;
	wire [8-1:0] node8279;
	wire [8-1:0] node8280;
	wire [8-1:0] node8281;
	wire [8-1:0] node8282;
	wire [8-1:0] node8284;
	wire [8-1:0] node8287;
	wire [8-1:0] node8288;
	wire [8-1:0] node8290;
	wire [8-1:0] node8293;
	wire [8-1:0] node8295;
	wire [8-1:0] node8298;
	wire [8-1:0] node8299;
	wire [8-1:0] node8300;
	wire [8-1:0] node8302;
	wire [8-1:0] node8305;
	wire [8-1:0] node8306;
	wire [8-1:0] node8308;
	wire [8-1:0] node8311;
	wire [8-1:0] node8313;
	wire [8-1:0] node8316;
	wire [8-1:0] node8317;
	wire [8-1:0] node8319;
	wire [8-1:0] node8322;
	wire [8-1:0] node8323;
	wire [8-1:0] node8325;
	wire [8-1:0] node8328;
	wire [8-1:0] node8330;
	wire [8-1:0] node8333;
	wire [8-1:0] node8334;
	wire [8-1:0] node8335;
	wire [8-1:0] node8336;
	wire [8-1:0] node8338;
	wire [8-1:0] node8341;
	wire [8-1:0] node8342;
	wire [8-1:0] node8344;
	wire [8-1:0] node8347;
	wire [8-1:0] node8349;
	wire [8-1:0] node8352;
	wire [8-1:0] node8353;
	wire [8-1:0] node8354;
	wire [8-1:0] node8356;
	wire [8-1:0] node8359;
	wire [8-1:0] node8360;
	wire [8-1:0] node8363;
	wire [8-1:0] node8365;
	wire [8-1:0] node8368;
	wire [8-1:0] node8369;
	wire [8-1:0] node8371;
	wire [8-1:0] node8374;
	wire [8-1:0] node8375;
	wire [8-1:0] node8377;
	wire [8-1:0] node8380;
	wire [8-1:0] node8382;
	wire [8-1:0] node8385;
	wire [8-1:0] node8386;
	wire [8-1:0] node8387;
	wire [8-1:0] node8389;
	wire [8-1:0] node8392;
	wire [8-1:0] node8393;
	wire [8-1:0] node8395;
	wire [8-1:0] node8398;
	wire [8-1:0] node8400;
	wire [8-1:0] node8403;
	wire [8-1:0] node8404;
	wire [8-1:0] node8405;
	wire [8-1:0] node8407;
	wire [8-1:0] node8410;
	wire [8-1:0] node8411;
	wire [8-1:0] node8413;
	wire [8-1:0] node8416;
	wire [8-1:0] node8418;
	wire [8-1:0] node8421;
	wire [8-1:0] node8422;
	wire [8-1:0] node8424;
	wire [8-1:0] node8427;
	wire [8-1:0] node8429;
	wire [8-1:0] node8431;
	wire [8-1:0] node8434;
	wire [8-1:0] node8435;
	wire [8-1:0] node8436;
	wire [8-1:0] node8437;
	wire [8-1:0] node8439;
	wire [8-1:0] node8441;
	wire [8-1:0] node8444;
	wire [8-1:0] node8445;
	wire [8-1:0] node8447;
	wire [8-1:0] node8449;
	wire [8-1:0] node8452;
	wire [8-1:0] node8453;
	wire [8-1:0] node8455;
	wire [8-1:0] node8458;
	wire [8-1:0] node8461;
	wire [8-1:0] node8462;
	wire [8-1:0] node8463;
	wire [8-1:0] node8465;
	wire [8-1:0] node8466;
	wire [8-1:0] node8470;
	wire [8-1:0] node8471;
	wire [8-1:0] node8473;
	wire [8-1:0] node8476;
	wire [8-1:0] node8477;
	wire [8-1:0] node8478;
	wire [8-1:0] node8481;
	wire [8-1:0] node8485;
	wire [8-1:0] node8486;
	wire [8-1:0] node8487;
	wire [8-1:0] node8488;
	wire [8-1:0] node8492;
	wire [8-1:0] node8493;
	wire [8-1:0] node8494;
	wire [8-1:0] node8498;
	wire [8-1:0] node8500;
	wire [8-1:0] node8503;
	wire [8-1:0] node8504;
	wire [8-1:0] node8507;
	wire [8-1:0] node8510;
	wire [8-1:0] node8511;
	wire [8-1:0] node8512;
	wire [8-1:0] node8513;
	wire [8-1:0] node8515;
	wire [8-1:0] node8517;
	wire [8-1:0] node8520;
	wire [8-1:0] node8521;
	wire [8-1:0] node8523;
	wire [8-1:0] node8524;
	wire [8-1:0] node8528;
	wire [8-1:0] node8531;
	wire [8-1:0] node8532;
	wire [8-1:0] node8533;
	wire [8-1:0] node8535;
	wire [8-1:0] node8538;
	wire [8-1:0] node8539;
	wire [8-1:0] node8540;
	wire [8-1:0] node8543;
	wire [8-1:0] node8547;
	wire [8-1:0] node8548;
	wire [8-1:0] node8549;
	wire [8-1:0] node8550;
	wire [8-1:0] node8552;
	wire [8-1:0] node8555;
	wire [8-1:0] node8557;
	wire [8-1:0] node8560;
	wire [8-1:0] node8561;
	wire [8-1:0] node8562;
	wire [8-1:0] node8566;
	wire [8-1:0] node8568;
	wire [8-1:0] node8571;
	wire [8-1:0] node8574;
	wire [8-1:0] node8575;
	wire [8-1:0] node8576;
	wire [8-1:0] node8577;
	wire [8-1:0] node8578;
	wire [8-1:0] node8582;
	wire [8-1:0] node8583;
	wire [8-1:0] node8584;
	wire [8-1:0] node8588;
	wire [8-1:0] node8590;
	wire [8-1:0] node8593;
	wire [8-1:0] node8594;
	wire [8-1:0] node8595;
	wire [8-1:0] node8597;
	wire [8-1:0] node8600;
	wire [8-1:0] node8601;
	wire [8-1:0] node8603;
	wire [8-1:0] node8607;
	wire [8-1:0] node8608;
	wire [8-1:0] node8609;
	wire [8-1:0] node8610;
	wire [8-1:0] node8614;
	wire [8-1:0] node8617;
	wire [8-1:0] node8618;
	wire [8-1:0] node8622;
	wire [8-1:0] node8623;
	wire [8-1:0] node8624;
	wire [8-1:0] node8627;
	wire [8-1:0] node8630;
	wire [8-1:0] node8631;
	wire [8-1:0] node8634;

	assign outp = (inp[7]) ? node4322 : node1;
		assign node1 = (inp[13]) ? node2091 : node2;
			assign node2 = (inp[4]) ? node398 : node3;
				assign node3 = (inp[11]) ? node127 : node4;
					assign node4 = (inp[0]) ? node72 : node5;
						assign node5 = (inp[8]) ? node29 : node6;
							assign node6 = (inp[2]) ? node14 : node7;
								assign node7 = (inp[1]) ? node9 : 8'b01111111;
									assign node9 = (inp[5]) ? node11 : 8'b00111110;
										assign node11 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node14 = (inp[1]) ? node20 : node15;
									assign node15 = (inp[6]) ? node17 : 8'b00101111;
										assign node17 = (inp[5]) ? 8'b01111111 : 8'b00101111;
									assign node20 = (inp[5]) ? node22 : 8'b00101110;
										assign node22 = (inp[6]) ? node26 : node23;
											assign node23 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node26 = (inp[3]) ? 8'b01111111 : 8'b00111110;
							assign node29 = (inp[1]) ? node45 : node30;
								assign node30 = (inp[2]) ? node36 : node31;
									assign node31 = (inp[5]) ? node33 : 8'b00111011;
										assign node33 = (inp[10]) ? 8'b01111111 : 8'b00111011;
									assign node36 = (inp[5]) ? node38 : 8'b00101011;
										assign node38 = (inp[10]) ? node42 : node39;
											assign node39 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node42 = (inp[6]) ? 8'b01111111 : 8'b00101111;
								assign node45 = (inp[5]) ? node49 : node46;
									assign node46 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node49 = (inp[10]) ? node61 : node50;
										assign node50 = (inp[3]) ? node56 : node51;
											assign node51 = (inp[6]) ? 8'b00111010 : node52;
												assign node52 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node56 = (inp[2]) ? node58 : 8'b00111011;
												assign node58 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node61 = (inp[3]) ? node67 : node62;
											assign node62 = (inp[6]) ? 8'b00111110 : node63;
												assign node63 = (inp[2]) ? 8'b00101110 : 8'b00111110;
											assign node67 = (inp[6]) ? 8'b01111111 : node68;
												assign node68 = (inp[2]) ? 8'b00101111 : 8'b01111111;
						assign node72 = (inp[5]) ? 8'b01111111 : node73;
							assign node73 = (inp[2]) ? node91 : node74;
								assign node74 = (inp[3]) ? node80 : node75;
									assign node75 = (inp[8]) ? node77 : 8'b01111111;
										assign node77 = (inp[10]) ? 8'b00111011 : 8'b01111111;
									assign node80 = (inp[1]) ? node86 : node81;
										assign node81 = (inp[10]) ? node83 : 8'b01111111;
											assign node83 = (inp[8]) ? 8'b00111011 : 8'b01111111;
										assign node86 = (inp[10]) ? node88 : 8'b00111110;
											assign node88 = (inp[8]) ? 8'b00111010 : 8'b00111110;
								assign node91 = (inp[6]) ? node109 : node92;
									assign node92 = (inp[3]) ? node98 : node93;
										assign node93 = (inp[8]) ? node95 : 8'b01111111;
											assign node95 = (inp[10]) ? 8'b00111011 : 8'b01111111;
										assign node98 = (inp[1]) ? node104 : node99;
											assign node99 = (inp[8]) ? node101 : 8'b01111111;
												assign node101 = (inp[10]) ? 8'b00111011 : 8'b01111111;
											assign node104 = (inp[10]) ? node106 : 8'b00111110;
												assign node106 = (inp[8]) ? 8'b00111010 : 8'b00111110;
									assign node109 = (inp[10]) ? node115 : node110;
										assign node110 = (inp[3]) ? node112 : 8'b00101111;
											assign node112 = (inp[1]) ? 8'b00101110 : 8'b00101111;
										assign node115 = (inp[8]) ? node121 : node116;
											assign node116 = (inp[1]) ? node118 : 8'b00101111;
												assign node118 = (inp[3]) ? 8'b00101110 : 8'b00101111;
											assign node121 = (inp[3]) ? node123 : 8'b00101011;
												assign node123 = (inp[1]) ? 8'b00101010 : 8'b00101011;
					assign node127 = (inp[8]) ? node219 : node128;
						assign node128 = (inp[1]) ? node156 : node129;
							assign node129 = (inp[2]) ? node133 : node130;
								assign node130 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node133 = (inp[12]) ? node145 : node134;
									assign node134 = (inp[0]) ? node140 : node135;
										assign node135 = (inp[6]) ? node137 : 8'b00111110;
											assign node137 = (inp[5]) ? 8'b00101110 : 8'b00111110;
										assign node140 = (inp[5]) ? 8'b00101110 : node141;
											assign node141 = (inp[6]) ? 8'b00111110 : 8'b00101110;
									assign node145 = (inp[0]) ? node151 : node146;
										assign node146 = (inp[5]) ? node148 : 8'b00101111;
											assign node148 = (inp[6]) ? 8'b00111110 : 8'b00101111;
										assign node151 = (inp[5]) ? 8'b00111110 : node152;
											assign node152 = (inp[6]) ? 8'b00101111 : 8'b00111110;
							assign node156 = (inp[12]) ? node188 : node157;
								assign node157 = (inp[2]) ? node169 : node158;
									assign node158 = (inp[0]) ? node164 : node159;
										assign node159 = (inp[3]) ? node161 : 8'b00101110;
											assign node161 = (inp[5]) ? 8'b00101011 : 8'b00101110;
										assign node164 = (inp[3]) ? node166 : 8'b00101011;
											assign node166 = (inp[5]) ? 8'b00101011 : 8'b00101110;
									assign node169 = (inp[5]) ? node179 : node170;
										assign node170 = (inp[0]) ? node172 : 8'b00111011;
											assign node172 = (inp[3]) ? node176 : node173;
												assign node173 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node176 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node179 = (inp[0]) ? 8'b00101010 : node180;
											assign node180 = (inp[3]) ? node184 : node181;
												assign node181 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node184 = (inp[6]) ? 8'b00101010 : 8'b00111010;
								assign node188 = (inp[5]) ? node204 : node189;
									assign node189 = (inp[2]) ? node195 : node190;
										assign node190 = (inp[3]) ? 8'b00111110 : node191;
											assign node191 = (inp[0]) ? 8'b00111011 : 8'b00111110;
										assign node195 = (inp[0]) ? node197 : 8'b00101110;
											assign node197 = (inp[6]) ? node201 : node198;
												assign node198 = (inp[9]) ? 8'b00111010 : 8'b00111011;
												assign node201 = (inp[3]) ? 8'b00101110 : 8'b00101011;
									assign node204 = (inp[2]) ? node210 : node205;
										assign node205 = (inp[3]) ? 8'b00111011 : node206;
											assign node206 = (inp[0]) ? 8'b00111011 : 8'b00111110;
										assign node210 = (inp[0]) ? 8'b00111010 : node211;
											assign node211 = (inp[6]) ? node215 : node212;
												assign node212 = (inp[3]) ? 8'b00101011 : 8'b00101110;
												assign node215 = (inp[3]) ? 8'b00111010 : 8'b00111011;
						assign node219 = (inp[12]) ? node307 : node220;
							assign node220 = (inp[2]) ? node252 : node221;
								assign node221 = (inp[0]) ? node237 : node222;
									assign node222 = (inp[1]) ? node228 : node223;
										assign node223 = (inp[5]) ? node225 : 8'b00101011;
											assign node225 = (inp[10]) ? 8'b00001111 : 8'b00101011;
										assign node228 = (inp[5]) ? node230 : 8'b00101010;
											assign node230 = (inp[3]) ? node234 : node231;
												assign node231 = (inp[10]) ? 8'b00001110 : 8'b00101010;
												assign node234 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node237 = (inp[1]) ? node243 : node238;
										assign node238 = (inp[5]) ? 8'b00001111 : node239;
											assign node239 = (inp[10]) ? 8'b00101011 : 8'b00001111;
										assign node243 = (inp[5]) ? 8'b00001011 : node244;
											assign node244 = (inp[3]) ? node248 : node245;
												assign node245 = (inp[10]) ? 8'b00001111 : 8'b00001011;
												assign node248 = (inp[10]) ? 8'b00101010 : 8'b00001110;
								assign node252 = (inp[1]) ? node272 : node253;
									assign node253 = (inp[0]) ? node263 : node254;
										assign node254 = (inp[5]) ? node256 : 8'b00111010;
											assign node256 = (inp[10]) ? node260 : node257;
												assign node257 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node260 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node263 = (inp[5]) ? 8'b00001110 : node264;
											assign node264 = (inp[10]) ? node268 : node265;
												assign node265 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node268 = (inp[6]) ? 8'b00111010 : 8'b00101010;
									assign node272 = (inp[5]) ? node290 : node273;
										assign node273 = (inp[0]) ? node275 : 8'b00011111;
											assign node275 = (inp[3]) ? node283 : node276;
												assign node276 = (inp[10]) ? node280 : node277;
													assign node277 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node280 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node283 = (inp[10]) ? node287 : node284;
													assign node284 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node287 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node290 = (inp[0]) ? 8'b00001010 : node291;
											assign node291 = (inp[6]) ? node299 : node292;
												assign node292 = (inp[10]) ? node296 : node293;
													assign node293 = (inp[3]) ? 8'b00011110 : 8'b00011111;
													assign node296 = (inp[3]) ? 8'b00011010 : 8'b00011011;
												assign node299 = (inp[10]) ? node303 : node300;
													assign node300 = (inp[3]) ? 8'b00001110 : 8'b00001111;
													assign node303 = (inp[3]) ? 8'b00001010 : 8'b00001011;
							assign node307 = (inp[2]) ? node341 : node308;
								assign node308 = (inp[0]) ? node326 : node309;
									assign node309 = (inp[5]) ? node313 : node310;
										assign node310 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node313 = (inp[10]) ? node319 : node314;
											assign node314 = (inp[1]) ? node316 : 8'b00111011;
												assign node316 = (inp[3]) ? 8'b00011111 : 8'b00111010;
											assign node319 = (inp[3]) ? node323 : node320;
												assign node320 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node323 = (inp[1]) ? 8'b00011011 : 8'b00011111;
									assign node326 = (inp[1]) ? node332 : node327;
										assign node327 = (inp[5]) ? 8'b00011111 : node328;
											assign node328 = (inp[10]) ? 8'b00111011 : 8'b00011111;
										assign node332 = (inp[5]) ? 8'b00011011 : node333;
											assign node333 = (inp[3]) ? node337 : node334;
												assign node334 = (inp[10]) ? 8'b00011111 : 8'b00011011;
												assign node337 = (inp[10]) ? 8'b00111010 : 8'b00011110;
								assign node341 = (inp[5]) ? node369 : node342;
									assign node342 = (inp[0]) ? node346 : node343;
										assign node343 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node346 = (inp[6]) ? node358 : node347;
											assign node347 = (inp[1]) ? node351 : node348;
												assign node348 = (inp[10]) ? 8'b00111010 : 8'b00011110;
												assign node351 = (inp[10]) ? node355 : node352;
													assign node352 = (inp[3]) ? 8'b00011011 : 8'b00011010;
													assign node355 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node358 = (inp[10]) ? node364 : node359;
												assign node359 = (inp[1]) ? node361 : 8'b00001111;
													assign node361 = (inp[3]) ? 8'b00001110 : 8'b00001011;
												assign node364 = (inp[1]) ? node366 : 8'b00101011;
													assign node366 = (inp[3]) ? 8'b00101010 : 8'b00001111;
									assign node369 = (inp[0]) ? node395 : node370;
										assign node370 = (inp[6]) ? node384 : node371;
											assign node371 = (inp[10]) ? node377 : node372;
												assign node372 = (inp[3]) ? node374 : 8'b00101010;
													assign node374 = (inp[1]) ? 8'b00001111 : 8'b00101011;
												assign node377 = (inp[3]) ? node381 : node378;
													assign node378 = (inp[1]) ? 8'b00001110 : 8'b00001111;
													assign node381 = (inp[1]) ? 8'b00001011 : 8'b00001111;
											assign node384 = (inp[1]) ? node388 : node385;
												assign node385 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node388 = (inp[10]) ? node392 : node389;
													assign node389 = (inp[3]) ? 8'b00011110 : 8'b00011111;
													assign node392 = (inp[3]) ? 8'b00011010 : 8'b00011011;
										assign node395 = (inp[1]) ? 8'b00011010 : 8'b00011110;
				assign node398 = (inp[9]) ? node1266 : node399;
					assign node399 = (inp[8]) ? node811 : node400;
						assign node400 = (inp[10]) ? node600 : node401;
							assign node401 = (inp[1]) ? node483 : node402;
								assign node402 = (inp[3]) ? node446 : node403;
									assign node403 = (inp[2]) ? node415 : node404;
										assign node404 = (inp[6]) ? node410 : node405;
											assign node405 = (inp[12]) ? 8'b00000010 : node406;
												assign node406 = (inp[11]) ? 8'b11110111 : 8'b10000010;
											assign node410 = (inp[12]) ? 8'b00011010 : node411;
												assign node411 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node415 = (inp[11]) ? node431 : node416;
											assign node416 = (inp[0]) ? node426 : node417;
												assign node417 = (inp[6]) ? node421 : node418;
													assign node418 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node421 = (inp[5]) ? 8'b10010000 : node422;
														assign node422 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node426 = (inp[5]) ? 8'b10010000 : node427;
													assign node427 = (inp[6]) ? 8'b10000010 : 8'b10010000;
											assign node431 = (inp[12]) ? node441 : node432;
												assign node432 = (inp[0]) ? node436 : node433;
													assign node433 = (inp[6]) ? 8'b10100101 : 8'b11110111;
													assign node436 = (inp[6]) ? node438 : 8'b10100101;
														assign node438 = (inp[5]) ? 8'b10100101 : 8'b11110111;
												assign node441 = (inp[5]) ? node443 : 8'b00000010;
													assign node443 = (inp[6]) ? 8'b11110101 : 8'b00000010;
									assign node446 = (inp[11]) ? node458 : node447;
										assign node447 = (inp[6]) ? node453 : node448;
											assign node448 = (inp[0]) ? node450 : 8'b00001011;
												assign node450 = (inp[2]) ? 8'b00011011 : 8'b00001011;
											assign node453 = (inp[5]) ? 8'b00011011 : node454;
												assign node454 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node458 = (inp[2]) ? node466 : node459;
											assign node459 = (inp[6]) ? node463 : node460;
												assign node460 = (inp[12]) ? 8'b00001011 : 8'b00011010;
												assign node463 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node466 = (inp[5]) ? node476 : node467;
												assign node467 = (inp[12]) ? node471 : node468;
													assign node468 = (inp[0]) ? 8'b00001010 : 8'b00011010;
													assign node471 = (inp[6]) ? 8'b00001011 : node472;
														assign node472 = (inp[0]) ? 8'b00011010 : 8'b00001011;
												assign node476 = (inp[12]) ? 8'b00011010 : node477;
													assign node477 = (inp[6]) ? 8'b00001010 : node478;
														assign node478 = (inp[0]) ? 8'b00001010 : 8'b00011010;
								assign node483 = (inp[11]) ? node529 : node484;
									assign node484 = (inp[5]) ? node508 : node485;
										assign node485 = (inp[6]) ? node499 : node486;
											assign node486 = (inp[0]) ? node490 : node487;
												assign node487 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node490 = (inp[3]) ? node494 : node491;
													assign node491 = (inp[2]) ? 8'b10010001 : 8'b10000001;
													assign node494 = (inp[2]) ? 8'b10010000 : node495;
														assign node495 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node499 = (inp[2]) ? node505 : node500;
												assign node500 = (inp[0]) ? node502 : 8'b00011010;
													assign node502 = (inp[3]) ? 8'b00011010 : 8'b10011001;
												assign node505 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node508 = (inp[6]) ? node518 : node509;
											assign node509 = (inp[0]) ? node515 : node510;
												assign node510 = (inp[3]) ? 8'b10000001 : node511;
													assign node511 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node515 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node518 = (inp[2]) ? node524 : node519;
												assign node519 = (inp[3]) ? 8'b10011001 : node520;
													assign node520 = (inp[0]) ? 8'b10011001 : 8'b00011010;
												assign node524 = (inp[3]) ? 8'b10010001 : node525;
													assign node525 = (inp[0]) ? 8'b10010001 : 8'b10010000;
									assign node529 = (inp[0]) ? node559 : node530;
										assign node530 = (inp[12]) ? node544 : node531;
											assign node531 = (inp[6]) ? node537 : node532;
												assign node532 = (inp[5]) ? node534 : 8'b11110111;
													assign node534 = (inp[3]) ? 8'b10110100 : 8'b11110111;
												assign node537 = (inp[2]) ? node539 : 8'b00001010;
													assign node539 = (inp[5]) ? node541 : 8'b11110111;
														assign node541 = (inp[3]) ? 8'b10100100 : 8'b10100101;
											assign node544 = (inp[5]) ? node550 : node545;
												assign node545 = (inp[2]) ? 8'b00000010 : node546;
													assign node546 = (inp[6]) ? 8'b00011010 : 8'b00000010;
												assign node550 = (inp[3]) ? node554 : node551;
													assign node551 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node554 = (inp[6]) ? node556 : 8'b10100101;
														assign node556 = (inp[2]) ? 8'b10110100 : 8'b11111101;
										assign node559 = (inp[2]) ? node581 : node560;
											assign node560 = (inp[6]) ? node570 : node561;
												assign node561 = (inp[12]) ? node565 : node562;
													assign node562 = (inp[5]) ? 8'b10110100 : 8'b11110111;
													assign node565 = (inp[3]) ? node567 : 8'b10100101;
														assign node567 = (inp[5]) ? 8'b10100101 : 8'b00000010;
												assign node570 = (inp[12]) ? node576 : node571;
													assign node571 = (inp[3]) ? node573 : 8'b10101101;
														assign node573 = (inp[5]) ? 8'b10101101 : 8'b00001010;
													assign node576 = (inp[3]) ? node578 : 8'b11111101;
														assign node578 = (inp[5]) ? 8'b11111101 : 8'b00011010;
											assign node581 = (inp[5]) ? node597 : node582;
												assign node582 = (inp[3]) ? node590 : node583;
													assign node583 = (inp[6]) ? node587 : node584;
														assign node584 = (inp[12]) ? 8'b10110100 : 8'b10100100;
														assign node587 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node590 = (inp[6]) ? node594 : node591;
														assign node591 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node594 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node597 = (inp[12]) ? 8'b10110100 : 8'b10100100;
							assign node600 = (inp[11]) ? node676 : node601;
								assign node601 = (inp[3]) ? node649 : node602;
									assign node602 = (inp[0]) ? node610 : node603;
										assign node603 = (inp[6]) ? node605 : 8'b00001110;
											assign node605 = (inp[5]) ? 8'b00011110 : node606;
												assign node606 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node610 = (inp[1]) ? node628 : node611;
											assign node611 = (inp[5]) ? node623 : node612;
												assign node612 = (inp[12]) ? node618 : node613;
													assign node613 = (inp[2]) ? 8'b00001110 : node614;
														assign node614 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node618 = (inp[2]) ? node620 : 8'b00011110;
														assign node620 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node623 = (inp[6]) ? 8'b00011110 : node624;
													assign node624 = (inp[2]) ? 8'b00011110 : 8'b00001110;
											assign node628 = (inp[5]) ? node644 : node629;
												assign node629 = (inp[12]) ? node637 : node630;
													assign node630 = (inp[6]) ? node634 : node631;
														assign node631 = (inp[2]) ? 8'b00011111 : 8'b00001111;
														assign node634 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node637 = (inp[6]) ? node641 : node638;
														assign node638 = (inp[2]) ? 8'b00011111 : 8'b00001111;
														assign node641 = (inp[2]) ? 8'b00001111 : 8'b00011111;
												assign node644 = (inp[2]) ? 8'b00011111 : node645;
													assign node645 = (inp[6]) ? 8'b00011111 : 8'b00001111;
									assign node649 = (inp[5]) ? node669 : node650;
										assign node650 = (inp[1]) ? node660 : node651;
											assign node651 = (inp[2]) ? node655 : node652;
												assign node652 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node655 = (inp[0]) ? node657 : 8'b00001111;
													assign node657 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node660 = (inp[0]) ? node662 : 8'b00001110;
												assign node662 = (inp[6]) ? node666 : node663;
													assign node663 = (inp[2]) ? 8'b00011110 : 8'b00001110;
													assign node666 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node669 = (inp[6]) ? 8'b00011111 : node670;
											assign node670 = (inp[0]) ? node672 : 8'b00001111;
												assign node672 = (inp[2]) ? 8'b00011111 : 8'b00001111;
								assign node676 = (inp[1]) ? node730 : node677;
									assign node677 = (inp[3]) ? node709 : node678;
										assign node678 = (inp[2]) ? node686 : node679;
											assign node679 = (inp[12]) ? node683 : node680;
												assign node680 = (inp[6]) ? 8'b00001110 : 8'b00011011;
												assign node683 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node686 = (inp[12]) ? node698 : node687;
												assign node687 = (inp[0]) ? node693 : node688;
													assign node688 = (inp[6]) ? node690 : 8'b00011011;
														assign node690 = (inp[5]) ? 8'b00001011 : 8'b00011011;
													assign node693 = (inp[5]) ? 8'b00001011 : node694;
														assign node694 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node698 = (inp[5]) ? node704 : node699;
													assign node699 = (inp[0]) ? node701 : 8'b00001110;
														assign node701 = (inp[6]) ? 8'b00001110 : 8'b00011011;
													assign node704 = (inp[6]) ? 8'b00011011 : node705;
														assign node705 = (inp[0]) ? 8'b00011011 : 8'b00001110;
										assign node709 = (inp[12]) ? node721 : node710;
											assign node710 = (inp[6]) ? node716 : node711;
												assign node711 = (inp[2]) ? node713 : 8'b00011110;
													assign node713 = (inp[0]) ? 8'b00001110 : 8'b00011110;
												assign node716 = (inp[2]) ? node718 : 8'b00001111;
													assign node718 = (inp[5]) ? 8'b00001110 : 8'b00011110;
											assign node721 = (inp[6]) ? node727 : node722;
												assign node722 = (inp[2]) ? node724 : 8'b00001111;
													assign node724 = (inp[0]) ? 8'b00011110 : 8'b00001111;
												assign node727 = (inp[2]) ? 8'b00001111 : 8'b00011111;
									assign node730 = (inp[5]) ? node772 : node731;
										assign node731 = (inp[12]) ? node751 : node732;
											assign node732 = (inp[6]) ? node742 : node733;
												assign node733 = (inp[0]) ? node735 : 8'b00011011;
													assign node735 = (inp[3]) ? node739 : node736;
														assign node736 = (inp[2]) ? 8'b00001010 : 8'b00011010;
														assign node739 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node742 = (inp[2]) ? node748 : node743;
													assign node743 = (inp[0]) ? node745 : 8'b00001110;
														assign node745 = (inp[3]) ? 8'b00001110 : 8'b00001011;
													assign node748 = (inp[0]) ? 8'b00011010 : 8'b00011011;
											assign node751 = (inp[0]) ? node757 : node752;
												assign node752 = (inp[6]) ? node754 : 8'b00001110;
													assign node754 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node757 = (inp[3]) ? node765 : node758;
													assign node758 = (inp[2]) ? node762 : node759;
														assign node759 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node762 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node765 = (inp[6]) ? node769 : node766;
														assign node766 = (inp[2]) ? 8'b00011011 : 8'b00001110;
														assign node769 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node772 = (inp[2]) ? node794 : node773;
											assign node773 = (inp[3]) ? node787 : node774;
												assign node774 = (inp[0]) ? node780 : node775;
													assign node775 = (inp[6]) ? node777 : 8'b00011011;
														assign node777 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node780 = (inp[12]) ? node784 : node781;
														assign node781 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node784 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node787 = (inp[6]) ? node791 : node788;
													assign node788 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node791 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node794 = (inp[0]) ? node808 : node795;
												assign node795 = (inp[3]) ? node801 : node796;
													assign node796 = (inp[12]) ? 8'b00011011 : node797;
														assign node797 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node801 = (inp[6]) ? node805 : node802;
														assign node802 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node805 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node808 = (inp[12]) ? 8'b00011010 : 8'b00001010;
						assign node811 = (inp[0]) ? node1011 : node812;
							assign node812 = (inp[5]) ? node866 : node813;
								assign node813 = (inp[12]) ? node849 : node814;
									assign node814 = (inp[11]) ? node832 : node815;
										assign node815 = (inp[1]) ? node827 : node816;
											assign node816 = (inp[3]) ? node822 : node817;
												assign node817 = (inp[6]) ? node819 : 8'b10000010;
													assign node819 = (inp[2]) ? 8'b10000010 : 8'b00011010;
												assign node822 = (inp[6]) ? node824 : 8'b00001011;
													assign node824 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node827 = (inp[2]) ? 8'b10000010 : node828;
												assign node828 = (inp[6]) ? 8'b00011010 : 8'b10000010;
										assign node832 = (inp[6]) ? node838 : node833;
											assign node833 = (inp[1]) ? 8'b11110111 : node834;
												assign node834 = (inp[3]) ? 8'b00011010 : 8'b11110111;
											assign node838 = (inp[2]) ? node844 : node839;
												assign node839 = (inp[3]) ? node841 : 8'b00001010;
													assign node841 = (inp[1]) ? 8'b00001010 : 8'b00001011;
												assign node844 = (inp[1]) ? 8'b11110111 : node845;
													assign node845 = (inp[3]) ? 8'b00011010 : 8'b11110111;
									assign node849 = (inp[2]) ? node861 : node850;
										assign node850 = (inp[6]) ? node856 : node851;
											assign node851 = (inp[3]) ? node853 : 8'b00000010;
												assign node853 = (inp[1]) ? 8'b00000010 : 8'b00001011;
											assign node856 = (inp[1]) ? 8'b00011010 : node857;
												assign node857 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node861 = (inp[3]) ? node863 : 8'b00000010;
											assign node863 = (inp[1]) ? 8'b00000010 : 8'b00001011;
								assign node866 = (inp[10]) ? node942 : node867;
									assign node867 = (inp[1]) ? node899 : node868;
										assign node868 = (inp[3]) ? node884 : node869;
											assign node869 = (inp[6]) ? node875 : node870;
												assign node870 = (inp[12]) ? 8'b00000010 : node871;
													assign node871 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node875 = (inp[2]) ? node881 : node876;
													assign node876 = (inp[11]) ? node878 : 8'b00011010;
														assign node878 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node881 = (inp[11]) ? 8'b11110101 : 8'b10010000;
											assign node884 = (inp[6]) ? node890 : node885;
												assign node885 = (inp[12]) ? 8'b00001011 : node886;
													assign node886 = (inp[11]) ? 8'b00011010 : 8'b00001011;
												assign node890 = (inp[11]) ? node892 : 8'b00011011;
													assign node892 = (inp[2]) ? node896 : node893;
														assign node893 = (inp[12]) ? 8'b00011011 : 8'b00001011;
														assign node896 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node899 = (inp[3]) ? node925 : node900;
											assign node900 = (inp[2]) ? node912 : node901;
												assign node901 = (inp[6]) ? node907 : node902;
													assign node902 = (inp[12]) ? 8'b00000010 : node903;
														assign node903 = (inp[11]) ? 8'b11110111 : 8'b10000010;
													assign node907 = (inp[11]) ? node909 : 8'b00011010;
														assign node909 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node912 = (inp[11]) ? node918 : node913;
													assign node913 = (inp[6]) ? 8'b10010000 : node914;
														assign node914 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node918 = (inp[6]) ? node922 : node919;
														assign node919 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node922 = (inp[12]) ? 8'b11110101 : 8'b10100101;
											assign node925 = (inp[11]) ? node931 : node926;
												assign node926 = (inp[6]) ? node928 : 8'b10000001;
													assign node928 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node931 = (inp[2]) ? node937 : node932;
													assign node932 = (inp[6]) ? 8'b10101101 : node933;
														assign node933 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node937 = (inp[12]) ? node939 : 8'b10110100;
														assign node939 = (inp[6]) ? 8'b10110100 : 8'b10100101;
									assign node942 = (inp[11]) ? node958 : node943;
										assign node943 = (inp[3]) ? node949 : node944;
											assign node944 = (inp[6]) ? node946 : 8'b10000100;
												assign node946 = (inp[2]) ? 8'b10010100 : 8'b10011100;
											assign node949 = (inp[6]) ? node953 : node950;
												assign node950 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node953 = (inp[2]) ? node955 : 8'b10011101;
													assign node955 = (inp[1]) ? 8'b10010101 : 8'b10011101;
										assign node958 = (inp[1]) ? node982 : node959;
											assign node959 = (inp[3]) ? node969 : node960;
												assign node960 = (inp[2]) ? node964 : node961;
													assign node961 = (inp[12]) ? 8'b10100100 : 8'b10101100;
													assign node964 = (inp[12]) ? 8'b10110001 : node965;
														assign node965 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node969 = (inp[2]) ? node975 : node970;
													assign node970 = (inp[12]) ? 8'b11111101 : node971;
														assign node971 = (inp[6]) ? 8'b10101101 : 8'b10111100;
													assign node975 = (inp[6]) ? node979 : node976;
														assign node976 = (inp[12]) ? 8'b10101101 : 8'b10111100;
														assign node979 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node982 = (inp[3]) ? node996 : node983;
												assign node983 = (inp[2]) ? node991 : node984;
													assign node984 = (inp[6]) ? node988 : node985;
														assign node985 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node988 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node991 = (inp[6]) ? node993 : 8'b10100100;
														assign node993 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node996 = (inp[2]) ? node1004 : node997;
													assign node997 = (inp[6]) ? node1001 : node998;
														assign node998 = (inp[12]) ? 8'b10100001 : 8'b10110000;
														assign node1001 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node1004 = (inp[6]) ? node1008 : node1005;
														assign node1005 = (inp[12]) ? 8'b10100001 : 8'b10110000;
														assign node1008 = (inp[12]) ? 8'b10110000 : 8'b10100000;
							assign node1011 = (inp[11]) ? node1113 : node1012;
								assign node1012 = (inp[5]) ? node1086 : node1013;
									assign node1013 = (inp[10]) ? node1047 : node1014;
										assign node1014 = (inp[2]) ? node1036 : node1015;
											assign node1015 = (inp[6]) ? node1023 : node1016;
												assign node1016 = (inp[3]) ? node1020 : node1017;
													assign node1017 = (inp[1]) ? 8'b10000101 : 8'b10000100;
													assign node1020 = (inp[1]) ? 8'b10000100 : 8'b10001101;
												assign node1023 = (inp[12]) ? node1029 : node1024;
													assign node1024 = (inp[3]) ? 8'b10011100 : node1025;
														assign node1025 = (inp[1]) ? 8'b10011101 : 8'b10011100;
													assign node1029 = (inp[1]) ? node1033 : node1030;
														assign node1030 = (inp[3]) ? 8'b10011101 : 8'b10011100;
														assign node1033 = (inp[3]) ? 8'b10011100 : 8'b10011101;
											assign node1036 = (inp[6]) ? node1040 : node1037;
												assign node1037 = (inp[3]) ? 8'b10010100 : 8'b10010101;
												assign node1040 = (inp[3]) ? node1044 : node1041;
													assign node1041 = (inp[1]) ? 8'b10000101 : 8'b10000100;
													assign node1044 = (inp[1]) ? 8'b10000100 : 8'b10001101;
										assign node1047 = (inp[1]) ? node1067 : node1048;
											assign node1048 = (inp[3]) ? node1054 : node1049;
												assign node1049 = (inp[2]) ? 8'b10010000 : node1050;
													assign node1050 = (inp[6]) ? 8'b00011010 : 8'b00000010;
												assign node1054 = (inp[12]) ? node1062 : node1055;
													assign node1055 = (inp[6]) ? node1059 : node1056;
														assign node1056 = (inp[2]) ? 8'b00011011 : 8'b00001011;
														assign node1059 = (inp[2]) ? 8'b00001011 : 8'b00011011;
													assign node1062 = (inp[6]) ? node1064 : 8'b00001011;
														assign node1064 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1067 = (inp[3]) ? node1075 : node1068;
												assign node1068 = (inp[2]) ? node1072 : node1069;
													assign node1069 = (inp[6]) ? 8'b10011001 : 8'b10000001;
													assign node1072 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node1075 = (inp[6]) ? node1081 : node1076;
													assign node1076 = (inp[2]) ? 8'b10010000 : node1077;
														assign node1077 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node1081 = (inp[2]) ? node1083 : 8'b00011010;
														assign node1083 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node1086 = (inp[6]) ? node1100 : node1087;
										assign node1087 = (inp[2]) ? node1093 : node1088;
											assign node1088 = (inp[1]) ? 8'b10000101 : node1089;
												assign node1089 = (inp[3]) ? 8'b10001101 : 8'b10000100;
											assign node1093 = (inp[3]) ? node1097 : node1094;
												assign node1094 = (inp[1]) ? 8'b10010101 : 8'b10010100;
												assign node1097 = (inp[1]) ? 8'b10010101 : 8'b10011101;
										assign node1100 = (inp[2]) ? node1106 : node1101;
											assign node1101 = (inp[1]) ? 8'b10011101 : node1102;
												assign node1102 = (inp[3]) ? 8'b10011101 : 8'b10011100;
											assign node1106 = (inp[3]) ? node1110 : node1107;
												assign node1107 = (inp[1]) ? 8'b10010101 : 8'b10010100;
												assign node1110 = (inp[1]) ? 8'b10010101 : 8'b10011101;
								assign node1113 = (inp[1]) ? node1191 : node1114;
									assign node1114 = (inp[3]) ? node1152 : node1115;
										assign node1115 = (inp[2]) ? node1133 : node1116;
											assign node1116 = (inp[6]) ? node1128 : node1117;
												assign node1117 = (inp[12]) ? node1123 : node1118;
													assign node1118 = (inp[5]) ? 8'b10110001 : node1119;
														assign node1119 = (inp[10]) ? 8'b11110111 : 8'b10110001;
													assign node1123 = (inp[10]) ? node1125 : 8'b10100100;
														assign node1125 = (inp[5]) ? 8'b10100100 : 8'b00000010;
												assign node1128 = (inp[12]) ? node1130 : 8'b10101100;
													assign node1130 = (inp[10]) ? 8'b00011010 : 8'b10111100;
											assign node1133 = (inp[5]) ? node1149 : node1134;
												assign node1134 = (inp[10]) ? node1142 : node1135;
													assign node1135 = (inp[6]) ? node1139 : node1136;
														assign node1136 = (inp[12]) ? 8'b10110001 : 8'b10100001;
														assign node1139 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node1142 = (inp[6]) ? node1146 : node1143;
														assign node1143 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node1146 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node1149 = (inp[12]) ? 8'b10110001 : 8'b10100001;
										assign node1152 = (inp[5]) ? node1180 : node1153;
											assign node1153 = (inp[10]) ? node1167 : node1154;
												assign node1154 = (inp[6]) ? node1162 : node1155;
													assign node1155 = (inp[2]) ? node1159 : node1156;
														assign node1156 = (inp[12]) ? 8'b10101101 : 8'b10111100;
														assign node1159 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node1162 = (inp[12]) ? node1164 : 8'b10101101;
														assign node1164 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node1167 = (inp[6]) ? node1175 : node1168;
													assign node1168 = (inp[12]) ? node1172 : node1169;
														assign node1169 = (inp[2]) ? 8'b00001010 : 8'b00011010;
														assign node1172 = (inp[2]) ? 8'b00011010 : 8'b00001011;
													assign node1175 = (inp[2]) ? 8'b00001011 : node1176;
														assign node1176 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node1180 = (inp[2]) ? node1188 : node1181;
												assign node1181 = (inp[12]) ? node1185 : node1182;
													assign node1182 = (inp[6]) ? 8'b10101101 : 8'b10111100;
													assign node1185 = (inp[6]) ? 8'b11111101 : 8'b10101101;
												assign node1188 = (inp[12]) ? 8'b10111100 : 8'b10101100;
									assign node1191 = (inp[2]) ? node1231 : node1192;
										assign node1192 = (inp[6]) ? node1214 : node1193;
											assign node1193 = (inp[12]) ? node1203 : node1194;
												assign node1194 = (inp[5]) ? 8'b10110000 : node1195;
													assign node1195 = (inp[10]) ? node1199 : node1196;
														assign node1196 = (inp[3]) ? 8'b10110001 : 8'b10110000;
														assign node1199 = (inp[3]) ? 8'b11110111 : 8'b10110100;
												assign node1203 = (inp[3]) ? node1209 : node1204;
													assign node1204 = (inp[10]) ? node1206 : 8'b10100001;
														assign node1206 = (inp[5]) ? 8'b10100001 : 8'b10100101;
													assign node1209 = (inp[10]) ? node1211 : 8'b10100100;
														assign node1211 = (inp[5]) ? 8'b10100001 : 8'b00000010;
											assign node1214 = (inp[12]) ? node1222 : node1215;
												assign node1215 = (inp[5]) ? 8'b10101001 : node1216;
													assign node1216 = (inp[10]) ? 8'b00001010 : node1217;
														assign node1217 = (inp[3]) ? 8'b10101100 : 8'b10101001;
												assign node1222 = (inp[5]) ? 8'b10111001 : node1223;
													assign node1223 = (inp[3]) ? node1227 : node1224;
														assign node1224 = (inp[10]) ? 8'b11111101 : 8'b10111001;
														assign node1227 = (inp[10]) ? 8'b00011010 : 8'b10111100;
										assign node1231 = (inp[5]) ? node1263 : node1232;
											assign node1232 = (inp[10]) ? node1248 : node1233;
												assign node1233 = (inp[3]) ? node1241 : node1234;
													assign node1234 = (inp[12]) ? node1238 : node1235;
														assign node1235 = (inp[6]) ? 8'b10110000 : 8'b10100000;
														assign node1238 = (inp[6]) ? 8'b10100001 : 8'b10110000;
													assign node1241 = (inp[12]) ? node1245 : node1242;
														assign node1242 = (inp[6]) ? 8'b10110001 : 8'b10100001;
														assign node1245 = (inp[6]) ? 8'b10100100 : 8'b10110001;
												assign node1248 = (inp[3]) ? node1256 : node1249;
													assign node1249 = (inp[6]) ? node1253 : node1250;
														assign node1250 = (inp[12]) ? 8'b10110100 : 8'b10100100;
														assign node1253 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node1256 = (inp[6]) ? node1260 : node1257;
														assign node1257 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node1260 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node1263 = (inp[12]) ? 8'b10110000 : 8'b10100000;
					assign node1266 = (inp[11]) ? node1558 : node1267;
						assign node1267 = (inp[6]) ? node1397 : node1268;
							assign node1268 = (inp[0]) ? node1292 : node1269;
								assign node1269 = (inp[3]) ? node1277 : node1270;
									assign node1270 = (inp[10]) ? node1272 : 8'b00101010;
										assign node1272 = (inp[5]) ? 8'b00101110 : node1273;
											assign node1273 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node1277 = (inp[10]) ? node1283 : node1278;
										assign node1278 = (inp[5]) ? 8'b00101011 : node1279;
											assign node1279 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node1283 = (inp[5]) ? 8'b00101111 : node1284;
											assign node1284 = (inp[1]) ? node1288 : node1285;
												assign node1285 = (inp[8]) ? 8'b00101011 : 8'b00101111;
												assign node1288 = (inp[8]) ? 8'b00101010 : 8'b00101110;
								assign node1292 = (inp[2]) ? node1332 : node1293;
									assign node1293 = (inp[3]) ? node1313 : node1294;
										assign node1294 = (inp[1]) ? node1304 : node1295;
											assign node1295 = (inp[10]) ? node1299 : node1296;
												assign node1296 = (inp[8]) ? 8'b00101110 : 8'b00101010;
												assign node1299 = (inp[8]) ? node1301 : 8'b00101110;
													assign node1301 = (inp[5]) ? 8'b00101110 : 8'b00101010;
											assign node1304 = (inp[8]) ? node1308 : node1305;
												assign node1305 = (inp[10]) ? 8'b00101111 : 8'b00101011;
												assign node1308 = (inp[5]) ? 8'b00101111 : node1309;
													assign node1309 = (inp[10]) ? 8'b00101011 : 8'b00101111;
										assign node1313 = (inp[5]) ? node1327 : node1314;
											assign node1314 = (inp[1]) ? node1322 : node1315;
												assign node1315 = (inp[8]) ? node1319 : node1316;
													assign node1316 = (inp[10]) ? 8'b00101111 : 8'b00101011;
													assign node1319 = (inp[10]) ? 8'b00101011 : 8'b00101111;
												assign node1322 = (inp[8]) ? node1324 : 8'b00101110;
													assign node1324 = (inp[10]) ? 8'b00101010 : 8'b00101110;
											assign node1327 = (inp[8]) ? 8'b00101111 : node1328;
												assign node1328 = (inp[10]) ? 8'b00101111 : 8'b00101011;
									assign node1332 = (inp[5]) ? node1380 : node1333;
										assign node1333 = (inp[3]) ? node1355 : node1334;
											assign node1334 = (inp[1]) ? node1342 : node1335;
												assign node1335 = (inp[10]) ? node1339 : node1336;
													assign node1336 = (inp[8]) ? 8'b00111110 : 8'b00111010;
													assign node1339 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node1342 = (inp[12]) ? node1348 : node1343;
													assign node1343 = (inp[10]) ? 8'b01111111 : node1344;
														assign node1344 = (inp[8]) ? 8'b01111111 : 8'b00111011;
													assign node1348 = (inp[10]) ? node1352 : node1349;
														assign node1349 = (inp[8]) ? 8'b01111111 : 8'b00111011;
														assign node1352 = (inp[8]) ? 8'b00111011 : 8'b01111111;
											assign node1355 = (inp[1]) ? node1365 : node1356;
												assign node1356 = (inp[12]) ? 8'b00111011 : node1357;
													assign node1357 = (inp[10]) ? node1361 : node1358;
														assign node1358 = (inp[8]) ? 8'b01111111 : 8'b00111011;
														assign node1361 = (inp[8]) ? 8'b00111011 : 8'b01111111;
												assign node1365 = (inp[12]) ? node1373 : node1366;
													assign node1366 = (inp[8]) ? node1370 : node1367;
														assign node1367 = (inp[10]) ? 8'b00111110 : 8'b00111010;
														assign node1370 = (inp[10]) ? 8'b00111010 : 8'b00111110;
													assign node1373 = (inp[10]) ? node1377 : node1374;
														assign node1374 = (inp[8]) ? 8'b00111110 : 8'b00111010;
														assign node1377 = (inp[8]) ? 8'b00111010 : 8'b00111110;
										assign node1380 = (inp[1]) ? node1392 : node1381;
											assign node1381 = (inp[3]) ? node1387 : node1382;
												assign node1382 = (inp[10]) ? 8'b00111110 : node1383;
													assign node1383 = (inp[8]) ? 8'b00111110 : 8'b00111010;
												assign node1387 = (inp[10]) ? 8'b01111111 : node1388;
													assign node1388 = (inp[8]) ? 8'b01111111 : 8'b00111011;
											assign node1392 = (inp[10]) ? 8'b01111111 : node1393;
												assign node1393 = (inp[8]) ? 8'b01111111 : 8'b00111011;
							assign node1397 = (inp[5]) ? node1535 : node1398;
								assign node1398 = (inp[2]) ? node1472 : node1399;
									assign node1399 = (inp[0]) ? node1417 : node1400;
										assign node1400 = (inp[1]) ? node1412 : node1401;
											assign node1401 = (inp[3]) ? node1407 : node1402;
												assign node1402 = (inp[8]) ? 8'b00111010 : node1403;
													assign node1403 = (inp[10]) ? 8'b00111110 : 8'b00111010;
												assign node1407 = (inp[10]) ? node1409 : 8'b00111011;
													assign node1409 = (inp[8]) ? 8'b00111011 : 8'b01111111;
											assign node1412 = (inp[8]) ? 8'b00111010 : node1413;
												assign node1413 = (inp[10]) ? 8'b00111110 : 8'b00111010;
										assign node1417 = (inp[12]) ? node1445 : node1418;
											assign node1418 = (inp[8]) ? node1434 : node1419;
												assign node1419 = (inp[10]) ? node1427 : node1420;
													assign node1420 = (inp[1]) ? node1424 : node1421;
														assign node1421 = (inp[3]) ? 8'b00111011 : 8'b00111010;
														assign node1424 = (inp[3]) ? 8'b00111010 : 8'b00111011;
													assign node1427 = (inp[1]) ? node1431 : node1428;
														assign node1428 = (inp[3]) ? 8'b01111111 : 8'b00111110;
														assign node1431 = (inp[3]) ? 8'b00111110 : 8'b01111111;
												assign node1434 = (inp[10]) ? node1440 : node1435;
													assign node1435 = (inp[1]) ? 8'b01111111 : node1436;
														assign node1436 = (inp[3]) ? 8'b01111111 : 8'b00111110;
													assign node1440 = (inp[1]) ? node1442 : 8'b00111011;
														assign node1442 = (inp[3]) ? 8'b00111010 : 8'b00111011;
											assign node1445 = (inp[3]) ? node1459 : node1446;
												assign node1446 = (inp[1]) ? node1454 : node1447;
													assign node1447 = (inp[8]) ? node1451 : node1448;
														assign node1448 = (inp[10]) ? 8'b00111110 : 8'b00111010;
														assign node1451 = (inp[10]) ? 8'b00111010 : 8'b00111110;
													assign node1454 = (inp[10]) ? node1456 : 8'b01111111;
														assign node1456 = (inp[8]) ? 8'b00111011 : 8'b01111111;
												assign node1459 = (inp[1]) ? node1465 : node1460;
													assign node1460 = (inp[8]) ? node1462 : 8'b00111011;
														assign node1462 = (inp[10]) ? 8'b00111011 : 8'b01111111;
													assign node1465 = (inp[10]) ? node1469 : node1466;
														assign node1466 = (inp[8]) ? 8'b00111110 : 8'b00111010;
														assign node1469 = (inp[8]) ? 8'b00111010 : 8'b00111110;
									assign node1472 = (inp[0]) ? node1490 : node1473;
										assign node1473 = (inp[10]) ? node1479 : node1474;
											assign node1474 = (inp[3]) ? node1476 : 8'b00101010;
												assign node1476 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node1479 = (inp[8]) ? node1485 : node1480;
												assign node1480 = (inp[1]) ? 8'b00101110 : node1481;
													assign node1481 = (inp[3]) ? 8'b00101111 : 8'b00101110;
												assign node1485 = (inp[1]) ? 8'b00101010 : node1486;
													assign node1486 = (inp[3]) ? 8'b00101011 : 8'b00101010;
										assign node1490 = (inp[3]) ? node1512 : node1491;
											assign node1491 = (inp[1]) ? node1499 : node1492;
												assign node1492 = (inp[8]) ? node1496 : node1493;
													assign node1493 = (inp[10]) ? 8'b00101110 : 8'b00101010;
													assign node1496 = (inp[10]) ? 8'b00101010 : 8'b00101110;
												assign node1499 = (inp[12]) ? node1507 : node1500;
													assign node1500 = (inp[8]) ? node1504 : node1501;
														assign node1501 = (inp[10]) ? 8'b00101111 : 8'b00101011;
														assign node1504 = (inp[10]) ? 8'b00101011 : 8'b00101111;
													assign node1507 = (inp[10]) ? node1509 : 8'b00101111;
														assign node1509 = (inp[8]) ? 8'b00101011 : 8'b00101111;
											assign node1512 = (inp[1]) ? node1520 : node1513;
												assign node1513 = (inp[10]) ? node1517 : node1514;
													assign node1514 = (inp[8]) ? 8'b00101111 : 8'b00101011;
													assign node1517 = (inp[8]) ? 8'b00101011 : 8'b00101111;
												assign node1520 = (inp[12]) ? node1528 : node1521;
													assign node1521 = (inp[8]) ? node1525 : node1522;
														assign node1522 = (inp[10]) ? 8'b00101110 : 8'b00101010;
														assign node1525 = (inp[10]) ? 8'b00101010 : 8'b00101110;
													assign node1528 = (inp[8]) ? node1532 : node1529;
														assign node1529 = (inp[10]) ? 8'b00101110 : 8'b00101010;
														assign node1532 = (inp[10]) ? 8'b00101010 : 8'b00101110;
								assign node1535 = (inp[3]) ? node1551 : node1536;
									assign node1536 = (inp[10]) ? node1546 : node1537;
										assign node1537 = (inp[0]) ? node1539 : 8'b00111010;
											assign node1539 = (inp[8]) ? node1543 : node1540;
												assign node1540 = (inp[1]) ? 8'b00111011 : 8'b00111010;
												assign node1543 = (inp[1]) ? 8'b01111111 : 8'b00111110;
										assign node1546 = (inp[1]) ? node1548 : 8'b00111110;
											assign node1548 = (inp[0]) ? 8'b01111111 : 8'b00111110;
									assign node1551 = (inp[10]) ? 8'b01111111 : node1552;
										assign node1552 = (inp[8]) ? node1554 : 8'b00111011;
											assign node1554 = (inp[0]) ? 8'b01111111 : 8'b00111011;
						assign node1558 = (inp[8]) ? node1828 : node1559;
							assign node1559 = (inp[10]) ? node1697 : node1560;
								assign node1560 = (inp[1]) ? node1616 : node1561;
									assign node1561 = (inp[3]) ? node1593 : node1562;
										assign node1562 = (inp[2]) ? node1570 : node1563;
											assign node1563 = (inp[12]) ? node1567 : node1564;
												assign node1564 = (inp[6]) ? 8'b00101010 : 8'b00011111;
												assign node1567 = (inp[6]) ? 8'b00111010 : 8'b00101010;
											assign node1570 = (inp[12]) ? node1582 : node1571;
												assign node1571 = (inp[0]) ? node1577 : node1572;
													assign node1572 = (inp[5]) ? node1574 : 8'b00011111;
														assign node1574 = (inp[6]) ? 8'b00001111 : 8'b00011111;
													assign node1577 = (inp[6]) ? node1579 : 8'b00001111;
														assign node1579 = (inp[5]) ? 8'b00001111 : 8'b00011111;
												assign node1582 = (inp[0]) ? node1588 : node1583;
													assign node1583 = (inp[6]) ? node1585 : 8'b00101010;
														assign node1585 = (inp[5]) ? 8'b00011111 : 8'b00101010;
													assign node1588 = (inp[6]) ? node1590 : 8'b00011111;
														assign node1590 = (inp[5]) ? 8'b00011111 : 8'b00101010;
										assign node1593 = (inp[2]) ? node1601 : node1594;
											assign node1594 = (inp[6]) ? node1598 : node1595;
												assign node1595 = (inp[12]) ? 8'b00101011 : 8'b00111010;
												assign node1598 = (inp[12]) ? 8'b00111011 : 8'b00101011;
											assign node1601 = (inp[12]) ? node1607 : node1602;
												assign node1602 = (inp[5]) ? node1604 : 8'b00111010;
													assign node1604 = (inp[0]) ? 8'b00101010 : 8'b00111010;
												assign node1607 = (inp[5]) ? node1611 : node1608;
													assign node1608 = (inp[6]) ? 8'b00101011 : 8'b00111010;
													assign node1611 = (inp[6]) ? 8'b00111010 : node1612;
														assign node1612 = (inp[0]) ? 8'b00111010 : 8'b00101011;
									assign node1616 = (inp[12]) ? node1658 : node1617;
										assign node1617 = (inp[6]) ? node1635 : node1618;
											assign node1618 = (inp[0]) ? node1624 : node1619;
												assign node1619 = (inp[3]) ? node1621 : 8'b00011111;
													assign node1621 = (inp[5]) ? 8'b00011110 : 8'b00011111;
												assign node1624 = (inp[2]) ? node1630 : node1625;
													assign node1625 = (inp[5]) ? 8'b00011110 : node1626;
														assign node1626 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node1630 = (inp[3]) ? node1632 : 8'b00001110;
														assign node1632 = (inp[5]) ? 8'b00001110 : 8'b00001111;
											assign node1635 = (inp[2]) ? node1647 : node1636;
												assign node1636 = (inp[0]) ? node1642 : node1637;
													assign node1637 = (inp[5]) ? node1639 : 8'b00101010;
														assign node1639 = (inp[3]) ? 8'b00001111 : 8'b00101010;
													assign node1642 = (inp[3]) ? node1644 : 8'b00001111;
														assign node1644 = (inp[5]) ? 8'b00001111 : 8'b00101010;
												assign node1647 = (inp[5]) ? node1653 : node1648;
													assign node1648 = (inp[0]) ? node1650 : 8'b00011111;
														assign node1650 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node1653 = (inp[0]) ? 8'b00001110 : node1654;
														assign node1654 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node1658 = (inp[5]) ? node1678 : node1659;
											assign node1659 = (inp[0]) ? node1665 : node1660;
												assign node1660 = (inp[2]) ? 8'b00101010 : node1661;
													assign node1661 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node1665 = (inp[3]) ? node1673 : node1666;
													assign node1666 = (inp[2]) ? node1670 : node1667;
														assign node1667 = (inp[6]) ? 8'b00011111 : 8'b00001111;
														assign node1670 = (inp[6]) ? 8'b00001111 : 8'b00011110;
													assign node1673 = (inp[6]) ? node1675 : 8'b00101010;
														assign node1675 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node1678 = (inp[6]) ? node1686 : node1679;
												assign node1679 = (inp[0]) ? node1683 : node1680;
													assign node1680 = (inp[3]) ? 8'b00001111 : 8'b00101010;
													assign node1683 = (inp[2]) ? 8'b00011110 : 8'b00001111;
												assign node1686 = (inp[2]) ? node1692 : node1687;
													assign node1687 = (inp[0]) ? 8'b00011111 : node1688;
														assign node1688 = (inp[3]) ? 8'b00011111 : 8'b00111010;
													assign node1692 = (inp[0]) ? 8'b00011110 : node1693;
														assign node1693 = (inp[3]) ? 8'b00011110 : 8'b00011111;
								assign node1697 = (inp[1]) ? node1757 : node1698;
									assign node1698 = (inp[3]) ? node1726 : node1699;
										assign node1699 = (inp[2]) ? node1707 : node1700;
											assign node1700 = (inp[12]) ? node1704 : node1701;
												assign node1701 = (inp[6]) ? 8'b00101110 : 8'b00111011;
												assign node1704 = (inp[6]) ? 8'b00111110 : 8'b00101110;
											assign node1707 = (inp[12]) ? node1715 : node1708;
												assign node1708 = (inp[0]) ? 8'b00101011 : node1709;
													assign node1709 = (inp[6]) ? node1711 : 8'b00111011;
														assign node1711 = (inp[5]) ? 8'b00101011 : 8'b00111011;
												assign node1715 = (inp[0]) ? node1721 : node1716;
													assign node1716 = (inp[6]) ? node1718 : 8'b00101110;
														assign node1718 = (inp[5]) ? 8'b00111011 : 8'b00101110;
													assign node1721 = (inp[6]) ? node1723 : 8'b00111011;
														assign node1723 = (inp[5]) ? 8'b00111011 : 8'b00101110;
										assign node1726 = (inp[2]) ? node1734 : node1727;
											assign node1727 = (inp[6]) ? node1731 : node1728;
												assign node1728 = (inp[12]) ? 8'b00101111 : 8'b00111110;
												assign node1731 = (inp[12]) ? 8'b01111111 : 8'b00101111;
											assign node1734 = (inp[12]) ? node1746 : node1735;
												assign node1735 = (inp[0]) ? node1741 : node1736;
													assign node1736 = (inp[5]) ? node1738 : 8'b00111110;
														assign node1738 = (inp[6]) ? 8'b00101110 : 8'b00111110;
													assign node1741 = (inp[5]) ? 8'b00101110 : node1742;
														assign node1742 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node1746 = (inp[0]) ? node1752 : node1747;
													assign node1747 = (inp[5]) ? node1749 : 8'b00101111;
														assign node1749 = (inp[6]) ? 8'b00111110 : 8'b00101111;
													assign node1752 = (inp[6]) ? node1754 : 8'b00111110;
														assign node1754 = (inp[5]) ? 8'b00111110 : 8'b00101111;
									assign node1757 = (inp[12]) ? node1793 : node1758;
										assign node1758 = (inp[6]) ? node1774 : node1759;
											assign node1759 = (inp[0]) ? node1765 : node1760;
												assign node1760 = (inp[3]) ? node1762 : 8'b00111011;
													assign node1762 = (inp[5]) ? 8'b00111010 : 8'b00111011;
												assign node1765 = (inp[2]) ? node1769 : node1766;
													assign node1766 = (inp[5]) ? 8'b00111010 : 8'b00111011;
													assign node1769 = (inp[3]) ? node1771 : 8'b00101010;
														assign node1771 = (inp[5]) ? 8'b00101010 : 8'b00101011;
											assign node1774 = (inp[2]) ? node1786 : node1775;
												assign node1775 = (inp[5]) ? node1781 : node1776;
													assign node1776 = (inp[0]) ? node1778 : 8'b00101110;
														assign node1778 = (inp[3]) ? 8'b00101110 : 8'b00101011;
													assign node1781 = (inp[3]) ? 8'b00101011 : node1782;
														assign node1782 = (inp[0]) ? 8'b00101011 : 8'b00101110;
												assign node1786 = (inp[5]) ? 8'b00101010 : node1787;
													assign node1787 = (inp[3]) ? 8'b00111011 : node1788;
														assign node1788 = (inp[0]) ? 8'b00111010 : 8'b00111011;
										assign node1793 = (inp[0]) ? node1811 : node1794;
											assign node1794 = (inp[5]) ? node1800 : node1795;
												assign node1795 = (inp[2]) ? 8'b00101110 : node1796;
													assign node1796 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node1800 = (inp[6]) ? node1804 : node1801;
													assign node1801 = (inp[3]) ? 8'b00101011 : 8'b00101110;
													assign node1804 = (inp[3]) ? node1808 : node1805;
														assign node1805 = (inp[2]) ? 8'b00111011 : 8'b00111110;
														assign node1808 = (inp[2]) ? 8'b00111010 : 8'b00111011;
											assign node1811 = (inp[2]) ? node1819 : node1812;
												assign node1812 = (inp[6]) ? node1814 : 8'b00101011;
													assign node1814 = (inp[5]) ? 8'b00111011 : node1815;
														assign node1815 = (inp[3]) ? 8'b00111110 : 8'b00111011;
												assign node1819 = (inp[5]) ? 8'b00111010 : node1820;
													assign node1820 = (inp[6]) ? node1824 : node1821;
														assign node1821 = (inp[3]) ? 8'b00111011 : 8'b00111010;
														assign node1824 = (inp[3]) ? 8'b00101110 : 8'b00101011;
							assign node1828 = (inp[0]) ? node1932 : node1829;
								assign node1829 = (inp[12]) ? node1879 : node1830;
									assign node1830 = (inp[6]) ? node1848 : node1831;
										assign node1831 = (inp[3]) ? node1837 : node1832;
											assign node1832 = (inp[10]) ? node1834 : 8'b00011111;
												assign node1834 = (inp[5]) ? 8'b00011011 : 8'b00011111;
											assign node1837 = (inp[1]) ? node1843 : node1838;
												assign node1838 = (inp[5]) ? node1840 : 8'b00111010;
													assign node1840 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node1843 = (inp[5]) ? node1845 : 8'b00011111;
													assign node1845 = (inp[10]) ? 8'b00011010 : 8'b00011110;
										assign node1848 = (inp[2]) ? node1866 : node1849;
											assign node1849 = (inp[5]) ? node1855 : node1850;
												assign node1850 = (inp[1]) ? 8'b00101010 : node1851;
													assign node1851 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node1855 = (inp[3]) ? node1859 : node1856;
													assign node1856 = (inp[10]) ? 8'b00001110 : 8'b00101010;
													assign node1859 = (inp[1]) ? node1863 : node1860;
														assign node1860 = (inp[10]) ? 8'b00001111 : 8'b00101011;
														assign node1863 = (inp[10]) ? 8'b00001011 : 8'b00001111;
											assign node1866 = (inp[5]) ? node1872 : node1867;
												assign node1867 = (inp[1]) ? 8'b00011111 : node1868;
													assign node1868 = (inp[3]) ? 8'b00111010 : 8'b00011111;
												assign node1872 = (inp[3]) ? node1876 : node1873;
													assign node1873 = (inp[10]) ? 8'b00001011 : 8'b00001111;
													assign node1876 = (inp[1]) ? 8'b00001010 : 8'b00101010;
									assign node1879 = (inp[5]) ? node1897 : node1880;
										assign node1880 = (inp[6]) ? node1886 : node1881;
											assign node1881 = (inp[1]) ? 8'b00101010 : node1882;
												assign node1882 = (inp[3]) ? 8'b00101011 : 8'b00101010;
											assign node1886 = (inp[2]) ? node1892 : node1887;
												assign node1887 = (inp[1]) ? 8'b00111010 : node1888;
													assign node1888 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node1892 = (inp[1]) ? 8'b00101010 : node1893;
													assign node1893 = (inp[3]) ? 8'b00101011 : 8'b00101010;
										assign node1897 = (inp[6]) ? node1909 : node1898;
											assign node1898 = (inp[10]) ? node1904 : node1899;
												assign node1899 = (inp[3]) ? node1901 : 8'b00101010;
													assign node1901 = (inp[1]) ? 8'b00001111 : 8'b00101011;
												assign node1904 = (inp[3]) ? node1906 : 8'b00001110;
													assign node1906 = (inp[1]) ? 8'b00001011 : 8'b00001111;
											assign node1909 = (inp[10]) ? node1925 : node1910;
												assign node1910 = (inp[1]) ? node1918 : node1911;
													assign node1911 = (inp[3]) ? node1915 : node1912;
														assign node1912 = (inp[2]) ? 8'b00011111 : 8'b00111010;
														assign node1915 = (inp[2]) ? 8'b00111010 : 8'b00111011;
													assign node1918 = (inp[3]) ? node1922 : node1919;
														assign node1919 = (inp[2]) ? 8'b00011111 : 8'b00111010;
														assign node1922 = (inp[2]) ? 8'b00011110 : 8'b00011111;
												assign node1925 = (inp[2]) ? node1929 : node1926;
													assign node1926 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node1929 = (inp[3]) ? 8'b00011110 : 8'b00011011;
								assign node1932 = (inp[1]) ? node2024 : node1933;
									assign node1933 = (inp[10]) ? node1973 : node1934;
										assign node1934 = (inp[3]) ? node1954 : node1935;
											assign node1935 = (inp[2]) ? node1943 : node1936;
												assign node1936 = (inp[12]) ? node1940 : node1937;
													assign node1937 = (inp[6]) ? 8'b00001110 : 8'b00011011;
													assign node1940 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node1943 = (inp[12]) ? node1949 : node1944;
													assign node1944 = (inp[6]) ? node1946 : 8'b00001011;
														assign node1946 = (inp[5]) ? 8'b00001011 : 8'b00011011;
													assign node1949 = (inp[5]) ? 8'b00011011 : node1950;
														assign node1950 = (inp[6]) ? 8'b00001110 : 8'b00011011;
											assign node1954 = (inp[2]) ? node1962 : node1955;
												assign node1955 = (inp[12]) ? node1959 : node1956;
													assign node1956 = (inp[6]) ? 8'b00001111 : 8'b00011110;
													assign node1959 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node1962 = (inp[12]) ? node1968 : node1963;
													assign node1963 = (inp[6]) ? node1965 : 8'b00001110;
														assign node1965 = (inp[5]) ? 8'b00001110 : 8'b00011110;
													assign node1968 = (inp[6]) ? node1970 : 8'b00011110;
														assign node1970 = (inp[5]) ? 8'b00011110 : 8'b00001111;
										assign node1973 = (inp[5]) ? node2003 : node1974;
											assign node1974 = (inp[3]) ? node1990 : node1975;
												assign node1975 = (inp[6]) ? node1983 : node1976;
													assign node1976 = (inp[2]) ? node1980 : node1977;
														assign node1977 = (inp[12]) ? 8'b00101010 : 8'b00011111;
														assign node1980 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node1983 = (inp[2]) ? node1987 : node1984;
														assign node1984 = (inp[12]) ? 8'b00111010 : 8'b00101010;
														assign node1987 = (inp[12]) ? 8'b00101010 : 8'b00011111;
												assign node1990 = (inp[12]) ? node1998 : node1991;
													assign node1991 = (inp[2]) ? node1995 : node1992;
														assign node1992 = (inp[6]) ? 8'b00101011 : 8'b00111010;
														assign node1995 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node1998 = (inp[2]) ? 8'b00101011 : node1999;
														assign node1999 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node2003 = (inp[3]) ? node2015 : node2004;
												assign node2004 = (inp[2]) ? node2012 : node2005;
													assign node2005 = (inp[12]) ? node2009 : node2006;
														assign node2006 = (inp[6]) ? 8'b00001110 : 8'b00011011;
														assign node2009 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node2012 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2015 = (inp[2]) ? node2021 : node2016;
													assign node2016 = (inp[12]) ? 8'b00001111 : node2017;
														assign node2017 = (inp[6]) ? 8'b00001111 : 8'b00011110;
													assign node2021 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node2024 = (inp[5]) ? node2080 : node2025;
										assign node2025 = (inp[10]) ? node2051 : node2026;
											assign node2026 = (inp[3]) ? node2042 : node2027;
												assign node2027 = (inp[6]) ? node2035 : node2028;
													assign node2028 = (inp[2]) ? node2032 : node2029;
														assign node2029 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node2032 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2035 = (inp[12]) ? node2039 : node2036;
														assign node2036 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node2039 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node2042 = (inp[6]) ? node2044 : 8'b00011011;
													assign node2044 = (inp[12]) ? node2048 : node2045;
														assign node2045 = (inp[2]) ? 8'b00011011 : 8'b00001110;
														assign node2048 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node2051 = (inp[3]) ? node2065 : node2052;
												assign node2052 = (inp[12]) ? node2060 : node2053;
													assign node2053 = (inp[6]) ? node2057 : node2054;
														assign node2054 = (inp[2]) ? 8'b00001110 : 8'b00011110;
														assign node2057 = (inp[2]) ? 8'b00011110 : 8'b00001111;
													assign node2060 = (inp[6]) ? node2062 : 8'b00001111;
														assign node2062 = (inp[2]) ? 8'b00001111 : 8'b00011111;
												assign node2065 = (inp[2]) ? node2073 : node2066;
													assign node2066 = (inp[6]) ? node2070 : node2067;
														assign node2067 = (inp[12]) ? 8'b00101010 : 8'b00011111;
														assign node2070 = (inp[12]) ? 8'b00111010 : 8'b00101010;
													assign node2073 = (inp[12]) ? node2077 : node2074;
														assign node2074 = (inp[6]) ? 8'b00011111 : 8'b00001111;
														assign node2077 = (inp[6]) ? 8'b00101010 : 8'b00011111;
										assign node2080 = (inp[2]) ? node2088 : node2081;
											assign node2081 = (inp[6]) ? node2085 : node2082;
												assign node2082 = (inp[12]) ? 8'b00001011 : 8'b00011010;
												assign node2085 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node2088 = (inp[12]) ? 8'b00011010 : 8'b00001010;
			assign node2091 = (inp[0]) ? node3103 : node2092;
				assign node2092 = (inp[5]) ? node2290 : node2093;
					assign node2093 = (inp[8]) ? node2219 : node2094;
						assign node2094 = (inp[4]) ? node2118 : node2095;
							assign node2095 = (inp[1]) ? node2107 : node2096;
								assign node2096 = (inp[2]) ? node2102 : node2097;
									assign node2097 = (inp[12]) ? 8'b00011111 : node2098;
										assign node2098 = (inp[11]) ? 8'b00001111 : 8'b00011111;
									assign node2102 = (inp[11]) ? node2104 : 8'b00001111;
										assign node2104 = (inp[12]) ? 8'b00001111 : 8'b00011110;
								assign node2107 = (inp[2]) ? node2113 : node2108;
									assign node2108 = (inp[12]) ? 8'b00011110 : node2109;
										assign node2109 = (inp[11]) ? 8'b00001110 : 8'b00011110;
									assign node2113 = (inp[11]) ? node2115 : 8'b00001110;
										assign node2115 = (inp[12]) ? 8'b00001110 : 8'b00011011;
							assign node2118 = (inp[10]) ? node2168 : node2119;
								assign node2119 = (inp[12]) ? node2151 : node2120;
									assign node2120 = (inp[11]) ? node2134 : node2121;
										assign node2121 = (inp[2]) ? node2129 : node2122;
											assign node2122 = (inp[6]) ? node2124 : 8'b10000010;
												assign node2124 = (inp[1]) ? 8'b00011010 : node2125;
													assign node2125 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node2129 = (inp[3]) ? node2131 : 8'b10000010;
												assign node2131 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node2134 = (inp[3]) ? node2140 : node2135;
											assign node2135 = (inp[2]) ? 8'b11110111 : node2136;
												assign node2136 = (inp[6]) ? 8'b00001010 : 8'b11110111;
											assign node2140 = (inp[1]) ? node2146 : node2141;
												assign node2141 = (inp[6]) ? node2143 : 8'b00011010;
													assign node2143 = (inp[2]) ? 8'b00011010 : 8'b00001011;
												assign node2146 = (inp[2]) ? 8'b11110111 : node2147;
													assign node2147 = (inp[6]) ? 8'b00001010 : 8'b11110111;
									assign node2151 = (inp[6]) ? node2157 : node2152;
										assign node2152 = (inp[1]) ? 8'b00000010 : node2153;
											assign node2153 = (inp[3]) ? 8'b00001011 : 8'b00000010;
										assign node2157 = (inp[2]) ? node2163 : node2158;
											assign node2158 = (inp[1]) ? 8'b00011010 : node2159;
												assign node2159 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node2163 = (inp[1]) ? 8'b00000010 : node2164;
												assign node2164 = (inp[3]) ? 8'b00001011 : 8'b00000010;
								assign node2168 = (inp[12]) ? node2202 : node2169;
									assign node2169 = (inp[11]) ? node2185 : node2170;
										assign node2170 = (inp[6]) ? node2176 : node2171;
											assign node2171 = (inp[1]) ? 8'b00001110 : node2172;
												assign node2172 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node2176 = (inp[2]) ? node2182 : node2177;
												assign node2177 = (inp[3]) ? node2179 : 8'b00011110;
													assign node2179 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node2182 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node2185 = (inp[2]) ? node2197 : node2186;
											assign node2186 = (inp[6]) ? node2192 : node2187;
												assign node2187 = (inp[1]) ? 8'b00011011 : node2188;
													assign node2188 = (inp[3]) ? 8'b00011110 : 8'b00011011;
												assign node2192 = (inp[3]) ? node2194 : 8'b00001110;
													assign node2194 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node2197 = (inp[3]) ? node2199 : 8'b00011011;
												assign node2199 = (inp[1]) ? 8'b00011011 : 8'b00011110;
									assign node2202 = (inp[2]) ? node2214 : node2203;
										assign node2203 = (inp[6]) ? node2209 : node2204;
											assign node2204 = (inp[3]) ? node2206 : 8'b00001110;
												assign node2206 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node2209 = (inp[3]) ? node2211 : 8'b00011110;
												assign node2211 = (inp[1]) ? 8'b00011110 : 8'b00011111;
										assign node2214 = (inp[3]) ? node2216 : 8'b00001110;
											assign node2216 = (inp[1]) ? 8'b00001110 : 8'b00001111;
						assign node2219 = (inp[1]) ? node2267 : node2220;
							assign node2220 = (inp[4]) ? node2232 : node2221;
								assign node2221 = (inp[2]) ? node2227 : node2222;
									assign node2222 = (inp[12]) ? 8'b00011011 : node2223;
										assign node2223 = (inp[11]) ? 8'b00001011 : 8'b00011011;
									assign node2227 = (inp[12]) ? 8'b00001011 : node2228;
										assign node2228 = (inp[11]) ? 8'b00011010 : 8'b00001011;
								assign node2232 = (inp[3]) ? node2250 : node2233;
									assign node2233 = (inp[12]) ? node2245 : node2234;
										assign node2234 = (inp[11]) ? node2240 : node2235;
											assign node2235 = (inp[6]) ? node2237 : 8'b10000010;
												assign node2237 = (inp[2]) ? 8'b10000010 : 8'b00011010;
											assign node2240 = (inp[6]) ? node2242 : 8'b11110111;
												assign node2242 = (inp[2]) ? 8'b11110111 : 8'b00001010;
										assign node2245 = (inp[2]) ? 8'b00000010 : node2246;
											assign node2246 = (inp[6]) ? 8'b00011010 : 8'b00000010;
									assign node2250 = (inp[11]) ? node2256 : node2251;
										assign node2251 = (inp[6]) ? node2253 : 8'b00001011;
											assign node2253 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node2256 = (inp[12]) ? node2262 : node2257;
											assign node2257 = (inp[6]) ? node2259 : 8'b00011010;
												assign node2259 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node2262 = (inp[6]) ? node2264 : 8'b00001011;
												assign node2264 = (inp[2]) ? 8'b00001011 : 8'b00011011;
							assign node2267 = (inp[2]) ? node2285 : node2268;
								assign node2268 = (inp[4]) ? node2274 : node2269;
									assign node2269 = (inp[12]) ? 8'b00011010 : node2270;
										assign node2270 = (inp[11]) ? 8'b00001010 : 8'b00011010;
									assign node2274 = (inp[6]) ? node2280 : node2275;
										assign node2275 = (inp[12]) ? 8'b00000010 : node2276;
											assign node2276 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node2280 = (inp[12]) ? 8'b00011010 : node2281;
											assign node2281 = (inp[11]) ? 8'b00001010 : 8'b00011010;
								assign node2285 = (inp[12]) ? 8'b00000010 : node2286;
									assign node2286 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node2290 = (inp[9]) ? node2698 : node2291;
						assign node2291 = (inp[8]) ? node2475 : node2292;
							assign node2292 = (inp[4]) ? node2346 : node2293;
								assign node2293 = (inp[11]) ? node2311 : node2294;
									assign node2294 = (inp[6]) ? node2306 : node2295;
										assign node2295 = (inp[2]) ? node2301 : node2296;
											assign node2296 = (inp[3]) ? 8'b00011111 : node2297;
												assign node2297 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node2301 = (inp[1]) ? node2303 : 8'b00001111;
												assign node2303 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node2306 = (inp[1]) ? node2308 : 8'b00011111;
											assign node2308 = (inp[3]) ? 8'b00011111 : 8'b00011110;
									assign node2311 = (inp[1]) ? node2323 : node2312;
										assign node2312 = (inp[2]) ? node2316 : node2313;
											assign node2313 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node2316 = (inp[12]) ? node2320 : node2317;
												assign node2317 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node2320 = (inp[6]) ? 8'b00011110 : 8'b00001111;
										assign node2323 = (inp[3]) ? node2335 : node2324;
											assign node2324 = (inp[2]) ? node2328 : node2325;
												assign node2325 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2328 = (inp[12]) ? node2332 : node2329;
													assign node2329 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node2332 = (inp[6]) ? 8'b00011011 : 8'b00001110;
											assign node2335 = (inp[2]) ? node2339 : node2336;
												assign node2336 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2339 = (inp[12]) ? node2343 : node2340;
													assign node2340 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node2343 = (inp[6]) ? 8'b00011010 : 8'b00001011;
								assign node2346 = (inp[10]) ? node2418 : node2347;
									assign node2347 = (inp[11]) ? node2365 : node2348;
										assign node2348 = (inp[6]) ? node2356 : node2349;
											assign node2349 = (inp[3]) ? node2353 : node2350;
												assign node2350 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node2353 = (inp[1]) ? 8'b10000001 : 8'b00001011;
											assign node2356 = (inp[3]) ? node2360 : node2357;
												assign node2357 = (inp[2]) ? 8'b10010000 : 8'b00011010;
												assign node2360 = (inp[1]) ? node2362 : 8'b00011011;
													assign node2362 = (inp[2]) ? 8'b10010001 : 8'b10011001;
										assign node2365 = (inp[1]) ? node2389 : node2366;
											assign node2366 = (inp[3]) ? node2376 : node2367;
												assign node2367 = (inp[6]) ? node2371 : node2368;
													assign node2368 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node2371 = (inp[2]) ? node2373 : 8'b00001010;
														assign node2373 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node2376 = (inp[2]) ? node2384 : node2377;
													assign node2377 = (inp[6]) ? node2381 : node2378;
														assign node2378 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node2381 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node2384 = (inp[12]) ? node2386 : 8'b00011010;
														assign node2386 = (inp[6]) ? 8'b00011010 : 8'b00001011;
											assign node2389 = (inp[3]) ? node2403 : node2390;
												assign node2390 = (inp[2]) ? node2396 : node2391;
													assign node2391 = (inp[6]) ? node2393 : 8'b00000010;
														assign node2393 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2396 = (inp[6]) ? node2400 : node2397;
														assign node2397 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node2400 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node2403 = (inp[2]) ? node2411 : node2404;
													assign node2404 = (inp[6]) ? node2408 : node2405;
														assign node2405 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node2408 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node2411 = (inp[12]) ? node2415 : node2412;
														assign node2412 = (inp[6]) ? 8'b10100100 : 8'b10110100;
														assign node2415 = (inp[6]) ? 8'b10110100 : 8'b10100101;
									assign node2418 = (inp[11]) ? node2426 : node2419;
										assign node2419 = (inp[3]) ? node2423 : node2420;
											assign node2420 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node2423 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node2426 = (inp[1]) ? node2452 : node2427;
											assign node2427 = (inp[3]) ? node2441 : node2428;
												assign node2428 = (inp[2]) ? node2436 : node2429;
													assign node2429 = (inp[6]) ? node2433 : node2430;
														assign node2430 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node2433 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node2436 = (inp[12]) ? 8'b00011011 : node2437;
														assign node2437 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node2441 = (inp[12]) ? node2447 : node2442;
													assign node2442 = (inp[6]) ? node2444 : 8'b00011110;
														assign node2444 = (inp[2]) ? 8'b00001110 : 8'b00001111;
													assign node2447 = (inp[6]) ? node2449 : 8'b00001111;
														assign node2449 = (inp[2]) ? 8'b00011110 : 8'b00011111;
											assign node2452 = (inp[3]) ? node2464 : node2453;
												assign node2453 = (inp[12]) ? node2459 : node2454;
													assign node2454 = (inp[6]) ? node2456 : 8'b00011011;
														assign node2456 = (inp[2]) ? 8'b00001011 : 8'b00001110;
													assign node2459 = (inp[6]) ? node2461 : 8'b00001110;
														assign node2461 = (inp[2]) ? 8'b00011011 : 8'b00011110;
												assign node2464 = (inp[12]) ? node2470 : node2465;
													assign node2465 = (inp[6]) ? node2467 : 8'b00011010;
														assign node2467 = (inp[2]) ? 8'b00001010 : 8'b00001011;
													assign node2470 = (inp[6]) ? node2472 : 8'b00001011;
														assign node2472 = (inp[2]) ? 8'b00011010 : 8'b00011011;
							assign node2475 = (inp[10]) ? node2587 : node2476;
								assign node2476 = (inp[1]) ? node2526 : node2477;
									assign node2477 = (inp[4]) ? node2495 : node2478;
										assign node2478 = (inp[11]) ? node2484 : node2479;
											assign node2479 = (inp[6]) ? 8'b00011011 : node2480;
												assign node2480 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node2484 = (inp[2]) ? node2488 : node2485;
												assign node2485 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2488 = (inp[6]) ? node2492 : node2489;
													assign node2489 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node2492 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node2495 = (inp[3]) ? node2511 : node2496;
											assign node2496 = (inp[6]) ? node2502 : node2497;
												assign node2497 = (inp[12]) ? 8'b00000010 : node2498;
													assign node2498 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node2502 = (inp[2]) ? node2508 : node2503;
													assign node2503 = (inp[11]) ? node2505 : 8'b00011010;
														assign node2505 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2508 = (inp[11]) ? 8'b11110101 : 8'b10010000;
											assign node2511 = (inp[11]) ? node2515 : node2512;
												assign node2512 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node2515 = (inp[12]) ? node2521 : node2516;
													assign node2516 = (inp[6]) ? node2518 : 8'b00011010;
														assign node2518 = (inp[2]) ? 8'b00001010 : 8'b00001011;
													assign node2521 = (inp[6]) ? node2523 : 8'b00001011;
														assign node2523 = (inp[2]) ? 8'b00011010 : 8'b00011011;
									assign node2526 = (inp[3]) ? node2558 : node2527;
										assign node2527 = (inp[2]) ? node2545 : node2528;
											assign node2528 = (inp[6]) ? node2540 : node2529;
												assign node2529 = (inp[4]) ? node2535 : node2530;
													assign node2530 = (inp[12]) ? 8'b00011010 : node2531;
														assign node2531 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node2535 = (inp[12]) ? 8'b00000010 : node2536;
														assign node2536 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node2540 = (inp[11]) ? node2542 : 8'b00011010;
													assign node2542 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node2545 = (inp[11]) ? node2551 : node2546;
												assign node2546 = (inp[6]) ? 8'b10010000 : node2547;
													assign node2547 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node2551 = (inp[6]) ? node2555 : node2552;
													assign node2552 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node2555 = (inp[12]) ? 8'b11110101 : 8'b10100101;
										assign node2558 = (inp[11]) ? node2568 : node2559;
											assign node2559 = (inp[6]) ? node2565 : node2560;
												assign node2560 = (inp[4]) ? 8'b10000001 : node2561;
													assign node2561 = (inp[2]) ? 8'b10000001 : 8'b10011001;
												assign node2565 = (inp[2]) ? 8'b10010001 : 8'b10011001;
											assign node2568 = (inp[2]) ? node2580 : node2569;
												assign node2569 = (inp[12]) ? node2575 : node2570;
													assign node2570 = (inp[4]) ? node2572 : 8'b10101101;
														assign node2572 = (inp[6]) ? 8'b10101101 : 8'b10110100;
													assign node2575 = (inp[6]) ? 8'b11111101 : node2576;
														assign node2576 = (inp[4]) ? 8'b10100101 : 8'b11111101;
												assign node2580 = (inp[6]) ? node2584 : node2581;
													assign node2581 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node2584 = (inp[12]) ? 8'b10110100 : 8'b10100100;
								assign node2587 = (inp[11]) ? node2625 : node2588;
									assign node2588 = (inp[3]) ? node2608 : node2589;
										assign node2589 = (inp[6]) ? node2597 : node2590;
											assign node2590 = (inp[4]) ? 8'b10000100 : node2591;
												assign node2591 = (inp[2]) ? 8'b10000100 : node2592;
													assign node2592 = (inp[1]) ? 8'b10011100 : 8'b10011101;
											assign node2597 = (inp[2]) ? node2603 : node2598;
												assign node2598 = (inp[4]) ? 8'b10011100 : node2599;
													assign node2599 = (inp[1]) ? 8'b10011100 : 8'b10011101;
												assign node2603 = (inp[1]) ? 8'b10010100 : node2604;
													assign node2604 = (inp[4]) ? 8'b10010100 : 8'b10011101;
										assign node2608 = (inp[6]) ? node2620 : node2609;
											assign node2609 = (inp[1]) ? node2615 : node2610;
												assign node2610 = (inp[4]) ? 8'b10001101 : node2611;
													assign node2611 = (inp[2]) ? 8'b10001101 : 8'b10011101;
												assign node2615 = (inp[4]) ? 8'b10000101 : node2616;
													assign node2616 = (inp[2]) ? 8'b10000101 : 8'b10011101;
											assign node2620 = (inp[2]) ? node2622 : 8'b10011101;
												assign node2622 = (inp[1]) ? 8'b10010101 : 8'b10011101;
									assign node2625 = (inp[1]) ? node2661 : node2626;
										assign node2626 = (inp[4]) ? node2638 : node2627;
											assign node2627 = (inp[2]) ? node2631 : node2628;
												assign node2628 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node2631 = (inp[6]) ? node2635 : node2632;
													assign node2632 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node2635 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node2638 = (inp[3]) ? node2652 : node2639;
												assign node2639 = (inp[2]) ? node2647 : node2640;
													assign node2640 = (inp[6]) ? node2644 : node2641;
														assign node2641 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node2644 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node2647 = (inp[12]) ? 8'b10110001 : node2648;
														assign node2648 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node2652 = (inp[12]) ? node2658 : node2653;
													assign node2653 = (inp[6]) ? node2655 : 8'b10111100;
														assign node2655 = (inp[2]) ? 8'b10101100 : 8'b10101101;
													assign node2658 = (inp[6]) ? 8'b11111101 : 8'b10101101;
										assign node2661 = (inp[2]) ? node2683 : node2662;
											assign node2662 = (inp[3]) ? node2672 : node2663;
												assign node2663 = (inp[4]) ? node2667 : node2664;
													assign node2664 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node2667 = (inp[12]) ? node2669 : 8'b10110001;
														assign node2669 = (inp[6]) ? 8'b10111100 : 8'b10100100;
												assign node2672 = (inp[6]) ? node2680 : node2673;
													assign node2673 = (inp[4]) ? node2677 : node2674;
														assign node2674 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node2677 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node2680 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node2683 = (inp[3]) ? node2691 : node2684;
												assign node2684 = (inp[6]) ? node2688 : node2685;
													assign node2685 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node2688 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node2691 = (inp[6]) ? node2695 : node2692;
													assign node2692 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node2695 = (inp[12]) ? 8'b10110000 : 8'b10100000;
						assign node2698 = (inp[11]) ? node2804 : node2699;
							assign node2699 = (inp[10]) ? node2757 : node2700;
								assign node2700 = (inp[3]) ? node2730 : node2701;
									assign node2701 = (inp[4]) ? node2725 : node2702;
										assign node2702 = (inp[8]) ? node2714 : node2703;
											assign node2703 = (inp[1]) ? node2709 : node2704;
												assign node2704 = (inp[2]) ? node2706 : 8'b11111101;
													assign node2706 = (inp[6]) ? 8'b11111101 : 8'b10101101;
												assign node2709 = (inp[2]) ? node2711 : 8'b10111100;
													assign node2711 = (inp[6]) ? 8'b10111100 : 8'b10101100;
											assign node2714 = (inp[1]) ? node2720 : node2715;
												assign node2715 = (inp[2]) ? node2717 : 8'b10111001;
													assign node2717 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node2720 = (inp[2]) ? node2722 : 8'b10111000;
													assign node2722 = (inp[6]) ? 8'b10110000 : 8'b10100000;
										assign node2725 = (inp[6]) ? node2727 : 8'b10100000;
											assign node2727 = (inp[2]) ? 8'b10110000 : 8'b10111000;
									assign node2730 = (inp[6]) ? node2744 : node2731;
										assign node2731 = (inp[4]) ? node2741 : node2732;
											assign node2732 = (inp[8]) ? node2736 : node2733;
												assign node2733 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node2736 = (inp[2]) ? node2738 : 8'b10111001;
													assign node2738 = (inp[1]) ? 8'b10100001 : 8'b10101001;
											assign node2741 = (inp[1]) ? 8'b10100001 : 8'b10101001;
										assign node2744 = (inp[8]) ? node2752 : node2745;
											assign node2745 = (inp[4]) ? node2747 : 8'b11111101;
												assign node2747 = (inp[2]) ? node2749 : 8'b10111001;
													assign node2749 = (inp[1]) ? 8'b10110001 : 8'b10111001;
											assign node2752 = (inp[2]) ? node2754 : 8'b10111001;
												assign node2754 = (inp[1]) ? 8'b10110001 : 8'b10111001;
								assign node2757 = (inp[3]) ? node2783 : node2758;
									assign node2758 = (inp[4]) ? node2774 : node2759;
										assign node2759 = (inp[1]) ? node2765 : node2760;
											assign node2760 = (inp[6]) ? 8'b11111101 : node2761;
												assign node2761 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node2765 = (inp[2]) ? node2767 : 8'b10111100;
												assign node2767 = (inp[8]) ? node2771 : node2768;
													assign node2768 = (inp[6]) ? 8'b10111100 : 8'b10101100;
													assign node2771 = (inp[6]) ? 8'b10110100 : 8'b10100100;
										assign node2774 = (inp[6]) ? node2778 : node2775;
											assign node2775 = (inp[8]) ? 8'b10100100 : 8'b10101100;
											assign node2778 = (inp[2]) ? node2780 : 8'b10111100;
												assign node2780 = (inp[8]) ? 8'b10110100 : 8'b10111100;
									assign node2783 = (inp[6]) ? node2797 : node2784;
										assign node2784 = (inp[2]) ? node2792 : node2785;
											assign node2785 = (inp[4]) ? node2787 : 8'b11111101;
												assign node2787 = (inp[8]) ? node2789 : 8'b10101101;
													assign node2789 = (inp[1]) ? 8'b10100101 : 8'b10101101;
											assign node2792 = (inp[1]) ? node2794 : 8'b10101101;
												assign node2794 = (inp[8]) ? 8'b10100101 : 8'b10101101;
										assign node2797 = (inp[8]) ? node2799 : 8'b11111101;
											assign node2799 = (inp[1]) ? node2801 : 8'b11111101;
												assign node2801 = (inp[2]) ? 8'b11110101 : 8'b11111101;
							assign node2804 = (inp[8]) ? node2952 : node2805;
								assign node2805 = (inp[4]) ? node2841 : node2806;
									assign node2806 = (inp[1]) ? node2818 : node2807;
										assign node2807 = (inp[2]) ? node2811 : node2808;
											assign node2808 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node2811 = (inp[12]) ? node2815 : node2812;
												assign node2812 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node2815 = (inp[6]) ? 8'b10111100 : 8'b10101101;
										assign node2818 = (inp[3]) ? node2830 : node2819;
											assign node2819 = (inp[2]) ? node2823 : node2820;
												assign node2820 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2823 = (inp[12]) ? node2827 : node2824;
													assign node2824 = (inp[6]) ? 8'b10101001 : 8'b10111001;
													assign node2827 = (inp[6]) ? 8'b10111001 : 8'b10101100;
											assign node2830 = (inp[2]) ? node2834 : node2831;
												assign node2831 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2834 = (inp[6]) ? node2838 : node2835;
													assign node2835 = (inp[12]) ? 8'b10101001 : 8'b10111000;
													assign node2838 = (inp[12]) ? 8'b10111000 : 8'b10101000;
									assign node2841 = (inp[10]) ? node2897 : node2842;
										assign node2842 = (inp[1]) ? node2870 : node2843;
											assign node2843 = (inp[3]) ? node2859 : node2844;
												assign node2844 = (inp[2]) ? node2852 : node2845;
													assign node2845 = (inp[6]) ? node2849 : node2846;
														assign node2846 = (inp[12]) ? 8'b10100000 : 8'b10010101;
														assign node2849 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node2852 = (inp[12]) ? node2856 : node2853;
														assign node2853 = (inp[6]) ? 8'b10000101 : 8'b10010101;
														assign node2856 = (inp[6]) ? 8'b10010101 : 8'b10100000;
												assign node2859 = (inp[2]) ? node2865 : node2860;
													assign node2860 = (inp[12]) ? 8'b10101001 : node2861;
														assign node2861 = (inp[6]) ? 8'b10101001 : 8'b10111000;
													assign node2865 = (inp[12]) ? 8'b10111000 : node2866;
														assign node2866 = (inp[6]) ? 8'b10101000 : 8'b10111000;
											assign node2870 = (inp[2]) ? node2884 : node2871;
												assign node2871 = (inp[6]) ? node2879 : node2872;
													assign node2872 = (inp[12]) ? node2876 : node2873;
														assign node2873 = (inp[3]) ? 8'b10010100 : 8'b10010101;
														assign node2876 = (inp[3]) ? 8'b10000101 : 8'b10100000;
													assign node2879 = (inp[3]) ? 8'b10011101 : node2880;
														assign node2880 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node2884 = (inp[3]) ? node2890 : node2885;
													assign node2885 = (inp[12]) ? 8'b10010101 : node2886;
														assign node2886 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node2890 = (inp[12]) ? node2894 : node2891;
														assign node2891 = (inp[6]) ? 8'b10000100 : 8'b10010100;
														assign node2894 = (inp[6]) ? 8'b10010100 : 8'b10000101;
										assign node2897 = (inp[1]) ? node2929 : node2898;
											assign node2898 = (inp[3]) ? node2914 : node2899;
												assign node2899 = (inp[2]) ? node2907 : node2900;
													assign node2900 = (inp[6]) ? node2904 : node2901;
														assign node2901 = (inp[12]) ? 8'b10101100 : 8'b10111001;
														assign node2904 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node2907 = (inp[6]) ? node2911 : node2908;
														assign node2908 = (inp[12]) ? 8'b10101100 : 8'b10111001;
														assign node2911 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2914 = (inp[2]) ? node2922 : node2915;
													assign node2915 = (inp[12]) ? node2919 : node2916;
														assign node2916 = (inp[6]) ? 8'b10101101 : 8'b10111100;
														assign node2919 = (inp[6]) ? 8'b11111101 : 8'b10101101;
													assign node2922 = (inp[12]) ? node2926 : node2923;
														assign node2923 = (inp[6]) ? 8'b10101100 : 8'b10111100;
														assign node2926 = (inp[6]) ? 8'b10111100 : 8'b10101101;
											assign node2929 = (inp[3]) ? node2941 : node2930;
												assign node2930 = (inp[2]) ? node2938 : node2931;
													assign node2931 = (inp[12]) ? node2935 : node2932;
														assign node2932 = (inp[6]) ? 8'b10101100 : 8'b10111001;
														assign node2935 = (inp[6]) ? 8'b10111100 : 8'b10101100;
													assign node2938 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node2941 = (inp[12]) ? node2947 : node2942;
													assign node2942 = (inp[6]) ? node2944 : 8'b10111000;
														assign node2944 = (inp[2]) ? 8'b10101000 : 8'b10101001;
													assign node2947 = (inp[6]) ? node2949 : 8'b10101001;
														assign node2949 = (inp[2]) ? 8'b10111000 : 8'b10111001;
								assign node2952 = (inp[10]) ? node3030 : node2953;
									assign node2953 = (inp[1]) ? node2991 : node2954;
										assign node2954 = (inp[4]) ? node2966 : node2955;
											assign node2955 = (inp[2]) ? node2959 : node2956;
												assign node2956 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2959 = (inp[12]) ? node2963 : node2960;
													assign node2960 = (inp[6]) ? 8'b10101000 : 8'b10111000;
													assign node2963 = (inp[3]) ? 8'b10111000 : 8'b10101001;
											assign node2966 = (inp[3]) ? node2982 : node2967;
												assign node2967 = (inp[2]) ? node2975 : node2968;
													assign node2968 = (inp[6]) ? node2972 : node2969;
														assign node2969 = (inp[12]) ? 8'b10100000 : 8'b10010101;
														assign node2972 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node2975 = (inp[6]) ? node2979 : node2976;
														assign node2976 = (inp[12]) ? 8'b10100000 : 8'b10010101;
														assign node2979 = (inp[12]) ? 8'b10010101 : 8'b10000101;
												assign node2982 = (inp[12]) ? node2988 : node2983;
													assign node2983 = (inp[6]) ? node2985 : 8'b10111000;
														assign node2985 = (inp[2]) ? 8'b10101000 : 8'b10101001;
													assign node2988 = (inp[6]) ? 8'b10111001 : 8'b10101001;
										assign node2991 = (inp[3]) ? node3011 : node2992;
											assign node2992 = (inp[2]) ? node3004 : node2993;
												assign node2993 = (inp[12]) ? node2999 : node2994;
													assign node2994 = (inp[4]) ? node2996 : 8'b10101000;
														assign node2996 = (inp[6]) ? 8'b10101000 : 8'b10010101;
													assign node2999 = (inp[4]) ? node3001 : 8'b10111000;
														assign node3001 = (inp[6]) ? 8'b10111000 : 8'b10100000;
												assign node3004 = (inp[12]) ? node3008 : node3005;
													assign node3005 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node3008 = (inp[6]) ? 8'b10010101 : 8'b10100000;
											assign node3011 = (inp[2]) ? node3023 : node3012;
												assign node3012 = (inp[6]) ? node3020 : node3013;
													assign node3013 = (inp[4]) ? node3017 : node3014;
														assign node3014 = (inp[12]) ? 8'b10011101 : 8'b10001101;
														assign node3017 = (inp[12]) ? 8'b10000101 : 8'b10010100;
													assign node3020 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node3023 = (inp[6]) ? node3027 : node3024;
													assign node3024 = (inp[12]) ? 8'b10000101 : 8'b10010100;
													assign node3027 = (inp[12]) ? 8'b10010100 : 8'b10000100;
									assign node3030 = (inp[1]) ? node3066 : node3031;
										assign node3031 = (inp[2]) ? node3047 : node3032;
											assign node3032 = (inp[4]) ? node3036 : node3033;
												assign node3033 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node3036 = (inp[3]) ? node3042 : node3037;
													assign node3037 = (inp[6]) ? node3039 : 8'b10000100;
														assign node3039 = (inp[12]) ? 8'b10011100 : 8'b10001100;
													assign node3042 = (inp[12]) ? 8'b10001101 : node3043;
														assign node3043 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node3047 = (inp[4]) ? node3055 : node3048;
												assign node3048 = (inp[6]) ? node3052 : node3049;
													assign node3049 = (inp[12]) ? 8'b10001101 : 8'b10011100;
													assign node3052 = (inp[12]) ? 8'b10011100 : 8'b10001100;
												assign node3055 = (inp[3]) ? node3061 : node3056;
													assign node3056 = (inp[12]) ? node3058 : 8'b10010001;
														assign node3058 = (inp[6]) ? 8'b10010001 : 8'b10000100;
													assign node3061 = (inp[12]) ? 8'b10011100 : node3062;
														assign node3062 = (inp[6]) ? 8'b10001100 : 8'b10011100;
										assign node3066 = (inp[2]) ? node3088 : node3067;
											assign node3067 = (inp[3]) ? node3077 : node3068;
												assign node3068 = (inp[6]) ? node3074 : node3069;
													assign node3069 = (inp[12]) ? node3071 : 8'b10010001;
														assign node3071 = (inp[4]) ? 8'b10000100 : 8'b10011100;
													assign node3074 = (inp[12]) ? 8'b10011100 : 8'b10001100;
												assign node3077 = (inp[12]) ? node3083 : node3078;
													assign node3078 = (inp[4]) ? node3080 : 8'b10001001;
														assign node3080 = (inp[6]) ? 8'b10001001 : 8'b10010000;
													assign node3083 = (inp[6]) ? 8'b10011001 : node3084;
														assign node3084 = (inp[4]) ? 8'b10000001 : 8'b10011001;
											assign node3088 = (inp[3]) ? node3096 : node3089;
												assign node3089 = (inp[12]) ? node3093 : node3090;
													assign node3090 = (inp[6]) ? 8'b10000001 : 8'b10010001;
													assign node3093 = (inp[6]) ? 8'b10010001 : 8'b10000100;
												assign node3096 = (inp[12]) ? node3100 : node3097;
													assign node3097 = (inp[6]) ? 8'b10000000 : 8'b10010000;
													assign node3100 = (inp[6]) ? 8'b10010000 : 8'b10000001;
				assign node3103 = (inp[11]) ? node3589 : node3104;
					assign node3104 = (inp[5]) ? node3500 : node3105;
						assign node3105 = (inp[9]) ? node3299 : node3106;
							assign node3106 = (inp[4]) ? node3160 : node3107;
								assign node3107 = (inp[1]) ? node3125 : node3108;
									assign node3108 = (inp[8]) ? node3114 : node3109;
										assign node3109 = (inp[6]) ? node3111 : 8'b11111101;
											assign node3111 = (inp[2]) ? 8'b10101101 : 8'b11111101;
										assign node3114 = (inp[10]) ? node3120 : node3115;
											assign node3115 = (inp[6]) ? node3117 : 8'b11111101;
												assign node3117 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node3120 = (inp[2]) ? node3122 : 8'b10111001;
												assign node3122 = (inp[6]) ? 8'b10101001 : 8'b10111001;
									assign node3125 = (inp[3]) ? node3143 : node3126;
										assign node3126 = (inp[2]) ? node3132 : node3127;
											assign node3127 = (inp[8]) ? node3129 : 8'b11111101;
												assign node3129 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node3132 = (inp[6]) ? node3138 : node3133;
												assign node3133 = (inp[8]) ? node3135 : 8'b11111101;
													assign node3135 = (inp[10]) ? 8'b10110001 : 8'b11110101;
												assign node3138 = (inp[8]) ? node3140 : 8'b10101101;
													assign node3140 = (inp[10]) ? 8'b10100001 : 8'b10100101;
										assign node3143 = (inp[2]) ? node3149 : node3144;
											assign node3144 = (inp[10]) ? node3146 : 8'b10111100;
												assign node3146 = (inp[8]) ? 8'b10111000 : 8'b10111100;
											assign node3149 = (inp[8]) ? node3153 : node3150;
												assign node3150 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node3153 = (inp[10]) ? node3157 : node3154;
													assign node3154 = (inp[6]) ? 8'b10100100 : 8'b10110100;
													assign node3157 = (inp[6]) ? 8'b10100000 : 8'b10110000;
								assign node3160 = (inp[3]) ? node3230 : node3161;
									assign node3161 = (inp[1]) ? node3191 : node3162;
										assign node3162 = (inp[6]) ? node3178 : node3163;
											assign node3163 = (inp[2]) ? node3171 : node3164;
												assign node3164 = (inp[8]) ? node3168 : node3165;
													assign node3165 = (inp[10]) ? 8'b10101100 : 8'b10100000;
													assign node3168 = (inp[10]) ? 8'b10100000 : 8'b10100100;
												assign node3171 = (inp[10]) ? node3175 : node3172;
													assign node3172 = (inp[8]) ? 8'b10110100 : 8'b10110000;
													assign node3175 = (inp[8]) ? 8'b10110000 : 8'b10111100;
											assign node3178 = (inp[2]) ? node3184 : node3179;
												assign node3179 = (inp[10]) ? 8'b10111000 : node3180;
													assign node3180 = (inp[8]) ? 8'b10111100 : 8'b10111000;
												assign node3184 = (inp[10]) ? node3188 : node3185;
													assign node3185 = (inp[8]) ? 8'b10100100 : 8'b10100000;
													assign node3188 = (inp[8]) ? 8'b10100000 : 8'b10101100;
										assign node3191 = (inp[8]) ? node3215 : node3192;
											assign node3192 = (inp[10]) ? node3200 : node3193;
												assign node3193 = (inp[2]) ? node3197 : node3194;
													assign node3194 = (inp[6]) ? 8'b10111001 : 8'b10100001;
													assign node3197 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node3200 = (inp[12]) ? node3208 : node3201;
													assign node3201 = (inp[2]) ? node3205 : node3202;
														assign node3202 = (inp[6]) ? 8'b11111101 : 8'b10101101;
														assign node3205 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node3208 = (inp[2]) ? node3212 : node3209;
														assign node3209 = (inp[6]) ? 8'b11111101 : 8'b10101101;
														assign node3212 = (inp[6]) ? 8'b10101101 : 8'b11111101;
											assign node3215 = (inp[10]) ? node3223 : node3216;
												assign node3216 = (inp[6]) ? node3220 : node3217;
													assign node3217 = (inp[2]) ? 8'b11110101 : 8'b10100101;
													assign node3220 = (inp[2]) ? 8'b10100101 : 8'b11111101;
												assign node3223 = (inp[2]) ? node3227 : node3224;
													assign node3224 = (inp[6]) ? 8'b10111001 : 8'b10100001;
													assign node3227 = (inp[6]) ? 8'b10100001 : 8'b10110001;
									assign node3230 = (inp[1]) ? node3268 : node3231;
										assign node3231 = (inp[8]) ? node3245 : node3232;
											assign node3232 = (inp[10]) ? node3238 : node3233;
												assign node3233 = (inp[2]) ? 8'b10111001 : node3234;
													assign node3234 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node3238 = (inp[2]) ? node3242 : node3239;
													assign node3239 = (inp[6]) ? 8'b11111101 : 8'b10101101;
													assign node3242 = (inp[6]) ? 8'b10101101 : 8'b11111101;
											assign node3245 = (inp[10]) ? node3261 : node3246;
												assign node3246 = (inp[12]) ? node3254 : node3247;
													assign node3247 = (inp[2]) ? node3251 : node3248;
														assign node3248 = (inp[6]) ? 8'b11111101 : 8'b10101101;
														assign node3251 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node3254 = (inp[2]) ? node3258 : node3255;
														assign node3255 = (inp[6]) ? 8'b11111101 : 8'b10101101;
														assign node3258 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node3261 = (inp[2]) ? node3265 : node3262;
													assign node3262 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node3265 = (inp[6]) ? 8'b10101001 : 8'b10111001;
										assign node3268 = (inp[10]) ? node3284 : node3269;
											assign node3269 = (inp[8]) ? node3277 : node3270;
												assign node3270 = (inp[2]) ? node3274 : node3271;
													assign node3271 = (inp[6]) ? 8'b10111000 : 8'b10100000;
													assign node3274 = (inp[6]) ? 8'b10100000 : 8'b10110000;
												assign node3277 = (inp[2]) ? node3281 : node3278;
													assign node3278 = (inp[6]) ? 8'b10111100 : 8'b10100100;
													assign node3281 = (inp[6]) ? 8'b10100100 : 8'b10110100;
											assign node3284 = (inp[8]) ? node3292 : node3285;
												assign node3285 = (inp[6]) ? node3289 : node3286;
													assign node3286 = (inp[2]) ? 8'b10111100 : 8'b10101100;
													assign node3289 = (inp[2]) ? 8'b10101100 : 8'b10111100;
												assign node3292 = (inp[6]) ? node3296 : node3293;
													assign node3293 = (inp[2]) ? 8'b10110000 : 8'b10100000;
													assign node3296 = (inp[2]) ? 8'b10100000 : 8'b10111000;
							assign node3299 = (inp[8]) ? node3401 : node3300;
								assign node3300 = (inp[4]) ? node3318 : node3301;
									assign node3301 = (inp[2]) ? node3307 : node3302;
										assign node3302 = (inp[1]) ? node3304 : 8'b00011111;
											assign node3304 = (inp[3]) ? 8'b00011110 : 8'b00011111;
										assign node3307 = (inp[6]) ? node3313 : node3308;
											assign node3308 = (inp[3]) ? node3310 : 8'b00011111;
												assign node3310 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node3313 = (inp[3]) ? node3315 : 8'b00001111;
												assign node3315 = (inp[1]) ? 8'b00001110 : 8'b00001111;
									assign node3318 = (inp[10]) ? node3356 : node3319;
										assign node3319 = (inp[1]) ? node3339 : node3320;
											assign node3320 = (inp[3]) ? node3332 : node3321;
												assign node3321 = (inp[12]) ? node3327 : node3322;
													assign node3322 = (inp[2]) ? node3324 : 8'b10000010;
														assign node3324 = (inp[6]) ? 8'b10000010 : 8'b10010000;
													assign node3327 = (inp[2]) ? 8'b00000010 : node3328;
														assign node3328 = (inp[6]) ? 8'b00011010 : 8'b00000010;
												assign node3332 = (inp[6]) ? node3336 : node3333;
													assign node3333 = (inp[2]) ? 8'b00011011 : 8'b00001011;
													assign node3336 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node3339 = (inp[3]) ? node3347 : node3340;
												assign node3340 = (inp[2]) ? node3344 : node3341;
													assign node3341 = (inp[6]) ? 8'b10011001 : 8'b10000001;
													assign node3344 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node3347 = (inp[2]) ? node3353 : node3348;
													assign node3348 = (inp[6]) ? 8'b00011010 : node3349;
														assign node3349 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node3353 = (inp[6]) ? 8'b10000010 : 8'b10010000;
										assign node3356 = (inp[2]) ? node3386 : node3357;
											assign node3357 = (inp[6]) ? node3371 : node3358;
												assign node3358 = (inp[12]) ? node3364 : node3359;
													assign node3359 = (inp[1]) ? node3361 : 8'b00001111;
														assign node3361 = (inp[3]) ? 8'b00001110 : 8'b00001111;
													assign node3364 = (inp[3]) ? node3368 : node3365;
														assign node3365 = (inp[1]) ? 8'b00001111 : 8'b00001110;
														assign node3368 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node3371 = (inp[12]) ? node3379 : node3372;
													assign node3372 = (inp[3]) ? node3376 : node3373;
														assign node3373 = (inp[1]) ? 8'b00011111 : 8'b00011110;
														assign node3376 = (inp[1]) ? 8'b00011110 : 8'b00011111;
													assign node3379 = (inp[3]) ? node3383 : node3380;
														assign node3380 = (inp[1]) ? 8'b00011111 : 8'b00011110;
														assign node3383 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node3386 = (inp[6]) ? node3394 : node3387;
												assign node3387 = (inp[3]) ? node3391 : node3388;
													assign node3388 = (inp[1]) ? 8'b00011111 : 8'b00011110;
													assign node3391 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node3394 = (inp[3]) ? node3398 : node3395;
													assign node3395 = (inp[1]) ? 8'b00001111 : 8'b00001110;
													assign node3398 = (inp[1]) ? 8'b00001110 : 8'b00001111;
								assign node3401 = (inp[10]) ? node3443 : node3402;
									assign node3402 = (inp[2]) ? node3424 : node3403;
										assign node3403 = (inp[4]) ? node3409 : node3404;
											assign node3404 = (inp[1]) ? node3406 : 8'b10011101;
												assign node3406 = (inp[3]) ? 8'b10011100 : 8'b10011101;
											assign node3409 = (inp[6]) ? node3417 : node3410;
												assign node3410 = (inp[3]) ? node3414 : node3411;
													assign node3411 = (inp[1]) ? 8'b10000101 : 8'b10000100;
													assign node3414 = (inp[1]) ? 8'b10000100 : 8'b10001101;
												assign node3417 = (inp[3]) ? node3421 : node3418;
													assign node3418 = (inp[1]) ? 8'b10011101 : 8'b10011100;
													assign node3421 = (inp[1]) ? 8'b10011100 : 8'b10011101;
										assign node3424 = (inp[6]) ? node3434 : node3425;
											assign node3425 = (inp[1]) ? node3431 : node3426;
												assign node3426 = (inp[3]) ? 8'b10011101 : node3427;
													assign node3427 = (inp[4]) ? 8'b10010100 : 8'b10011101;
												assign node3431 = (inp[3]) ? 8'b10010100 : 8'b10010101;
											assign node3434 = (inp[1]) ? node3440 : node3435;
												assign node3435 = (inp[3]) ? 8'b10001101 : node3436;
													assign node3436 = (inp[4]) ? 8'b10000100 : 8'b10001101;
												assign node3440 = (inp[3]) ? 8'b10000100 : 8'b10000101;
									assign node3443 = (inp[1]) ? node3477 : node3444;
										assign node3444 = (inp[4]) ? node3450 : node3445;
											assign node3445 = (inp[2]) ? node3447 : 8'b00011011;
												assign node3447 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node3450 = (inp[3]) ? node3462 : node3451;
												assign node3451 = (inp[2]) ? node3457 : node3452;
													assign node3452 = (inp[6]) ? 8'b00011010 : node3453;
														assign node3453 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node3457 = (inp[6]) ? node3459 : 8'b10010000;
														assign node3459 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3462 = (inp[12]) ? node3470 : node3463;
													assign node3463 = (inp[6]) ? node3467 : node3464;
														assign node3464 = (inp[2]) ? 8'b00011011 : 8'b00001011;
														assign node3467 = (inp[2]) ? 8'b00001011 : 8'b00011011;
													assign node3470 = (inp[2]) ? node3474 : node3471;
														assign node3471 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node3474 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node3477 = (inp[3]) ? node3487 : node3478;
											assign node3478 = (inp[2]) ? node3484 : node3479;
												assign node3479 = (inp[6]) ? 8'b10011001 : node3480;
													assign node3480 = (inp[4]) ? 8'b10000001 : 8'b10011001;
												assign node3484 = (inp[6]) ? 8'b10000001 : 8'b10010001;
											assign node3487 = (inp[2]) ? node3495 : node3488;
												assign node3488 = (inp[6]) ? 8'b00011010 : node3489;
													assign node3489 = (inp[4]) ? node3491 : 8'b00011010;
														assign node3491 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3495 = (inp[6]) ? node3497 : 8'b10010000;
													assign node3497 = (inp[12]) ? 8'b00000010 : 8'b10000010;
						assign node3500 = (inp[4]) ? node3508 : node3501;
							assign node3501 = (inp[1]) ? node3503 : 8'b11111101;
								assign node3503 = (inp[8]) ? node3505 : 8'b11111101;
									assign node3505 = (inp[2]) ? 8'b11110101 : 8'b11111101;
							assign node3508 = (inp[3]) ? node3554 : node3509;
								assign node3509 = (inp[1]) ? node3529 : node3510;
									assign node3510 = (inp[2]) ? node3524 : node3511;
										assign node3511 = (inp[6]) ? node3519 : node3512;
											assign node3512 = (inp[10]) ? node3516 : node3513;
												assign node3513 = (inp[8]) ? 8'b10100100 : 8'b10100000;
												assign node3516 = (inp[8]) ? 8'b10100100 : 8'b10101100;
											assign node3519 = (inp[10]) ? 8'b10111100 : node3520;
												assign node3520 = (inp[8]) ? 8'b10111100 : 8'b10111000;
										assign node3524 = (inp[8]) ? 8'b10110100 : node3525;
											assign node3525 = (inp[10]) ? 8'b10111100 : 8'b10110000;
									assign node3529 = (inp[6]) ? node3543 : node3530;
										assign node3530 = (inp[2]) ? node3536 : node3531;
											assign node3531 = (inp[8]) ? 8'b10100101 : node3532;
												assign node3532 = (inp[10]) ? 8'b10101101 : 8'b10100001;
											assign node3536 = (inp[10]) ? node3540 : node3537;
												assign node3537 = (inp[8]) ? 8'b11110101 : 8'b10110001;
												assign node3540 = (inp[8]) ? 8'b11110101 : 8'b11111101;
										assign node3543 = (inp[2]) ? node3549 : node3544;
											assign node3544 = (inp[8]) ? 8'b11111101 : node3545;
												assign node3545 = (inp[10]) ? 8'b11111101 : 8'b10111001;
											assign node3549 = (inp[8]) ? 8'b11110101 : node3550;
												assign node3550 = (inp[10]) ? 8'b11111101 : 8'b10110001;
								assign node3554 = (inp[6]) ? node3576 : node3555;
									assign node3555 = (inp[2]) ? node3567 : node3556;
										assign node3556 = (inp[1]) ? node3562 : node3557;
											assign node3557 = (inp[8]) ? 8'b10101101 : node3558;
												assign node3558 = (inp[10]) ? 8'b10101101 : 8'b10101001;
											assign node3562 = (inp[8]) ? 8'b10100101 : node3563;
												assign node3563 = (inp[10]) ? 8'b10101101 : 8'b10100001;
										assign node3567 = (inp[8]) ? node3573 : node3568;
											assign node3568 = (inp[10]) ? 8'b11111101 : node3569;
												assign node3569 = (inp[1]) ? 8'b10110001 : 8'b10111001;
											assign node3573 = (inp[1]) ? 8'b11110101 : 8'b11111101;
									assign node3576 = (inp[8]) ? node3584 : node3577;
										assign node3577 = (inp[10]) ? 8'b11111101 : node3578;
											assign node3578 = (inp[2]) ? node3580 : 8'b10111001;
												assign node3580 = (inp[1]) ? 8'b10110001 : 8'b10111001;
										assign node3584 = (inp[2]) ? node3586 : 8'b11111101;
											assign node3586 = (inp[1]) ? 8'b11110101 : 8'b11111101;
					assign node3589 = (inp[8]) ? node3983 : node3590;
						assign node3590 = (inp[5]) ? node3890 : node3591;
							assign node3591 = (inp[9]) ? node3739 : node3592;
								assign node3592 = (inp[4]) ? node3628 : node3593;
									assign node3593 = (inp[1]) ? node3605 : node3594;
										assign node3594 = (inp[2]) ? node3598 : node3595;
											assign node3595 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node3598 = (inp[12]) ? node3602 : node3599;
												assign node3599 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node3602 = (inp[6]) ? 8'b10101101 : 8'b10111100;
										assign node3605 = (inp[3]) ? node3617 : node3606;
											assign node3606 = (inp[2]) ? node3610 : node3607;
												assign node3607 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node3610 = (inp[6]) ? node3614 : node3611;
													assign node3611 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node3614 = (inp[12]) ? 8'b10101001 : 8'b10111000;
											assign node3617 = (inp[2]) ? node3621 : node3618;
												assign node3618 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node3621 = (inp[12]) ? node3625 : node3622;
													assign node3622 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node3625 = (inp[6]) ? 8'b10101100 : 8'b10111001;
									assign node3628 = (inp[10]) ? node3686 : node3629;
										assign node3629 = (inp[1]) ? node3659 : node3630;
											assign node3630 = (inp[3]) ? node3646 : node3631;
												assign node3631 = (inp[2]) ? node3639 : node3632;
													assign node3632 = (inp[6]) ? node3636 : node3633;
														assign node3633 = (inp[12]) ? 8'b10100000 : 8'b10010101;
														assign node3636 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node3639 = (inp[12]) ? node3643 : node3640;
														assign node3640 = (inp[6]) ? 8'b10010101 : 8'b10000101;
														assign node3643 = (inp[6]) ? 8'b10100000 : 8'b10010101;
												assign node3646 = (inp[12]) ? node3652 : node3647;
													assign node3647 = (inp[6]) ? 8'b10111000 : node3648;
														assign node3648 = (inp[2]) ? 8'b10101000 : 8'b10111000;
													assign node3652 = (inp[2]) ? node3656 : node3653;
														assign node3653 = (inp[6]) ? 8'b10111001 : 8'b10101001;
														assign node3656 = (inp[6]) ? 8'b10101001 : 8'b10111000;
											assign node3659 = (inp[3]) ? node3675 : node3660;
												assign node3660 = (inp[6]) ? node3668 : node3661;
													assign node3661 = (inp[12]) ? node3665 : node3662;
														assign node3662 = (inp[2]) ? 8'b10000100 : 8'b10010100;
														assign node3665 = (inp[2]) ? 8'b10010100 : 8'b10000101;
													assign node3668 = (inp[2]) ? node3672 : node3669;
														assign node3669 = (inp[12]) ? 8'b10011101 : 8'b10001101;
														assign node3672 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node3675 = (inp[12]) ? node3681 : node3676;
													assign node3676 = (inp[6]) ? 8'b10010101 : node3677;
														assign node3677 = (inp[2]) ? 8'b10000101 : 8'b10010101;
													assign node3681 = (inp[2]) ? node3683 : 8'b10100000;
														assign node3683 = (inp[6]) ? 8'b10100000 : 8'b10010101;
										assign node3686 = (inp[1]) ? node3712 : node3687;
											assign node3687 = (inp[3]) ? node3701 : node3688;
												assign node3688 = (inp[12]) ? node3694 : node3689;
													assign node3689 = (inp[2]) ? node3691 : 8'b10111001;
														assign node3691 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node3694 = (inp[2]) ? node3698 : node3695;
														assign node3695 = (inp[6]) ? 8'b10111100 : 8'b10101100;
														assign node3698 = (inp[6]) ? 8'b10101100 : 8'b10111001;
												assign node3701 = (inp[6]) ? node3707 : node3702;
													assign node3702 = (inp[2]) ? node3704 : 8'b10111100;
														assign node3704 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node3707 = (inp[12]) ? node3709 : 8'b10101101;
														assign node3709 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node3712 = (inp[3]) ? node3726 : node3713;
												assign node3713 = (inp[2]) ? node3721 : node3714;
													assign node3714 = (inp[12]) ? node3718 : node3715;
														assign node3715 = (inp[6]) ? 8'b10101001 : 8'b10111000;
														assign node3718 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node3721 = (inp[6]) ? 8'b10111000 : node3722;
														assign node3722 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node3726 = (inp[2]) ? node3734 : node3727;
													assign node3727 = (inp[6]) ? node3731 : node3728;
														assign node3728 = (inp[12]) ? 8'b10101100 : 8'b10111001;
														assign node3731 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node3734 = (inp[12]) ? 8'b10111001 : node3735;
														assign node3735 = (inp[6]) ? 8'b10111001 : 8'b10101001;
								assign node3739 = (inp[4]) ? node3775 : node3740;
									assign node3740 = (inp[1]) ? node3752 : node3741;
										assign node3741 = (inp[2]) ? node3745 : node3742;
											assign node3742 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node3745 = (inp[6]) ? node3749 : node3746;
												assign node3746 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node3749 = (inp[12]) ? 8'b00001111 : 8'b00011110;
										assign node3752 = (inp[3]) ? node3764 : node3753;
											assign node3753 = (inp[2]) ? node3757 : node3754;
												assign node3754 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node3757 = (inp[6]) ? node3761 : node3758;
													assign node3758 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3761 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node3764 = (inp[2]) ? node3768 : node3765;
												assign node3765 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node3768 = (inp[12]) ? node3772 : node3769;
													assign node3769 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node3772 = (inp[6]) ? 8'b00001110 : 8'b00011011;
									assign node3775 = (inp[10]) ? node3833 : node3776;
										assign node3776 = (inp[3]) ? node3804 : node3777;
											assign node3777 = (inp[1]) ? node3789 : node3778;
												assign node3778 = (inp[2]) ? node3782 : node3779;
													assign node3779 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node3782 = (inp[6]) ? node3786 : node3783;
														assign node3783 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node3786 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node3789 = (inp[2]) ? node3797 : node3790;
													assign node3790 = (inp[6]) ? node3794 : node3791;
														assign node3791 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node3794 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node3797 = (inp[12]) ? node3801 : node3798;
														assign node3798 = (inp[6]) ? 8'b10110100 : 8'b10100100;
														assign node3801 = (inp[6]) ? 8'b10100101 : 8'b10110100;
											assign node3804 = (inp[1]) ? node3820 : node3805;
												assign node3805 = (inp[12]) ? node3813 : node3806;
													assign node3806 = (inp[6]) ? node3810 : node3807;
														assign node3807 = (inp[2]) ? 8'b00001010 : 8'b00011010;
														assign node3810 = (inp[2]) ? 8'b00011010 : 8'b00001011;
													assign node3813 = (inp[2]) ? node3817 : node3814;
														assign node3814 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node3817 = (inp[6]) ? 8'b00001011 : 8'b00011010;
												assign node3820 = (inp[2]) ? node3826 : node3821;
													assign node3821 = (inp[6]) ? node3823 : 8'b00000010;
														assign node3823 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3826 = (inp[6]) ? node3830 : node3827;
														assign node3827 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node3830 = (inp[12]) ? 8'b00000010 : 8'b11110111;
										assign node3833 = (inp[1]) ? node3859 : node3834;
											assign node3834 = (inp[3]) ? node3850 : node3835;
												assign node3835 = (inp[2]) ? node3843 : node3836;
													assign node3836 = (inp[12]) ? node3840 : node3837;
														assign node3837 = (inp[6]) ? 8'b00001110 : 8'b00011011;
														assign node3840 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node3843 = (inp[6]) ? node3847 : node3844;
														assign node3844 = (inp[12]) ? 8'b00011011 : 8'b00001011;
														assign node3847 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node3850 = (inp[2]) ? node3852 : 8'b00001111;
													assign node3852 = (inp[12]) ? node3856 : node3853;
														assign node3853 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node3856 = (inp[6]) ? 8'b00001111 : 8'b00011110;
											assign node3859 = (inp[3]) ? node3875 : node3860;
												assign node3860 = (inp[12]) ? node3868 : node3861;
													assign node3861 = (inp[2]) ? node3865 : node3862;
														assign node3862 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node3865 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node3868 = (inp[6]) ? node3872 : node3869;
														assign node3869 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node3872 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node3875 = (inp[2]) ? node3883 : node3876;
													assign node3876 = (inp[6]) ? node3880 : node3877;
														assign node3877 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node3880 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node3883 = (inp[12]) ? node3887 : node3884;
														assign node3884 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node3887 = (inp[6]) ? 8'b00001110 : 8'b00011011;
							assign node3890 = (inp[12]) ? node3936 : node3891;
								assign node3891 = (inp[2]) ? node3921 : node3892;
									assign node3892 = (inp[4]) ? node3896 : node3893;
										assign node3893 = (inp[1]) ? 8'b10101001 : 8'b10101101;
										assign node3896 = (inp[6]) ? node3910 : node3897;
											assign node3897 = (inp[10]) ? node3903 : node3898;
												assign node3898 = (inp[1]) ? 8'b10010100 : node3899;
													assign node3899 = (inp[3]) ? 8'b10111000 : 8'b10010101;
												assign node3903 = (inp[3]) ? node3907 : node3904;
													assign node3904 = (inp[1]) ? 8'b10111000 : 8'b10111001;
													assign node3907 = (inp[1]) ? 8'b10111000 : 8'b10111100;
											assign node3910 = (inp[1]) ? node3918 : node3911;
												assign node3911 = (inp[3]) ? node3915 : node3912;
													assign node3912 = (inp[10]) ? 8'b10101100 : 8'b10101000;
													assign node3915 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node3918 = (inp[10]) ? 8'b10101001 : 8'b10001101;
									assign node3921 = (inp[1]) ? node3931 : node3922;
										assign node3922 = (inp[4]) ? node3924 : 8'b10101100;
											assign node3924 = (inp[3]) ? node3928 : node3925;
												assign node3925 = (inp[10]) ? 8'b10101001 : 8'b10000101;
												assign node3928 = (inp[10]) ? 8'b10101100 : 8'b10101000;
										assign node3931 = (inp[4]) ? node3933 : 8'b10101000;
											assign node3933 = (inp[10]) ? 8'b10101000 : 8'b10000100;
								assign node3936 = (inp[2]) ? node3964 : node3937;
									assign node3937 = (inp[1]) ? node3955 : node3938;
										assign node3938 = (inp[4]) ? node3940 : 8'b11111101;
											assign node3940 = (inp[10]) ? node3948 : node3941;
												assign node3941 = (inp[6]) ? node3945 : node3942;
													assign node3942 = (inp[3]) ? 8'b10101001 : 8'b10100000;
													assign node3945 = (inp[3]) ? 8'b10111001 : 8'b10111000;
												assign node3948 = (inp[3]) ? node3952 : node3949;
													assign node3949 = (inp[6]) ? 8'b10111100 : 8'b10101100;
													assign node3952 = (inp[6]) ? 8'b11111101 : 8'b10101101;
										assign node3955 = (inp[4]) ? node3957 : 8'b10111001;
											assign node3957 = (inp[10]) ? node3961 : node3958;
												assign node3958 = (inp[6]) ? 8'b10011101 : 8'b10000101;
												assign node3961 = (inp[6]) ? 8'b10111001 : 8'b10101001;
									assign node3964 = (inp[4]) ? node3968 : node3965;
										assign node3965 = (inp[1]) ? 8'b10111000 : 8'b10111100;
										assign node3968 = (inp[10]) ? node3976 : node3969;
											assign node3969 = (inp[3]) ? node3973 : node3970;
												assign node3970 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node3973 = (inp[1]) ? 8'b10010100 : 8'b10111000;
											assign node3976 = (inp[3]) ? node3980 : node3977;
												assign node3977 = (inp[1]) ? 8'b10111000 : 8'b10111001;
												assign node3980 = (inp[1]) ? 8'b10111000 : 8'b10111100;
						assign node3983 = (inp[1]) ? node4165 : node3984;
							assign node3984 = (inp[5]) ? node4134 : node3985;
								assign node3985 = (inp[10]) ? node4059 : node3986;
									assign node3986 = (inp[9]) ? node4022 : node3987;
										assign node3987 = (inp[4]) ? node3999 : node3988;
											assign node3988 = (inp[2]) ? node3992 : node3989;
												assign node3989 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node3992 = (inp[6]) ? node3996 : node3993;
													assign node3993 = (inp[12]) ? 8'b10011100 : 8'b10001100;
													assign node3996 = (inp[12]) ? 8'b10001101 : 8'b10011100;
											assign node3999 = (inp[3]) ? node4011 : node4000;
												assign node4000 = (inp[6]) ? node4008 : node4001;
													assign node4001 = (inp[12]) ? node4005 : node4002;
														assign node4002 = (inp[2]) ? 8'b10000001 : 8'b10010001;
														assign node4005 = (inp[2]) ? 8'b10010001 : 8'b10000100;
													assign node4008 = (inp[12]) ? 8'b10000100 : 8'b10001100;
												assign node4011 = (inp[12]) ? node4017 : node4012;
													assign node4012 = (inp[6]) ? 8'b10001101 : node4013;
														assign node4013 = (inp[2]) ? 8'b10001100 : 8'b10011100;
													assign node4017 = (inp[2]) ? 8'b10001101 : node4018;
														assign node4018 = (inp[6]) ? 8'b10011101 : 8'b10001101;
										assign node4022 = (inp[2]) ? node4040 : node4023;
											assign node4023 = (inp[12]) ? node4031 : node4024;
												assign node4024 = (inp[4]) ? node4026 : 8'b10101101;
													assign node4026 = (inp[6]) ? node4028 : 8'b10110001;
														assign node4028 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node4031 = (inp[4]) ? node4033 : 8'b11111101;
													assign node4033 = (inp[6]) ? node4037 : node4034;
														assign node4034 = (inp[3]) ? 8'b10101101 : 8'b10100100;
														assign node4037 = (inp[3]) ? 8'b11111101 : 8'b10111100;
											assign node4040 = (inp[3]) ? node4052 : node4041;
												assign node4041 = (inp[4]) ? node4047 : node4042;
													assign node4042 = (inp[6]) ? 8'b10101101 : node4043;
														assign node4043 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node4047 = (inp[6]) ? node4049 : 8'b10110001;
														assign node4049 = (inp[12]) ? 8'b10100100 : 8'b10110001;
												assign node4052 = (inp[12]) ? node4056 : node4053;
													assign node4053 = (inp[6]) ? 8'b10111100 : 8'b10101100;
													assign node4056 = (inp[6]) ? 8'b10101101 : 8'b10111100;
									assign node4059 = (inp[9]) ? node4099 : node4060;
										assign node4060 = (inp[4]) ? node4072 : node4061;
											assign node4061 = (inp[2]) ? node4065 : node4062;
												assign node4062 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node4065 = (inp[6]) ? node4069 : node4066;
													assign node4066 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node4069 = (inp[12]) ? 8'b10101001 : 8'b10111000;
											assign node4072 = (inp[3]) ? node4086 : node4073;
												assign node4073 = (inp[12]) ? node4081 : node4074;
													assign node4074 = (inp[6]) ? node4078 : node4075;
														assign node4075 = (inp[2]) ? 8'b10000101 : 8'b10010101;
														assign node4078 = (inp[2]) ? 8'b10010101 : 8'b10101000;
													assign node4081 = (inp[2]) ? 8'b10100000 : node4082;
														assign node4082 = (inp[6]) ? 8'b10111000 : 8'b10100000;
												assign node4086 = (inp[12]) ? node4094 : node4087;
													assign node4087 = (inp[6]) ? node4091 : node4088;
														assign node4088 = (inp[2]) ? 8'b10101000 : 8'b10111000;
														assign node4091 = (inp[2]) ? 8'b10111000 : 8'b10101001;
													assign node4094 = (inp[6]) ? node4096 : 8'b10101001;
														assign node4096 = (inp[2]) ? 8'b10101001 : 8'b10111001;
										assign node4099 = (inp[4]) ? node4111 : node4100;
											assign node4100 = (inp[2]) ? node4104 : node4101;
												assign node4101 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node4104 = (inp[12]) ? node4108 : node4105;
													assign node4105 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node4108 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node4111 = (inp[3]) ? node4127 : node4112;
												assign node4112 = (inp[2]) ? node4120 : node4113;
													assign node4113 = (inp[6]) ? node4117 : node4114;
														assign node4114 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node4117 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node4120 = (inp[6]) ? node4124 : node4121;
														assign node4121 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node4124 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node4127 = (inp[6]) ? node4129 : 8'b00011010;
													assign node4129 = (inp[2]) ? 8'b00001011 : node4130;
														assign node4130 = (inp[12]) ? 8'b00011011 : 8'b00001011;
								assign node4134 = (inp[12]) ? node4150 : node4135;
									assign node4135 = (inp[2]) ? node4145 : node4136;
										assign node4136 = (inp[4]) ? node4138 : 8'b10001101;
											assign node4138 = (inp[6]) ? node4142 : node4139;
												assign node4139 = (inp[3]) ? 8'b10011100 : 8'b10010001;
												assign node4142 = (inp[3]) ? 8'b10001101 : 8'b10001100;
										assign node4145 = (inp[3]) ? 8'b10001100 : node4146;
											assign node4146 = (inp[4]) ? 8'b10000001 : 8'b10001100;
									assign node4150 = (inp[2]) ? node4160 : node4151;
										assign node4151 = (inp[4]) ? node4153 : 8'b10011101;
											assign node4153 = (inp[6]) ? node4157 : node4154;
												assign node4154 = (inp[3]) ? 8'b10001101 : 8'b10000100;
												assign node4157 = (inp[3]) ? 8'b10011101 : 8'b10011100;
										assign node4160 = (inp[3]) ? 8'b10011100 : node4161;
											assign node4161 = (inp[4]) ? 8'b10010001 : 8'b10011100;
							assign node4165 = (inp[2]) ? node4255 : node4166;
								assign node4166 = (inp[5]) ? node4244 : node4167;
									assign node4167 = (inp[3]) ? node4209 : node4168;
										assign node4168 = (inp[10]) ? node4188 : node4169;
											assign node4169 = (inp[9]) ? node4177 : node4170;
												assign node4170 = (inp[12]) ? 8'b10011001 : node4171;
													assign node4171 = (inp[6]) ? 8'b10001001 : node4172;
														assign node4172 = (inp[4]) ? 8'b10010000 : 8'b10001001;
												assign node4177 = (inp[12]) ? node4183 : node4178;
													assign node4178 = (inp[4]) ? node4180 : 8'b10101001;
														assign node4180 = (inp[6]) ? 8'b10101001 : 8'b10110000;
													assign node4183 = (inp[6]) ? 8'b10111001 : node4184;
														assign node4184 = (inp[4]) ? 8'b10100001 : 8'b10111001;
											assign node4188 = (inp[9]) ? node4200 : node4189;
												assign node4189 = (inp[6]) ? node4197 : node4190;
													assign node4190 = (inp[4]) ? node4194 : node4191;
														assign node4191 = (inp[12]) ? 8'b10011101 : 8'b10001101;
														assign node4194 = (inp[12]) ? 8'b10000101 : 8'b10010100;
													assign node4197 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node4200 = (inp[12]) ? node4204 : node4201;
													assign node4201 = (inp[6]) ? 8'b10101101 : 8'b10110100;
													assign node4204 = (inp[6]) ? 8'b11111101 : node4205;
														assign node4205 = (inp[4]) ? 8'b10100101 : 8'b11111101;
										assign node4209 = (inp[10]) ? node4227 : node4210;
											assign node4210 = (inp[9]) ? node4220 : node4211;
												assign node4211 = (inp[4]) ? node4215 : node4212;
													assign node4212 = (inp[12]) ? 8'b10011100 : 8'b10001100;
													assign node4215 = (inp[6]) ? 8'b10001100 : node4216;
														assign node4216 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node4220 = (inp[12]) ? 8'b10111100 : node4221;
													assign node4221 = (inp[4]) ? node4223 : 8'b10101100;
														assign node4223 = (inp[6]) ? 8'b10101100 : 8'b10110001;
											assign node4227 = (inp[9]) ? node4235 : node4228;
												assign node4228 = (inp[6]) ? node4232 : node4229;
													assign node4229 = (inp[12]) ? 8'b10100000 : 8'b10010101;
													assign node4232 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node4235 = (inp[6]) ? node4241 : node4236;
													assign node4236 = (inp[4]) ? node4238 : 8'b00001010;
														assign node4238 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node4241 = (inp[12]) ? 8'b00011010 : 8'b00001010;
									assign node4244 = (inp[6]) ? node4252 : node4245;
										assign node4245 = (inp[4]) ? node4249 : node4246;
											assign node4246 = (inp[12]) ? 8'b10011001 : 8'b10001001;
											assign node4249 = (inp[12]) ? 8'b10000001 : 8'b10010000;
										assign node4252 = (inp[12]) ? 8'b10011001 : 8'b10001001;
								assign node4255 = (inp[5]) ? node4319 : node4256;
									assign node4256 = (inp[9]) ? node4288 : node4257;
										assign node4257 = (inp[10]) ? node4273 : node4258;
											assign node4258 = (inp[3]) ? node4266 : node4259;
												assign node4259 = (inp[6]) ? node4263 : node4260;
													assign node4260 = (inp[12]) ? 8'b10010000 : 8'b10000000;
													assign node4263 = (inp[12]) ? 8'b10000001 : 8'b10010000;
												assign node4266 = (inp[6]) ? node4270 : node4267;
													assign node4267 = (inp[12]) ? 8'b10010001 : 8'b10000001;
													assign node4270 = (inp[12]) ? 8'b10000100 : 8'b10010001;
											assign node4273 = (inp[3]) ? node4281 : node4274;
												assign node4274 = (inp[12]) ? node4278 : node4275;
													assign node4275 = (inp[6]) ? 8'b10010100 : 8'b10000100;
													assign node4278 = (inp[6]) ? 8'b10000101 : 8'b10010100;
												assign node4281 = (inp[12]) ? node4285 : node4282;
													assign node4282 = (inp[6]) ? 8'b10010101 : 8'b10000101;
													assign node4285 = (inp[6]) ? 8'b10100000 : 8'b10010101;
										assign node4288 = (inp[10]) ? node4304 : node4289;
											assign node4289 = (inp[3]) ? node4297 : node4290;
												assign node4290 = (inp[12]) ? node4294 : node4291;
													assign node4291 = (inp[6]) ? 8'b10110000 : 8'b10100000;
													assign node4294 = (inp[6]) ? 8'b10100001 : 8'b10110000;
												assign node4297 = (inp[6]) ? node4301 : node4298;
													assign node4298 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node4301 = (inp[12]) ? 8'b10100100 : 8'b10110001;
											assign node4304 = (inp[3]) ? node4312 : node4305;
												assign node4305 = (inp[12]) ? node4309 : node4306;
													assign node4306 = (inp[6]) ? 8'b10110100 : 8'b10100100;
													assign node4309 = (inp[6]) ? 8'b10100101 : 8'b10110100;
												assign node4312 = (inp[6]) ? node4316 : node4313;
													assign node4313 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node4316 = (inp[12]) ? 8'b00000010 : 8'b11110111;
									assign node4319 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node4322 = (inp[4]) ? node7518 : node4323;
			assign node4323 = (inp[13]) ? node5989 : node4324;
				assign node4324 = (inp[9]) ? node5144 : node4325;
					assign node4325 = (inp[11]) ? node4617 : node4326;
						assign node4326 = (inp[3]) ? node4482 : node4327;
							assign node4327 = (inp[0]) ? node4459 : node4328;
								assign node4328 = (inp[1]) ? node4402 : node4329;
									assign node4329 = (inp[5]) ? node4347 : node4330;
										assign node4330 = (inp[10]) ? node4342 : node4331;
											assign node4331 = (inp[8]) ? node4337 : node4332;
												assign node4332 = (inp[2]) ? 8'b00101111 : node4333;
													assign node4333 = (inp[6]) ? 8'b00101111 : 8'b01111111;
												assign node4337 = (inp[12]) ? 8'b00101011 : node4338;
													assign node4338 = (inp[6]) ? 8'b00101011 : 8'b00111011;
											assign node4342 = (inp[2]) ? 8'b00101011 : node4343;
												assign node4343 = (inp[6]) ? 8'b00101011 : 8'b00111011;
										assign node4347 = (inp[12]) ? node4377 : node4348;
											assign node4348 = (inp[2]) ? node4362 : node4349;
												assign node4349 = (inp[6]) ? node4355 : node4350;
													assign node4350 = (inp[10]) ? node4352 : 8'b00111011;
														assign node4352 = (inp[8]) ? 8'b01111111 : 8'b00111011;
													assign node4355 = (inp[10]) ? node4359 : node4356;
														assign node4356 = (inp[8]) ? 8'b00101011 : 8'b00101111;
														assign node4359 = (inp[8]) ? 8'b00101111 : 8'b00101011;
												assign node4362 = (inp[6]) ? node4370 : node4363;
													assign node4363 = (inp[10]) ? node4367 : node4364;
														assign node4364 = (inp[8]) ? 8'b00101011 : 8'b00101111;
														assign node4367 = (inp[8]) ? 8'b00101111 : 8'b00101011;
													assign node4370 = (inp[10]) ? node4374 : node4371;
														assign node4371 = (inp[8]) ? 8'b00111011 : 8'b01111111;
														assign node4374 = (inp[8]) ? 8'b01111111 : 8'b00111011;
											assign node4377 = (inp[2]) ? node4393 : node4378;
												assign node4378 = (inp[6]) ? node4386 : node4379;
													assign node4379 = (inp[8]) ? node4383 : node4380;
														assign node4380 = (inp[10]) ? 8'b00111011 : 8'b01111111;
														assign node4383 = (inp[10]) ? 8'b01111111 : 8'b00111011;
													assign node4386 = (inp[8]) ? node4390 : node4387;
														assign node4387 = (inp[10]) ? 8'b00101011 : 8'b00101111;
														assign node4390 = (inp[10]) ? 8'b00101111 : 8'b00101011;
												assign node4393 = (inp[6]) ? 8'b00111011 : node4394;
													assign node4394 = (inp[8]) ? node4398 : node4395;
														assign node4395 = (inp[10]) ? 8'b00101011 : 8'b00101111;
														assign node4398 = (inp[10]) ? 8'b00101111 : 8'b00101011;
									assign node4402 = (inp[5]) ? node4420 : node4403;
										assign node4403 = (inp[2]) ? node4415 : node4404;
											assign node4404 = (inp[6]) ? node4410 : node4405;
												assign node4405 = (inp[10]) ? 8'b00111010 : node4406;
													assign node4406 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node4410 = (inp[8]) ? 8'b00101010 : node4411;
													assign node4411 = (inp[10]) ? 8'b00101010 : 8'b00101110;
											assign node4415 = (inp[10]) ? 8'b00101010 : node4416;
												assign node4416 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node4420 = (inp[10]) ? node4444 : node4421;
											assign node4421 = (inp[8]) ? node4429 : node4422;
												assign node4422 = (inp[2]) ? node4426 : node4423;
													assign node4423 = (inp[6]) ? 8'b00101110 : 8'b00111110;
													assign node4426 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node4429 = (inp[12]) ? node4437 : node4430;
													assign node4430 = (inp[6]) ? node4434 : node4431;
														assign node4431 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node4434 = (inp[2]) ? 8'b00111010 : 8'b00101010;
													assign node4437 = (inp[6]) ? node4441 : node4438;
														assign node4438 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node4441 = (inp[2]) ? 8'b00111010 : 8'b00101010;
											assign node4444 = (inp[8]) ? node4452 : node4445;
												assign node4445 = (inp[6]) ? node4449 : node4446;
													assign node4446 = (inp[2]) ? 8'b00101010 : 8'b00111010;
													assign node4449 = (inp[2]) ? 8'b00111010 : 8'b00101010;
												assign node4452 = (inp[6]) ? node4456 : node4453;
													assign node4453 = (inp[2]) ? 8'b00101110 : 8'b00111110;
													assign node4456 = (inp[2]) ? 8'b00111110 : 8'b00101110;
								assign node4459 = (inp[6]) ? node4467 : node4460;
									assign node4460 = (inp[10]) ? node4462 : 8'b01111111;
										assign node4462 = (inp[8]) ? node4464 : 8'b00111011;
											assign node4464 = (inp[5]) ? 8'b01111111 : 8'b00111011;
									assign node4467 = (inp[10]) ? node4473 : node4468;
										assign node4468 = (inp[2]) ? node4470 : 8'b00101111;
											assign node4470 = (inp[5]) ? 8'b01111111 : 8'b00101111;
										assign node4473 = (inp[5]) ? node4475 : 8'b00101011;
											assign node4475 = (inp[2]) ? node4479 : node4476;
												assign node4476 = (inp[8]) ? 8'b00101111 : 8'b00101011;
												assign node4479 = (inp[8]) ? 8'b01111111 : 8'b00111011;
							assign node4482 = (inp[5]) ? node4506 : node4483;
								assign node4483 = (inp[6]) ? node4499 : node4484;
									assign node4484 = (inp[10]) ? node4494 : node4485;
										assign node4485 = (inp[0]) ? 8'b00111110 : node4486;
											assign node4486 = (inp[2]) ? node4490 : node4487;
												assign node4487 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node4490 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node4494 = (inp[2]) ? node4496 : 8'b00111010;
											assign node4496 = (inp[0]) ? 8'b00111010 : 8'b00101010;
									assign node4499 = (inp[10]) ? 8'b00101010 : node4500;
										assign node4500 = (inp[8]) ? node4502 : 8'b00101110;
											assign node4502 = (inp[0]) ? 8'b00101110 : 8'b00101010;
								assign node4506 = (inp[1]) ? node4570 : node4507;
									assign node4507 = (inp[0]) ? node4553 : node4508;
										assign node4508 = (inp[10]) ? node4532 : node4509;
											assign node4509 = (inp[8]) ? node4525 : node4510;
												assign node4510 = (inp[12]) ? node4518 : node4511;
													assign node4511 = (inp[6]) ? node4515 : node4512;
														assign node4512 = (inp[2]) ? 8'b00101110 : 8'b00111110;
														assign node4515 = (inp[2]) ? 8'b00111110 : 8'b00101110;
													assign node4518 = (inp[6]) ? node4522 : node4519;
														assign node4519 = (inp[2]) ? 8'b00101110 : 8'b00111110;
														assign node4522 = (inp[2]) ? 8'b00111110 : 8'b00101110;
												assign node4525 = (inp[6]) ? node4529 : node4526;
													assign node4526 = (inp[2]) ? 8'b00101010 : 8'b00111010;
													assign node4529 = (inp[2]) ? 8'b00111010 : 8'b00101010;
											assign node4532 = (inp[8]) ? node4546 : node4533;
												assign node4533 = (inp[12]) ? node4541 : node4534;
													assign node4534 = (inp[6]) ? node4538 : node4535;
														assign node4535 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node4538 = (inp[2]) ? 8'b00111010 : 8'b00101010;
													assign node4541 = (inp[2]) ? 8'b00101010 : node4542;
														assign node4542 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node4546 = (inp[6]) ? node4550 : node4547;
													assign node4547 = (inp[2]) ? 8'b00101110 : 8'b00111110;
													assign node4550 = (inp[2]) ? 8'b00111110 : 8'b00101110;
										assign node4553 = (inp[8]) ? node4565 : node4554;
											assign node4554 = (inp[10]) ? node4560 : node4555;
												assign node4555 = (inp[6]) ? node4557 : 8'b00111110;
													assign node4557 = (inp[2]) ? 8'b00111110 : 8'b00101110;
												assign node4560 = (inp[6]) ? node4562 : 8'b00111010;
													assign node4562 = (inp[2]) ? 8'b00111010 : 8'b00101010;
											assign node4565 = (inp[2]) ? 8'b00111110 : node4566;
												assign node4566 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node4570 = (inp[0]) ? node4604 : node4571;
										assign node4571 = (inp[8]) ? node4583 : node4572;
											assign node4572 = (inp[10]) ? node4580 : node4573;
												assign node4573 = (inp[6]) ? node4577 : node4574;
													assign node4574 = (inp[2]) ? 8'b00101111 : 8'b01111111;
													assign node4577 = (inp[2]) ? 8'b01111111 : 8'b00101111;
												assign node4580 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node4583 = (inp[10]) ? node4591 : node4584;
												assign node4584 = (inp[6]) ? node4588 : node4585;
													assign node4585 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node4588 = (inp[2]) ? 8'b00111011 : 8'b00101011;
												assign node4591 = (inp[12]) ? node4597 : node4592;
													assign node4592 = (inp[6]) ? node4594 : 8'b01111111;
														assign node4594 = (inp[2]) ? 8'b01111111 : 8'b00101111;
													assign node4597 = (inp[2]) ? node4601 : node4598;
														assign node4598 = (inp[6]) ? 8'b00101111 : 8'b01111111;
														assign node4601 = (inp[6]) ? 8'b01111111 : 8'b00101111;
										assign node4604 = (inp[2]) ? node4612 : node4605;
											assign node4605 = (inp[6]) ? node4607 : 8'b01111111;
												assign node4607 = (inp[8]) ? 8'b00101111 : node4608;
													assign node4608 = (inp[10]) ? 8'b00101011 : 8'b00101111;
											assign node4612 = (inp[10]) ? node4614 : 8'b01111111;
												assign node4614 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node4617 = (inp[8]) ? node4881 : node4618;
							assign node4618 = (inp[10]) ? node4750 : node4619;
								assign node4619 = (inp[1]) ? node4675 : node4620;
									assign node4620 = (inp[3]) ? node4648 : node4621;
										assign node4621 = (inp[2]) ? node4629 : node4622;
											assign node4622 = (inp[12]) ? node4626 : node4623;
												assign node4623 = (inp[6]) ? 8'b00111110 : 8'b00101111;
												assign node4626 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node4629 = (inp[12]) ? node4641 : node4630;
												assign node4630 = (inp[5]) ? node4636 : node4631;
													assign node4631 = (inp[6]) ? 8'b00111110 : node4632;
														assign node4632 = (inp[0]) ? 8'b00101110 : 8'b00111110;
													assign node4636 = (inp[6]) ? 8'b00101110 : node4637;
														assign node4637 = (inp[0]) ? 8'b00101110 : 8'b00111110;
												assign node4641 = (inp[5]) ? node4643 : 8'b00101111;
													assign node4643 = (inp[6]) ? 8'b00111110 : node4644;
														assign node4644 = (inp[0]) ? 8'b00111110 : 8'b00101111;
										assign node4648 = (inp[12]) ? node4660 : node4649;
											assign node4649 = (inp[6]) ? node4655 : node4650;
												assign node4650 = (inp[2]) ? node4652 : 8'b00101110;
													assign node4652 = (inp[0]) ? 8'b00101011 : 8'b00111011;
												assign node4655 = (inp[5]) ? node4657 : 8'b00111011;
													assign node4657 = (inp[2]) ? 8'b00101011 : 8'b00111011;
											assign node4660 = (inp[2]) ? node4664 : node4661;
												assign node4661 = (inp[6]) ? 8'b00101110 : 8'b00111110;
												assign node4664 = (inp[5]) ? node4670 : node4665;
													assign node4665 = (inp[0]) ? node4667 : 8'b00101110;
														assign node4667 = (inp[6]) ? 8'b00101110 : 8'b00111011;
													assign node4670 = (inp[0]) ? 8'b00111011 : node4671;
														assign node4671 = (inp[6]) ? 8'b00111011 : 8'b00101110;
									assign node4675 = (inp[0]) ? node4717 : node4676;
										assign node4676 = (inp[12]) ? node4696 : node4677;
											assign node4677 = (inp[5]) ? node4683 : node4678;
												assign node4678 = (inp[2]) ? 8'b00111011 : node4679;
													assign node4679 = (inp[6]) ? 8'b00111011 : 8'b00101110;
												assign node4683 = (inp[3]) ? node4691 : node4684;
													assign node4684 = (inp[6]) ? node4688 : node4685;
														assign node4685 = (inp[2]) ? 8'b00111011 : 8'b00101110;
														assign node4688 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node4691 = (inp[2]) ? node4693 : 8'b00101011;
														assign node4693 = (inp[6]) ? 8'b00101010 : 8'b00111010;
											assign node4696 = (inp[5]) ? node4702 : node4697;
												assign node4697 = (inp[6]) ? 8'b00101110 : node4698;
													assign node4698 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node4702 = (inp[3]) ? node4710 : node4703;
													assign node4703 = (inp[2]) ? node4707 : node4704;
														assign node4704 = (inp[6]) ? 8'b00101110 : 8'b00111110;
														assign node4707 = (inp[6]) ? 8'b00111011 : 8'b00101110;
													assign node4710 = (inp[2]) ? node4714 : node4711;
														assign node4711 = (inp[6]) ? 8'b00101011 : 8'b00111011;
														assign node4714 = (inp[6]) ? 8'b00111010 : 8'b00101011;
										assign node4717 = (inp[12]) ? node4731 : node4718;
											assign node4718 = (inp[6]) ? node4728 : node4719;
												assign node4719 = (inp[2]) ? node4723 : node4720;
													assign node4720 = (inp[5]) ? 8'b00101011 : 8'b00101110;
													assign node4723 = (inp[5]) ? 8'b00101010 : node4724;
														assign node4724 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node4728 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node4731 = (inp[6]) ? node4743 : node4732;
												assign node4732 = (inp[2]) ? node4738 : node4733;
													assign node4733 = (inp[5]) ? 8'b00111011 : node4734;
														assign node4734 = (inp[3]) ? 8'b00111110 : 8'b00111011;
													assign node4738 = (inp[3]) ? node4740 : 8'b00111010;
														assign node4740 = (inp[5]) ? 8'b00111010 : 8'b00111011;
												assign node4743 = (inp[2]) ? node4745 : 8'b00101011;
													assign node4745 = (inp[5]) ? 8'b00111010 : node4746;
														assign node4746 = (inp[3]) ? 8'b00101110 : 8'b00101011;
								assign node4750 = (inp[1]) ? node4802 : node4751;
									assign node4751 = (inp[3]) ? node4775 : node4752;
										assign node4752 = (inp[12]) ? node4764 : node4753;
											assign node4753 = (inp[6]) ? node4759 : node4754;
												assign node4754 = (inp[2]) ? node4756 : 8'b00101011;
													assign node4756 = (inp[0]) ? 8'b00101010 : 8'b00111010;
												assign node4759 = (inp[2]) ? node4761 : 8'b00111010;
													assign node4761 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node4764 = (inp[6]) ? node4770 : node4765;
												assign node4765 = (inp[2]) ? node4767 : 8'b00111011;
													assign node4767 = (inp[0]) ? 8'b00111010 : 8'b00101011;
												assign node4770 = (inp[2]) ? node4772 : 8'b00101011;
													assign node4772 = (inp[5]) ? 8'b00111010 : 8'b00101011;
										assign node4775 = (inp[12]) ? node4787 : node4776;
											assign node4776 = (inp[6]) ? node4782 : node4777;
												assign node4777 = (inp[2]) ? node4779 : 8'b00101010;
													assign node4779 = (inp[0]) ? 8'b00001111 : 8'b00011111;
												assign node4782 = (inp[5]) ? node4784 : 8'b00011111;
													assign node4784 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node4787 = (inp[2]) ? node4791 : node4788;
												assign node4788 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node4791 = (inp[5]) ? node4797 : node4792;
													assign node4792 = (inp[0]) ? node4794 : 8'b00101010;
														assign node4794 = (inp[6]) ? 8'b00101010 : 8'b00011111;
													assign node4797 = (inp[6]) ? 8'b00011111 : node4798;
														assign node4798 = (inp[0]) ? 8'b00011111 : 8'b00101010;
									assign node4802 = (inp[0]) ? node4842 : node4803;
										assign node4803 = (inp[12]) ? node4821 : node4804;
											assign node4804 = (inp[6]) ? node4812 : node4805;
												assign node4805 = (inp[2]) ? 8'b00011111 : node4806;
													assign node4806 = (inp[3]) ? node4808 : 8'b00101010;
														assign node4808 = (inp[5]) ? 8'b00001111 : 8'b00101010;
												assign node4812 = (inp[3]) ? node4818 : node4813;
													assign node4813 = (inp[5]) ? node4815 : 8'b00011111;
														assign node4815 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node4818 = (inp[5]) ? 8'b00011110 : 8'b00011111;
											assign node4821 = (inp[5]) ? node4827 : node4822;
												assign node4822 = (inp[2]) ? 8'b00101010 : node4823;
													assign node4823 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node4827 = (inp[3]) ? node4835 : node4828;
													assign node4828 = (inp[2]) ? node4832 : node4829;
														assign node4829 = (inp[6]) ? 8'b00101010 : 8'b00111010;
														assign node4832 = (inp[6]) ? 8'b00011111 : 8'b00101010;
													assign node4835 = (inp[2]) ? node4839 : node4836;
														assign node4836 = (inp[6]) ? 8'b00001111 : 8'b00011111;
														assign node4839 = (inp[6]) ? 8'b00011110 : 8'b00001111;
										assign node4842 = (inp[2]) ? node4864 : node4843;
											assign node4843 = (inp[3]) ? node4851 : node4844;
												assign node4844 = (inp[12]) ? node4848 : node4845;
													assign node4845 = (inp[6]) ? 8'b00011110 : 8'b00001111;
													assign node4848 = (inp[6]) ? 8'b00001111 : 8'b00011111;
												assign node4851 = (inp[5]) ? node4859 : node4852;
													assign node4852 = (inp[12]) ? node4856 : node4853;
														assign node4853 = (inp[6]) ? 8'b00011111 : 8'b00101010;
														assign node4856 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node4859 = (inp[12]) ? node4861 : 8'b00011110;
														assign node4861 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node4864 = (inp[5]) ? node4878 : node4865;
												assign node4865 = (inp[3]) ? node4873 : node4866;
													assign node4866 = (inp[12]) ? node4870 : node4867;
														assign node4867 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node4870 = (inp[6]) ? 8'b00001111 : 8'b00011110;
													assign node4873 = (inp[6]) ? 8'b00011111 : node4874;
														assign node4874 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node4878 = (inp[12]) ? 8'b00011110 : 8'b00001110;
							assign node4881 = (inp[5]) ? node4987 : node4882;
								assign node4882 = (inp[12]) ? node4934 : node4883;
									assign node4883 = (inp[6]) ? node4917 : node4884;
										assign node4884 = (inp[2]) ? node4900 : node4885;
											assign node4885 = (inp[0]) ? node4891 : node4886;
												assign node4886 = (inp[1]) ? 8'b00101010 : node4887;
													assign node4887 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node4891 = (inp[3]) ? node4897 : node4892;
													assign node4892 = (inp[1]) ? node4894 : 8'b00101011;
														assign node4894 = (inp[10]) ? 8'b00001111 : 8'b00001011;
													assign node4897 = (inp[10]) ? 8'b00101010 : 8'b00001110;
											assign node4900 = (inp[3]) ? node4912 : node4901;
												assign node4901 = (inp[0]) ? node4905 : node4902;
													assign node4902 = (inp[1]) ? 8'b00011111 : 8'b00111010;
													assign node4905 = (inp[1]) ? node4909 : node4906;
														assign node4906 = (inp[10]) ? 8'b00101010 : 8'b00001110;
														assign node4909 = (inp[10]) ? 8'b00001110 : 8'b00001010;
												assign node4912 = (inp[0]) ? node4914 : 8'b00011111;
													assign node4914 = (inp[10]) ? 8'b00001111 : 8'b00001011;
										assign node4917 = (inp[3]) ? node4929 : node4918;
											assign node4918 = (inp[1]) ? node4924 : node4919;
												assign node4919 = (inp[0]) ? node4921 : 8'b00111010;
													assign node4921 = (inp[10]) ? 8'b00111010 : 8'b00011110;
												assign node4924 = (inp[0]) ? node4926 : 8'b00011111;
													assign node4926 = (inp[10]) ? 8'b00011110 : 8'b00011010;
											assign node4929 = (inp[0]) ? node4931 : 8'b00011111;
												assign node4931 = (inp[10]) ? 8'b00011111 : 8'b00011011;
									assign node4934 = (inp[0]) ? node4950 : node4935;
										assign node4935 = (inp[2]) ? node4945 : node4936;
											assign node4936 = (inp[6]) ? node4942 : node4937;
												assign node4937 = (inp[1]) ? 8'b00111010 : node4938;
													assign node4938 = (inp[3]) ? 8'b00111010 : 8'b00111011;
												assign node4942 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node4945 = (inp[1]) ? 8'b00101010 : node4946;
												assign node4946 = (inp[3]) ? 8'b00101010 : 8'b00101011;
										assign node4950 = (inp[6]) ? node4976 : node4951;
											assign node4951 = (inp[10]) ? node4965 : node4952;
												assign node4952 = (inp[1]) ? node4960 : node4953;
													assign node4953 = (inp[2]) ? node4957 : node4954;
														assign node4954 = (inp[3]) ? 8'b00011110 : 8'b00011111;
														assign node4957 = (inp[3]) ? 8'b00011011 : 8'b00011110;
													assign node4960 = (inp[3]) ? 8'b00011011 : node4961;
														assign node4961 = (inp[2]) ? 8'b00011010 : 8'b00011011;
												assign node4965 = (inp[2]) ? node4971 : node4966;
													assign node4966 = (inp[3]) ? 8'b00111010 : node4967;
														assign node4967 = (inp[1]) ? 8'b00011111 : 8'b00111011;
													assign node4971 = (inp[3]) ? 8'b00011111 : node4972;
														assign node4972 = (inp[1]) ? 8'b00011110 : 8'b00111010;
											assign node4976 = (inp[3]) ? node4984 : node4977;
												assign node4977 = (inp[10]) ? node4981 : node4978;
													assign node4978 = (inp[1]) ? 8'b00001011 : 8'b00001111;
													assign node4981 = (inp[1]) ? 8'b00001111 : 8'b00101011;
												assign node4984 = (inp[10]) ? 8'b00101010 : 8'b00001110;
								assign node4987 = (inp[1]) ? node5075 : node4988;
									assign node4988 = (inp[10]) ? node5040 : node4989;
										assign node4989 = (inp[0]) ? node5019 : node4990;
											assign node4990 = (inp[3]) ? node5004 : node4991;
												assign node4991 = (inp[6]) ? node4997 : node4992;
													assign node4992 = (inp[12]) ? node4994 : 8'b00101011;
														assign node4994 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node4997 = (inp[12]) ? node5001 : node4998;
														assign node4998 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node5001 = (inp[2]) ? 8'b00111010 : 8'b00101011;
												assign node5004 = (inp[12]) ? node5012 : node5005;
													assign node5005 = (inp[6]) ? node5009 : node5006;
														assign node5006 = (inp[2]) ? 8'b00011111 : 8'b00101010;
														assign node5009 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node5012 = (inp[6]) ? node5016 : node5013;
														assign node5013 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node5016 = (inp[2]) ? 8'b00011111 : 8'b00101010;
											assign node5019 = (inp[12]) ? node5031 : node5020;
												assign node5020 = (inp[3]) ? node5026 : node5021;
													assign node5021 = (inp[6]) ? 8'b00011110 : node5022;
														assign node5022 = (inp[2]) ? 8'b00001110 : 8'b00001111;
													assign node5026 = (inp[2]) ? 8'b00001011 : node5027;
														assign node5027 = (inp[6]) ? 8'b00011011 : 8'b00001110;
												assign node5031 = (inp[2]) ? 8'b00011110 : node5032;
													assign node5032 = (inp[6]) ? node5036 : node5033;
														assign node5033 = (inp[3]) ? 8'b00011110 : 8'b00011111;
														assign node5036 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node5040 = (inp[3]) ? node5060 : node5041;
											assign node5041 = (inp[2]) ? node5049 : node5042;
												assign node5042 = (inp[6]) ? node5046 : node5043;
													assign node5043 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node5046 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node5049 = (inp[12]) ? node5055 : node5050;
													assign node5050 = (inp[6]) ? 8'b00001110 : node5051;
														assign node5051 = (inp[0]) ? 8'b00001110 : 8'b00011110;
													assign node5055 = (inp[0]) ? 8'b00011110 : node5056;
														assign node5056 = (inp[6]) ? 8'b00011110 : 8'b00001111;
											assign node5060 = (inp[2]) ? node5068 : node5061;
												assign node5061 = (inp[6]) ? node5065 : node5062;
													assign node5062 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node5065 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node5068 = (inp[12]) ? node5070 : 8'b00001011;
													assign node5070 = (inp[6]) ? 8'b00011011 : node5071;
														assign node5071 = (inp[0]) ? 8'b00011011 : 8'b00001110;
									assign node5075 = (inp[0]) ? node5133 : node5076;
										assign node5076 = (inp[10]) ? node5106 : node5077;
											assign node5077 = (inp[3]) ? node5091 : node5078;
												assign node5078 = (inp[2]) ? node5084 : node5079;
													assign node5079 = (inp[12]) ? node5081 : 8'b00101010;
														assign node5081 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node5084 = (inp[6]) ? node5088 : node5085;
														assign node5085 = (inp[12]) ? 8'b00101010 : 8'b00011111;
														assign node5088 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node5091 = (inp[12]) ? node5099 : node5092;
													assign node5092 = (inp[2]) ? node5096 : node5093;
														assign node5093 = (inp[6]) ? 8'b00011110 : 8'b00001111;
														assign node5096 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node5099 = (inp[2]) ? node5103 : node5100;
														assign node5100 = (inp[6]) ? 8'b00001111 : 8'b00011111;
														assign node5103 = (inp[6]) ? 8'b00011110 : 8'b00001111;
											assign node5106 = (inp[3]) ? node5118 : node5107;
												assign node5107 = (inp[6]) ? node5113 : node5108;
													assign node5108 = (inp[12]) ? node5110 : 8'b00011011;
														assign node5110 = (inp[2]) ? 8'b00001110 : 8'b00011110;
													assign node5113 = (inp[2]) ? node5115 : 8'b00011011;
														assign node5115 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node5118 = (inp[12]) ? node5126 : node5119;
													assign node5119 = (inp[6]) ? node5123 : node5120;
														assign node5120 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node5123 = (inp[2]) ? 8'b00001010 : 8'b00011010;
													assign node5126 = (inp[6]) ? node5130 : node5127;
														assign node5127 = (inp[2]) ? 8'b00001011 : 8'b00011011;
														assign node5130 = (inp[2]) ? 8'b00011010 : 8'b00001011;
										assign node5133 = (inp[2]) ? node5141 : node5134;
											assign node5134 = (inp[6]) ? node5138 : node5135;
												assign node5135 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node5138 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node5141 = (inp[12]) ? 8'b00011010 : 8'b00001010;
					assign node5144 = (inp[8]) ? node5550 : node5145;
						assign node5145 = (inp[10]) ? node5347 : node5146;
							assign node5146 = (inp[11]) ? node5210 : node5147;
								assign node5147 = (inp[6]) ? node5183 : node5148;
									assign node5148 = (inp[0]) ? node5176 : node5149;
										assign node5149 = (inp[2]) ? node5163 : node5150;
											assign node5150 = (inp[5]) ? node5156 : node5151;
												assign node5151 = (inp[1]) ? 8'b00011110 : node5152;
													assign node5152 = (inp[3]) ? 8'b00011110 : 8'b00011111;
												assign node5156 = (inp[3]) ? node5160 : node5157;
													assign node5157 = (inp[1]) ? 8'b00011110 : 8'b00011111;
													assign node5160 = (inp[1]) ? 8'b00011111 : 8'b00011110;
											assign node5163 = (inp[5]) ? node5169 : node5164;
												assign node5164 = (inp[3]) ? 8'b00001110 : node5165;
													assign node5165 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node5169 = (inp[12]) ? node5171 : 8'b00001111;
													assign node5171 = (inp[3]) ? 8'b00001111 : node5172;
														assign node5172 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node5176 = (inp[3]) ? node5178 : 8'b00011111;
											assign node5178 = (inp[1]) ? node5180 : 8'b00011110;
												assign node5180 = (inp[5]) ? 8'b00011111 : 8'b00011110;
									assign node5183 = (inp[3]) ? node5201 : node5184;
										assign node5184 = (inp[0]) ? node5196 : node5185;
											assign node5185 = (inp[1]) ? node5191 : node5186;
												assign node5186 = (inp[2]) ? node5188 : 8'b00001111;
													assign node5188 = (inp[5]) ? 8'b00011111 : 8'b00001111;
												assign node5191 = (inp[2]) ? node5193 : 8'b00001110;
													assign node5193 = (inp[5]) ? 8'b00011110 : 8'b00001110;
											assign node5196 = (inp[2]) ? node5198 : 8'b00001111;
												assign node5198 = (inp[5]) ? 8'b00011111 : 8'b00001111;
										assign node5201 = (inp[5]) ? node5203 : 8'b00001110;
											assign node5203 = (inp[2]) ? node5207 : node5204;
												assign node5204 = (inp[1]) ? 8'b00001111 : 8'b00001110;
												assign node5207 = (inp[1]) ? 8'b00011111 : 8'b00011110;
								assign node5210 = (inp[1]) ? node5270 : node5211;
									assign node5211 = (inp[3]) ? node5243 : node5212;
										assign node5212 = (inp[2]) ? node5220 : node5213;
											assign node5213 = (inp[12]) ? node5217 : node5214;
												assign node5214 = (inp[6]) ? 8'b00011110 : 8'b00001111;
												assign node5217 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node5220 = (inp[12]) ? node5232 : node5221;
												assign node5221 = (inp[0]) ? node5227 : node5222;
													assign node5222 = (inp[5]) ? node5224 : 8'b00011110;
														assign node5224 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node5227 = (inp[6]) ? node5229 : 8'b00001110;
														assign node5229 = (inp[5]) ? 8'b00001110 : 8'b00011110;
												assign node5232 = (inp[5]) ? node5238 : node5233;
													assign node5233 = (inp[6]) ? 8'b00001111 : node5234;
														assign node5234 = (inp[0]) ? 8'b00011110 : 8'b00001111;
													assign node5238 = (inp[6]) ? 8'b00011110 : node5239;
														assign node5239 = (inp[0]) ? 8'b00011110 : 8'b00001111;
										assign node5243 = (inp[2]) ? node5251 : node5244;
											assign node5244 = (inp[12]) ? node5248 : node5245;
												assign node5245 = (inp[6]) ? 8'b00011011 : 8'b00001110;
												assign node5248 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node5251 = (inp[12]) ? node5259 : node5252;
												assign node5252 = (inp[5]) ? node5254 : 8'b00011011;
													assign node5254 = (inp[6]) ? 8'b00001011 : node5255;
														assign node5255 = (inp[0]) ? 8'b00001011 : 8'b00011011;
												assign node5259 = (inp[5]) ? node5265 : node5260;
													assign node5260 = (inp[6]) ? 8'b00001110 : node5261;
														assign node5261 = (inp[0]) ? 8'b00011011 : 8'b00001110;
													assign node5265 = (inp[6]) ? 8'b00011011 : node5266;
														assign node5266 = (inp[0]) ? 8'b00011011 : 8'b00001110;
									assign node5270 = (inp[2]) ? node5310 : node5271;
										assign node5271 = (inp[5]) ? node5291 : node5272;
											assign node5272 = (inp[12]) ? node5280 : node5273;
												assign node5273 = (inp[6]) ? 8'b00011011 : node5274;
													assign node5274 = (inp[0]) ? node5276 : 8'b00001110;
														assign node5276 = (inp[3]) ? 8'b00001110 : 8'b00001011;
												assign node5280 = (inp[6]) ? node5286 : node5281;
													assign node5281 = (inp[0]) ? node5283 : 8'b00011110;
														assign node5283 = (inp[3]) ? 8'b00011110 : 8'b00011011;
													assign node5286 = (inp[0]) ? node5288 : 8'b00001110;
														assign node5288 = (inp[3]) ? 8'b00001110 : 8'b00001011;
											assign node5291 = (inp[0]) ? node5305 : node5292;
												assign node5292 = (inp[3]) ? node5300 : node5293;
													assign node5293 = (inp[6]) ? node5297 : node5294;
														assign node5294 = (inp[12]) ? 8'b00011110 : 8'b00001110;
														assign node5297 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node5300 = (inp[6]) ? 8'b00001011 : node5301;
														assign node5301 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node5305 = (inp[12]) ? node5307 : 8'b00001011;
													assign node5307 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node5310 = (inp[0]) ? node5332 : node5311;
											assign node5311 = (inp[12]) ? node5323 : node5312;
												assign node5312 = (inp[3]) ? node5318 : node5313;
													assign node5313 = (inp[5]) ? node5315 : 8'b00011011;
														assign node5315 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node5318 = (inp[5]) ? node5320 : 8'b00011011;
														assign node5320 = (inp[6]) ? 8'b00001010 : 8'b00011010;
												assign node5323 = (inp[5]) ? node5325 : 8'b00001110;
													assign node5325 = (inp[6]) ? node5329 : node5326;
														assign node5326 = (inp[3]) ? 8'b00001011 : 8'b00001110;
														assign node5329 = (inp[3]) ? 8'b00011010 : 8'b00011011;
											assign node5332 = (inp[12]) ? node5340 : node5333;
												assign node5333 = (inp[5]) ? 8'b00001010 : node5334;
													assign node5334 = (inp[3]) ? 8'b00011011 : node5335;
														assign node5335 = (inp[6]) ? 8'b00011010 : 8'b00001010;
												assign node5340 = (inp[5]) ? 8'b00011010 : node5341;
													assign node5341 = (inp[6]) ? 8'b00001011 : node5342;
														assign node5342 = (inp[3]) ? 8'b00011011 : 8'b00011010;
							assign node5347 = (inp[1]) ? node5435 : node5348;
								assign node5348 = (inp[3]) ? node5384 : node5349;
									assign node5349 = (inp[11]) ? node5361 : node5350;
										assign node5350 = (inp[6]) ? node5356 : node5351;
											assign node5351 = (inp[2]) ? node5353 : 8'b00011011;
												assign node5353 = (inp[0]) ? 8'b00011011 : 8'b00001011;
											assign node5356 = (inp[2]) ? node5358 : 8'b00001011;
												assign node5358 = (inp[5]) ? 8'b00011011 : 8'b00001011;
										assign node5361 = (inp[12]) ? node5373 : node5362;
											assign node5362 = (inp[6]) ? node5368 : node5363;
												assign node5363 = (inp[2]) ? node5365 : 8'b00001011;
													assign node5365 = (inp[0]) ? 8'b00001010 : 8'b00011010;
												assign node5368 = (inp[5]) ? node5370 : 8'b00011010;
													assign node5370 = (inp[2]) ? 8'b00001010 : 8'b00011010;
											assign node5373 = (inp[6]) ? node5379 : node5374;
												assign node5374 = (inp[2]) ? node5376 : 8'b00011011;
													assign node5376 = (inp[0]) ? 8'b00011010 : 8'b00001011;
												assign node5379 = (inp[2]) ? node5381 : 8'b00001011;
													assign node5381 = (inp[5]) ? 8'b00011010 : 8'b00001011;
									assign node5384 = (inp[11]) ? node5408 : node5385;
										assign node5385 = (inp[2]) ? node5391 : node5386;
											assign node5386 = (inp[6]) ? node5388 : 8'b00011010;
												assign node5388 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node5391 = (inp[0]) ? node5401 : node5392;
												assign node5392 = (inp[5]) ? node5396 : node5393;
													assign node5393 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5396 = (inp[6]) ? 8'b10010000 : node5397;
														assign node5397 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5401 = (inp[6]) ? node5403 : 8'b10010000;
													assign node5403 = (inp[5]) ? 8'b10010000 : node5404;
														assign node5404 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node5408 = (inp[2]) ? node5416 : node5409;
											assign node5409 = (inp[6]) ? node5413 : node5410;
												assign node5410 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node5413 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node5416 = (inp[12]) ? node5428 : node5417;
												assign node5417 = (inp[5]) ? node5423 : node5418;
													assign node5418 = (inp[0]) ? node5420 : 8'b11110111;
														assign node5420 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node5423 = (inp[0]) ? 8'b10100101 : node5424;
														assign node5424 = (inp[6]) ? 8'b10100101 : 8'b11110111;
												assign node5428 = (inp[5]) ? 8'b11110101 : node5429;
													assign node5429 = (inp[0]) ? node5431 : 8'b00000010;
														assign node5431 = (inp[6]) ? 8'b00000010 : 8'b11110101;
								assign node5435 = (inp[11]) ? node5481 : node5436;
									assign node5436 = (inp[5]) ? node5458 : node5437;
										assign node5437 = (inp[6]) ? node5451 : node5438;
											assign node5438 = (inp[2]) ? node5444 : node5439;
												assign node5439 = (inp[3]) ? 8'b00011010 : node5440;
													assign node5440 = (inp[0]) ? 8'b10011001 : 8'b00011010;
												assign node5444 = (inp[0]) ? node5448 : node5445;
													assign node5445 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5448 = (inp[12]) ? 8'b10010001 : 8'b10010000;
											assign node5451 = (inp[3]) ? node5455 : node5452;
												assign node5452 = (inp[0]) ? 8'b10000001 : 8'b10000010;
												assign node5455 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node5458 = (inp[0]) ? node5476 : node5459;
											assign node5459 = (inp[3]) ? node5469 : node5460;
												assign node5460 = (inp[6]) ? node5466 : node5461;
													assign node5461 = (inp[2]) ? node5463 : 8'b00011010;
														assign node5463 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5466 = (inp[2]) ? 8'b10010000 : 8'b10000010;
												assign node5469 = (inp[6]) ? node5473 : node5470;
													assign node5470 = (inp[2]) ? 8'b10000001 : 8'b10011001;
													assign node5473 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node5476 = (inp[2]) ? 8'b10010001 : node5477;
												assign node5477 = (inp[6]) ? 8'b10000001 : 8'b10011001;
									assign node5481 = (inp[5]) ? node5515 : node5482;
										assign node5482 = (inp[12]) ? node5500 : node5483;
											assign node5483 = (inp[6]) ? node5495 : node5484;
												assign node5484 = (inp[2]) ? node5490 : node5485;
													assign node5485 = (inp[0]) ? node5487 : 8'b00001010;
														assign node5487 = (inp[3]) ? 8'b00001010 : 8'b10101101;
													assign node5490 = (inp[0]) ? node5492 : 8'b11110111;
														assign node5492 = (inp[3]) ? 8'b10100101 : 8'b10100100;
												assign node5495 = (inp[3]) ? 8'b11110111 : node5496;
													assign node5496 = (inp[0]) ? 8'b10110100 : 8'b11110111;
											assign node5500 = (inp[0]) ? node5506 : node5501;
												assign node5501 = (inp[6]) ? 8'b00000010 : node5502;
													assign node5502 = (inp[2]) ? 8'b00000010 : 8'b00011010;
												assign node5506 = (inp[6]) ? node5512 : node5507;
													assign node5507 = (inp[2]) ? node5509 : 8'b11111101;
														assign node5509 = (inp[3]) ? 8'b11110101 : 8'b10110100;
													assign node5512 = (inp[3]) ? 8'b00000010 : 8'b10100101;
										assign node5515 = (inp[2]) ? node5531 : node5516;
											assign node5516 = (inp[6]) ? node5524 : node5517;
												assign node5517 = (inp[12]) ? node5519 : 8'b10101101;
													assign node5519 = (inp[0]) ? 8'b11111101 : node5520;
														assign node5520 = (inp[3]) ? 8'b11111101 : 8'b00011010;
												assign node5524 = (inp[12]) ? 8'b10100101 : node5525;
													assign node5525 = (inp[0]) ? 8'b10110100 : node5526;
														assign node5526 = (inp[3]) ? 8'b10110100 : 8'b11110111;
											assign node5531 = (inp[12]) ? node5539 : node5532;
												assign node5532 = (inp[0]) ? 8'b10100100 : node5533;
													assign node5533 = (inp[3]) ? node5535 : 8'b10100101;
														assign node5535 = (inp[6]) ? 8'b10100100 : 8'b10110100;
												assign node5539 = (inp[6]) ? node5545 : node5540;
													assign node5540 = (inp[3]) ? node5542 : 8'b00000010;
														assign node5542 = (inp[0]) ? 8'b10110100 : 8'b10100101;
													assign node5545 = (inp[3]) ? 8'b10110100 : node5546;
														assign node5546 = (inp[0]) ? 8'b10110100 : 8'b11110101;
						assign node5550 = (inp[5]) ? node5744 : node5551;
							assign node5551 = (inp[0]) ? node5605 : node5552;
								assign node5552 = (inp[12]) ? node5588 : node5553;
									assign node5553 = (inp[11]) ? node5571 : node5554;
										assign node5554 = (inp[6]) ? node5566 : node5555;
											assign node5555 = (inp[2]) ? node5561 : node5556;
												assign node5556 = (inp[3]) ? 8'b00011010 : node5557;
													assign node5557 = (inp[1]) ? 8'b00011010 : 8'b00011011;
												assign node5561 = (inp[1]) ? 8'b10000010 : node5562;
													assign node5562 = (inp[3]) ? 8'b10000010 : 8'b00001011;
											assign node5566 = (inp[1]) ? 8'b10000010 : node5567;
												assign node5567 = (inp[3]) ? 8'b10000010 : 8'b00001011;
										assign node5571 = (inp[6]) ? node5583 : node5572;
											assign node5572 = (inp[2]) ? node5578 : node5573;
												assign node5573 = (inp[1]) ? 8'b00001010 : node5574;
													assign node5574 = (inp[3]) ? 8'b00001010 : 8'b00001011;
												assign node5578 = (inp[3]) ? 8'b11110111 : node5579;
													assign node5579 = (inp[1]) ? 8'b11110111 : 8'b00011010;
											assign node5583 = (inp[1]) ? 8'b11110111 : node5584;
												assign node5584 = (inp[3]) ? 8'b11110111 : 8'b00011010;
									assign node5588 = (inp[6]) ? node5600 : node5589;
										assign node5589 = (inp[2]) ? node5595 : node5590;
											assign node5590 = (inp[3]) ? 8'b00011010 : node5591;
												assign node5591 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node5595 = (inp[3]) ? 8'b00000010 : node5596;
												assign node5596 = (inp[1]) ? 8'b00000010 : 8'b00001011;
										assign node5600 = (inp[1]) ? 8'b00000010 : node5601;
											assign node5601 = (inp[3]) ? 8'b00000010 : 8'b00001011;
								assign node5605 = (inp[10]) ? node5663 : node5606;
									assign node5606 = (inp[11]) ? node5622 : node5607;
										assign node5607 = (inp[6]) ? node5617 : node5608;
											assign node5608 = (inp[3]) ? node5614 : node5609;
												assign node5609 = (inp[1]) ? node5611 : 8'b10011101;
													assign node5611 = (inp[2]) ? 8'b10010101 : 8'b10011101;
												assign node5614 = (inp[2]) ? 8'b10010100 : 8'b10011100;
											assign node5617 = (inp[3]) ? 8'b10000100 : node5618;
												assign node5618 = (inp[1]) ? 8'b10000101 : 8'b10001101;
										assign node5622 = (inp[1]) ? node5642 : node5623;
											assign node5623 = (inp[3]) ? node5631 : node5624;
												assign node5624 = (inp[12]) ? node5628 : node5625;
													assign node5625 = (inp[2]) ? 8'b10101100 : 8'b10111100;
													assign node5628 = (inp[6]) ? 8'b10101101 : 8'b10111100;
												assign node5631 = (inp[2]) ? node5637 : node5632;
													assign node5632 = (inp[6]) ? 8'b10110001 : node5633;
														assign node5633 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node5637 = (inp[6]) ? 8'b10100100 : node5638;
														assign node5638 = (inp[12]) ? 8'b10110001 : 8'b10100001;
											assign node5642 = (inp[6]) ? node5656 : node5643;
												assign node5643 = (inp[2]) ? node5651 : node5644;
													assign node5644 = (inp[3]) ? node5648 : node5645;
														assign node5645 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node5648 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node5651 = (inp[3]) ? node5653 : 8'b10110000;
														assign node5653 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node5656 = (inp[12]) ? node5660 : node5657;
													assign node5657 = (inp[3]) ? 8'b10110001 : 8'b10110000;
													assign node5660 = (inp[3]) ? 8'b10100100 : 8'b10100001;
									assign node5663 = (inp[1]) ? node5705 : node5664;
										assign node5664 = (inp[3]) ? node5680 : node5665;
											assign node5665 = (inp[6]) ? node5675 : node5666;
												assign node5666 = (inp[11]) ? node5668 : 8'b00011011;
													assign node5668 = (inp[12]) ? node5672 : node5669;
														assign node5669 = (inp[2]) ? 8'b00001010 : 8'b00001011;
														assign node5672 = (inp[2]) ? 8'b00011010 : 8'b00011011;
												assign node5675 = (inp[12]) ? 8'b00001011 : node5676;
													assign node5676 = (inp[11]) ? 8'b00011010 : 8'b00001011;
											assign node5680 = (inp[2]) ? node5692 : node5681;
												assign node5681 = (inp[6]) ? node5687 : node5682;
													assign node5682 = (inp[12]) ? 8'b00011010 : node5683;
														assign node5683 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node5687 = (inp[12]) ? 8'b00000010 : node5688;
														assign node5688 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node5692 = (inp[11]) ? node5698 : node5693;
													assign node5693 = (inp[6]) ? node5695 : 8'b10010000;
														assign node5695 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5698 = (inp[6]) ? node5702 : node5699;
														assign node5699 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node5702 = (inp[12]) ? 8'b00000010 : 8'b11110111;
										assign node5705 = (inp[3]) ? node5723 : node5706;
											assign node5706 = (inp[11]) ? node5712 : node5707;
												assign node5707 = (inp[6]) ? 8'b10000001 : node5708;
													assign node5708 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node5712 = (inp[2]) ? node5716 : node5713;
													assign node5713 = (inp[6]) ? 8'b10100101 : 8'b11111101;
													assign node5716 = (inp[6]) ? node5720 : node5717;
														assign node5717 = (inp[12]) ? 8'b10110100 : 8'b10100100;
														assign node5720 = (inp[12]) ? 8'b10100101 : 8'b10110100;
											assign node5723 = (inp[2]) ? node5733 : node5724;
												assign node5724 = (inp[6]) ? node5730 : node5725;
													assign node5725 = (inp[12]) ? 8'b00011010 : node5726;
														assign node5726 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node5730 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5733 = (inp[11]) ? node5739 : node5734;
													assign node5734 = (inp[6]) ? node5736 : 8'b10010000;
														assign node5736 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5739 = (inp[6]) ? 8'b11110111 : node5740;
														assign node5740 = (inp[12]) ? 8'b11110101 : 8'b10100101;
							assign node5744 = (inp[11]) ? node5852 : node5745;
								assign node5745 = (inp[0]) ? node5823 : node5746;
									assign node5746 = (inp[10]) ? node5788 : node5747;
										assign node5747 = (inp[1]) ? node5771 : node5748;
											assign node5748 = (inp[3]) ? node5762 : node5749;
												assign node5749 = (inp[12]) ? node5755 : node5750;
													assign node5750 = (inp[2]) ? node5752 : 8'b00001011;
														assign node5752 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node5755 = (inp[2]) ? node5759 : node5756;
														assign node5756 = (inp[6]) ? 8'b00001011 : 8'b00011011;
														assign node5759 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node5762 = (inp[2]) ? node5768 : node5763;
													assign node5763 = (inp[6]) ? node5765 : 8'b00011010;
														assign node5765 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5768 = (inp[6]) ? 8'b10010000 : 8'b10000010;
											assign node5771 = (inp[3]) ? node5781 : node5772;
												assign node5772 = (inp[2]) ? node5778 : node5773;
													assign node5773 = (inp[6]) ? node5775 : 8'b00011010;
														assign node5775 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5778 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node5781 = (inp[2]) ? node5785 : node5782;
													assign node5782 = (inp[6]) ? 8'b10000001 : 8'b10011001;
													assign node5785 = (inp[6]) ? 8'b10010001 : 8'b10000001;
										assign node5788 = (inp[1]) ? node5804 : node5789;
											assign node5789 = (inp[3]) ? node5797 : node5790;
												assign node5790 = (inp[6]) ? node5794 : node5791;
													assign node5791 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node5794 = (inp[2]) ? 8'b10011101 : 8'b10001101;
												assign node5797 = (inp[2]) ? node5801 : node5798;
													assign node5798 = (inp[6]) ? 8'b10000100 : 8'b10011100;
													assign node5801 = (inp[6]) ? 8'b10010100 : 8'b10000100;
											assign node5804 = (inp[3]) ? node5812 : node5805;
												assign node5805 = (inp[6]) ? node5809 : node5806;
													assign node5806 = (inp[2]) ? 8'b10000100 : 8'b10011100;
													assign node5809 = (inp[2]) ? 8'b10010100 : 8'b10000100;
												assign node5812 = (inp[12]) ? node5818 : node5813;
													assign node5813 = (inp[6]) ? node5815 : 8'b10000101;
														assign node5815 = (inp[2]) ? 8'b10010101 : 8'b10000101;
													assign node5818 = (inp[6]) ? node5820 : 8'b10011101;
														assign node5820 = (inp[2]) ? 8'b10010101 : 8'b10000101;
									assign node5823 = (inp[6]) ? node5837 : node5824;
										assign node5824 = (inp[2]) ? node5830 : node5825;
											assign node5825 = (inp[3]) ? node5827 : 8'b10011101;
												assign node5827 = (inp[1]) ? 8'b10011101 : 8'b10011100;
											assign node5830 = (inp[3]) ? node5834 : node5831;
												assign node5831 = (inp[1]) ? 8'b10010101 : 8'b10011101;
												assign node5834 = (inp[1]) ? 8'b10010101 : 8'b10010100;
										assign node5837 = (inp[2]) ? node5845 : node5838;
											assign node5838 = (inp[3]) ? node5842 : node5839;
												assign node5839 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node5842 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node5845 = (inp[3]) ? node5849 : node5846;
												assign node5846 = (inp[1]) ? 8'b10010101 : 8'b10011101;
												assign node5849 = (inp[1]) ? 8'b10010101 : 8'b10010100;
								assign node5852 = (inp[1]) ? node5924 : node5853;
									assign node5853 = (inp[3]) ? node5891 : node5854;
										assign node5854 = (inp[0]) ? node5880 : node5855;
											assign node5855 = (inp[10]) ? node5867 : node5856;
												assign node5856 = (inp[2]) ? node5860 : node5857;
													assign node5857 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node5860 = (inp[12]) ? node5864 : node5861;
														assign node5861 = (inp[6]) ? 8'b00001010 : 8'b00011010;
														assign node5864 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node5867 = (inp[12]) ? node5873 : node5868;
													assign node5868 = (inp[6]) ? node5870 : 8'b10111100;
														assign node5870 = (inp[2]) ? 8'b10101100 : 8'b10111100;
													assign node5873 = (inp[6]) ? node5877 : node5874;
														assign node5874 = (inp[2]) ? 8'b10101101 : 8'b11111101;
														assign node5877 = (inp[2]) ? 8'b10111100 : 8'b10101101;
											assign node5880 = (inp[2]) ? node5888 : node5881;
												assign node5881 = (inp[12]) ? node5885 : node5882;
													assign node5882 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node5885 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node5888 = (inp[12]) ? 8'b10111100 : 8'b10101100;
										assign node5891 = (inp[2]) ? node5911 : node5892;
											assign node5892 = (inp[6]) ? node5904 : node5893;
												assign node5893 = (inp[0]) ? node5901 : node5894;
													assign node5894 = (inp[10]) ? node5898 : node5895;
														assign node5895 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node5898 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node5901 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node5904 = (inp[12]) ? node5906 : 8'b10110001;
													assign node5906 = (inp[0]) ? 8'b10100100 : node5907;
														assign node5907 = (inp[10]) ? 8'b10100100 : 8'b00000010;
											assign node5911 = (inp[0]) ? node5921 : node5912;
												assign node5912 = (inp[10]) ? node5916 : node5913;
													assign node5913 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node5916 = (inp[12]) ? node5918 : 8'b10110001;
														assign node5918 = (inp[6]) ? 8'b10110001 : 8'b10100100;
												assign node5921 = (inp[12]) ? 8'b10110001 : 8'b10100001;
									assign node5924 = (inp[2]) ? node5958 : node5925;
										assign node5925 = (inp[6]) ? node5943 : node5926;
											assign node5926 = (inp[12]) ? node5936 : node5927;
												assign node5927 = (inp[0]) ? 8'b10101001 : node5928;
													assign node5928 = (inp[3]) ? node5932 : node5929;
														assign node5929 = (inp[10]) ? 8'b10101100 : 8'b00001010;
														assign node5932 = (inp[10]) ? 8'b10101001 : 8'b10101101;
												assign node5936 = (inp[0]) ? 8'b10111001 : node5937;
													assign node5937 = (inp[10]) ? node5939 : 8'b11111101;
														assign node5939 = (inp[3]) ? 8'b10111001 : 8'b10111100;
											assign node5943 = (inp[12]) ? node5951 : node5944;
												assign node5944 = (inp[0]) ? 8'b10110000 : node5945;
													assign node5945 = (inp[10]) ? node5947 : 8'b11110111;
														assign node5947 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node5951 = (inp[0]) ? 8'b10100001 : node5952;
													assign node5952 = (inp[3]) ? node5954 : 8'b00000010;
														assign node5954 = (inp[10]) ? 8'b10100001 : 8'b10100101;
										assign node5958 = (inp[0]) ? node5986 : node5959;
											assign node5959 = (inp[10]) ? node5971 : node5960;
												assign node5960 = (inp[3]) ? node5966 : node5961;
													assign node5961 = (inp[6]) ? node5963 : 8'b11110111;
														assign node5963 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node5966 = (inp[12]) ? 8'b10100101 : node5967;
														assign node5967 = (inp[6]) ? 8'b10100100 : 8'b10110100;
												assign node5971 = (inp[3]) ? node5979 : node5972;
													assign node5972 = (inp[6]) ? node5976 : node5973;
														assign node5973 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node5976 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node5979 = (inp[6]) ? node5983 : node5980;
														assign node5980 = (inp[12]) ? 8'b10100001 : 8'b10110000;
														assign node5983 = (inp[12]) ? 8'b10110000 : 8'b10100000;
											assign node5986 = (inp[12]) ? 8'b10110000 : 8'b10100000;
				assign node5989 = (inp[5]) ? node6601 : node5990;
					assign node5990 = (inp[0]) ? node6152 : node5991;
						assign node5991 = (inp[12]) ? node6099 : node5992;
							assign node5992 = (inp[11]) ? node6046 : node5993;
								assign node5993 = (inp[1]) ? node6029 : node5994;
									assign node5994 = (inp[3]) ? node6012 : node5995;
										assign node5995 = (inp[6]) ? node6007 : node5996;
											assign node5996 = (inp[2]) ? node6002 : node5997;
												assign node5997 = (inp[8]) ? 8'b00011011 : node5998;
													assign node5998 = (inp[10]) ? 8'b00011011 : 8'b00011111;
												assign node6002 = (inp[10]) ? 8'b00001011 : node6003;
													assign node6003 = (inp[8]) ? 8'b00001011 : 8'b00001111;
											assign node6007 = (inp[8]) ? 8'b00001011 : node6008;
												assign node6008 = (inp[10]) ? 8'b00001011 : 8'b00001111;
										assign node6012 = (inp[8]) ? node6024 : node6013;
											assign node6013 = (inp[10]) ? node6019 : node6014;
												assign node6014 = (inp[6]) ? 8'b00001110 : node6015;
													assign node6015 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node6019 = (inp[2]) ? 8'b10000010 : node6020;
													assign node6020 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node6024 = (inp[6]) ? 8'b10000010 : node6025;
												assign node6025 = (inp[2]) ? 8'b10000010 : 8'b00011010;
									assign node6029 = (inp[6]) ? node6041 : node6030;
										assign node6030 = (inp[2]) ? node6036 : node6031;
											assign node6031 = (inp[10]) ? 8'b00011010 : node6032;
												assign node6032 = (inp[8]) ? 8'b00011010 : 8'b00011110;
											assign node6036 = (inp[8]) ? 8'b10000010 : node6037;
												assign node6037 = (inp[10]) ? 8'b10000010 : 8'b00001110;
										assign node6041 = (inp[10]) ? 8'b10000010 : node6042;
											assign node6042 = (inp[8]) ? 8'b10000010 : 8'b00001110;
								assign node6046 = (inp[2]) ? node6082 : node6047;
									assign node6047 = (inp[6]) ? node6065 : node6048;
										assign node6048 = (inp[10]) ? node6060 : node6049;
											assign node6049 = (inp[8]) ? node6055 : node6050;
												assign node6050 = (inp[1]) ? 8'b00001110 : node6051;
													assign node6051 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node6055 = (inp[1]) ? 8'b00001010 : node6056;
													assign node6056 = (inp[9]) ? 8'b00001011 : 8'b00001010;
											assign node6060 = (inp[1]) ? 8'b00001010 : node6061;
												assign node6061 = (inp[3]) ? 8'b00001010 : 8'b00001011;
										assign node6065 = (inp[8]) ? node6077 : node6066;
											assign node6066 = (inp[10]) ? node6072 : node6067;
												assign node6067 = (inp[1]) ? 8'b00011011 : node6068;
													assign node6068 = (inp[3]) ? 8'b00011011 : 8'b00011110;
												assign node6072 = (inp[3]) ? 8'b11110111 : node6073;
													assign node6073 = (inp[1]) ? 8'b11110111 : 8'b00011010;
											assign node6077 = (inp[3]) ? 8'b11110111 : node6078;
												assign node6078 = (inp[1]) ? 8'b11110111 : 8'b00011010;
									assign node6082 = (inp[3]) ? node6094 : node6083;
										assign node6083 = (inp[1]) ? node6089 : node6084;
											assign node6084 = (inp[8]) ? 8'b00011010 : node6085;
												assign node6085 = (inp[10]) ? 8'b00011010 : 8'b00011110;
											assign node6089 = (inp[8]) ? 8'b11110111 : node6090;
												assign node6090 = (inp[10]) ? 8'b11110111 : 8'b00011011;
										assign node6094 = (inp[10]) ? 8'b11110111 : node6095;
											assign node6095 = (inp[8]) ? 8'b11110111 : 8'b00011011;
							assign node6099 = (inp[6]) ? node6135 : node6100;
								assign node6100 = (inp[2]) ? node6118 : node6101;
									assign node6101 = (inp[10]) ? node6113 : node6102;
										assign node6102 = (inp[8]) ? node6108 : node6103;
											assign node6103 = (inp[3]) ? 8'b00011110 : node6104;
												assign node6104 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node6108 = (inp[3]) ? 8'b00011010 : node6109;
												assign node6109 = (inp[1]) ? 8'b00011010 : 8'b00011011;
										assign node6113 = (inp[1]) ? 8'b00011010 : node6114;
											assign node6114 = (inp[3]) ? 8'b00011010 : 8'b00011011;
									assign node6118 = (inp[3]) ? node6130 : node6119;
										assign node6119 = (inp[1]) ? node6125 : node6120;
											assign node6120 = (inp[8]) ? 8'b00001011 : node6121;
												assign node6121 = (inp[10]) ? 8'b00001011 : 8'b00001111;
											assign node6125 = (inp[10]) ? 8'b00000010 : node6126;
												assign node6126 = (inp[8]) ? 8'b00000010 : 8'b00001110;
										assign node6130 = (inp[8]) ? 8'b00000010 : node6131;
											assign node6131 = (inp[10]) ? 8'b00000010 : 8'b00001110;
								assign node6135 = (inp[8]) ? node6147 : node6136;
									assign node6136 = (inp[10]) ? node6142 : node6137;
										assign node6137 = (inp[1]) ? 8'b00001110 : node6138;
											assign node6138 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node6142 = (inp[3]) ? 8'b00000010 : node6143;
											assign node6143 = (inp[1]) ? 8'b00000010 : 8'b00001011;
									assign node6147 = (inp[3]) ? 8'b00000010 : node6148;
										assign node6148 = (inp[1]) ? 8'b00000010 : 8'b00001011;
						assign node6152 = (inp[9]) ? node6324 : node6153;
							assign node6153 = (inp[3]) ? node6263 : node6154;
								assign node6154 = (inp[11]) ? node6178 : node6155;
									assign node6155 = (inp[10]) ? node6169 : node6156;
										assign node6156 = (inp[6]) ? node6164 : node6157;
											assign node6157 = (inp[8]) ? node6159 : 8'b11111101;
												assign node6159 = (inp[2]) ? node6161 : 8'b11111101;
													assign node6161 = (inp[1]) ? 8'b11110101 : 8'b11111101;
											assign node6164 = (inp[8]) ? node6166 : 8'b10101101;
												assign node6166 = (inp[1]) ? 8'b10100101 : 8'b10101101;
										assign node6169 = (inp[6]) ? node6175 : node6170;
											assign node6170 = (inp[1]) ? node6172 : 8'b10111001;
												assign node6172 = (inp[2]) ? 8'b10110001 : 8'b10111001;
											assign node6175 = (inp[1]) ? 8'b10100001 : 8'b10101001;
									assign node6178 = (inp[1]) ? node6220 : node6179;
										assign node6179 = (inp[10]) ? node6209 : node6180;
											assign node6180 = (inp[8]) ? node6194 : node6181;
												assign node6181 = (inp[2]) ? node6187 : node6182;
													assign node6182 = (inp[12]) ? node6184 : 8'b10101101;
														assign node6184 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node6187 = (inp[12]) ? node6191 : node6188;
														assign node6188 = (inp[6]) ? 8'b10111100 : 8'b10101100;
														assign node6191 = (inp[6]) ? 8'b10101101 : 8'b10111100;
												assign node6194 = (inp[2]) ? node6202 : node6195;
													assign node6195 = (inp[12]) ? node6199 : node6196;
														assign node6196 = (inp[6]) ? 8'b10011100 : 8'b10001101;
														assign node6199 = (inp[6]) ? 8'b10001101 : 8'b10011101;
													assign node6202 = (inp[12]) ? node6206 : node6203;
														assign node6203 = (inp[6]) ? 8'b10011100 : 8'b10001100;
														assign node6206 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node6209 = (inp[12]) ? node6215 : node6210;
												assign node6210 = (inp[6]) ? 8'b10111000 : node6211;
													assign node6211 = (inp[2]) ? 8'b10101000 : 8'b10101001;
												assign node6215 = (inp[6]) ? 8'b10101001 : node6216;
													assign node6216 = (inp[2]) ? 8'b10111000 : 8'b10111001;
										assign node6220 = (inp[10]) ? node6248 : node6221;
											assign node6221 = (inp[8]) ? node6235 : node6222;
												assign node6222 = (inp[2]) ? node6228 : node6223;
													assign node6223 = (inp[6]) ? 8'b10101001 : node6224;
														assign node6224 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node6228 = (inp[12]) ? node6232 : node6229;
														assign node6229 = (inp[6]) ? 8'b10111000 : 8'b10101000;
														assign node6232 = (inp[6]) ? 8'b10101001 : 8'b10111000;
												assign node6235 = (inp[2]) ? node6241 : node6236;
													assign node6236 = (inp[6]) ? node6238 : 8'b10001001;
														assign node6238 = (inp[12]) ? 8'b10000001 : 8'b10010000;
													assign node6241 = (inp[6]) ? node6245 : node6242;
														assign node6242 = (inp[12]) ? 8'b10010000 : 8'b10000000;
														assign node6245 = (inp[12]) ? 8'b10000001 : 8'b10010000;
											assign node6248 = (inp[2]) ? node6256 : node6249;
												assign node6249 = (inp[6]) ? node6253 : node6250;
													assign node6250 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node6253 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node6256 = (inp[6]) ? node6260 : node6257;
													assign node6257 = (inp[12]) ? 8'b10010100 : 8'b10000100;
													assign node6260 = (inp[12]) ? 8'b10000101 : 8'b10010100;
								assign node6263 = (inp[11]) ? node6279 : node6264;
									assign node6264 = (inp[10]) ? node6274 : node6265;
										assign node6265 = (inp[6]) ? node6271 : node6266;
											assign node6266 = (inp[8]) ? node6268 : 8'b10111100;
												assign node6268 = (inp[2]) ? 8'b10110100 : 8'b10111100;
											assign node6271 = (inp[8]) ? 8'b10100100 : 8'b10101100;
										assign node6274 = (inp[6]) ? 8'b10100000 : node6275;
											assign node6275 = (inp[2]) ? 8'b10110000 : 8'b10111000;
									assign node6279 = (inp[2]) ? node6301 : node6280;
										assign node6280 = (inp[6]) ? node6292 : node6281;
											assign node6281 = (inp[10]) ? node6289 : node6282;
												assign node6282 = (inp[12]) ? node6286 : node6283;
													assign node6283 = (inp[8]) ? 8'b10001100 : 8'b10101100;
													assign node6286 = (inp[8]) ? 8'b10011100 : 8'b10111100;
												assign node6289 = (inp[12]) ? 8'b10111000 : 8'b10101000;
											assign node6292 = (inp[12]) ? node6296 : node6293;
												assign node6293 = (inp[10]) ? 8'b10010101 : 8'b10111001;
												assign node6296 = (inp[10]) ? 8'b10100000 : node6297;
													assign node6297 = (inp[8]) ? 8'b10000100 : 8'b10101100;
										assign node6301 = (inp[10]) ? node6317 : node6302;
											assign node6302 = (inp[8]) ? node6310 : node6303;
												assign node6303 = (inp[12]) ? node6307 : node6304;
													assign node6304 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node6307 = (inp[6]) ? 8'b10101100 : 8'b10111001;
												assign node6310 = (inp[6]) ? node6314 : node6311;
													assign node6311 = (inp[12]) ? 8'b10010001 : 8'b10000001;
													assign node6314 = (inp[12]) ? 8'b10000100 : 8'b10010001;
											assign node6317 = (inp[12]) ? node6321 : node6318;
												assign node6318 = (inp[6]) ? 8'b10010101 : 8'b10000101;
												assign node6321 = (inp[6]) ? 8'b10100000 : 8'b10010101;
							assign node6324 = (inp[8]) ? node6444 : node6325;
								assign node6325 = (inp[10]) ? node6375 : node6326;
									assign node6326 = (inp[6]) ? node6360 : node6327;
										assign node6327 = (inp[11]) ? node6331 : node6328;
											assign node6328 = (inp[3]) ? 8'b00011110 : 8'b00011111;
											assign node6331 = (inp[12]) ? node6345 : node6332;
												assign node6332 = (inp[1]) ? node6340 : node6333;
													assign node6333 = (inp[3]) ? node6337 : node6334;
														assign node6334 = (inp[2]) ? 8'b00001110 : 8'b00001111;
														assign node6337 = (inp[2]) ? 8'b00001011 : 8'b00001110;
													assign node6340 = (inp[3]) ? 8'b00001011 : node6341;
														assign node6341 = (inp[2]) ? 8'b00001010 : 8'b00001011;
												assign node6345 = (inp[1]) ? node6353 : node6346;
													assign node6346 = (inp[2]) ? node6350 : node6347;
														assign node6347 = (inp[3]) ? 8'b00011110 : 8'b00011111;
														assign node6350 = (inp[3]) ? 8'b00011011 : 8'b00011110;
													assign node6353 = (inp[3]) ? node6357 : node6354;
														assign node6354 = (inp[2]) ? 8'b00011010 : 8'b00011011;
														assign node6357 = (inp[2]) ? 8'b00011011 : 8'b00011110;
										assign node6360 = (inp[11]) ? node6364 : node6361;
											assign node6361 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node6364 = (inp[12]) ? node6370 : node6365;
												assign node6365 = (inp[3]) ? 8'b00011011 : node6366;
													assign node6366 = (inp[1]) ? 8'b00011010 : 8'b00011110;
												assign node6370 = (inp[3]) ? 8'b00001110 : node6371;
													assign node6371 = (inp[1]) ? 8'b00001011 : 8'b00001111;
									assign node6375 = (inp[11]) ? node6393 : node6376;
										assign node6376 = (inp[6]) ? node6386 : node6377;
											assign node6377 = (inp[2]) ? node6383 : node6378;
												assign node6378 = (inp[3]) ? 8'b00011010 : node6379;
													assign node6379 = (inp[1]) ? 8'b10011001 : 8'b00011011;
												assign node6383 = (inp[3]) ? 8'b10010000 : 8'b10010001;
											assign node6386 = (inp[3]) ? node6390 : node6387;
												assign node6387 = (inp[1]) ? 8'b10000001 : 8'b00001011;
												assign node6390 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node6393 = (inp[1]) ? node6413 : node6394;
											assign node6394 = (inp[3]) ? node6406 : node6395;
												assign node6395 = (inp[2]) ? node6401 : node6396;
													assign node6396 = (inp[6]) ? node6398 : 8'b00001011;
														assign node6398 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node6401 = (inp[12]) ? 8'b00011010 : node6402;
														assign node6402 = (inp[6]) ? 8'b00011010 : 8'b00001010;
												assign node6406 = (inp[12]) ? node6410 : node6407;
													assign node6407 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node6410 = (inp[6]) ? 8'b00000010 : 8'b11110101;
											assign node6413 = (inp[3]) ? node6429 : node6414;
												assign node6414 = (inp[2]) ? node6422 : node6415;
													assign node6415 = (inp[6]) ? node6419 : node6416;
														assign node6416 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node6419 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node6422 = (inp[12]) ? node6426 : node6423;
														assign node6423 = (inp[6]) ? 8'b10110100 : 8'b10100100;
														assign node6426 = (inp[6]) ? 8'b10100101 : 8'b10110100;
												assign node6429 = (inp[2]) ? node6437 : node6430;
													assign node6430 = (inp[6]) ? node6434 : node6431;
														assign node6431 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node6434 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node6437 = (inp[6]) ? node6441 : node6438;
														assign node6438 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node6441 = (inp[12]) ? 8'b00000010 : 8'b11110111;
								assign node6444 = (inp[10]) ? node6518 : node6445;
									assign node6445 = (inp[11]) ? node6459 : node6446;
										assign node6446 = (inp[3]) ? node6454 : node6447;
											assign node6447 = (inp[6]) ? node6451 : node6448;
												assign node6448 = (inp[1]) ? 8'b10010101 : 8'b10011101;
												assign node6451 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node6454 = (inp[6]) ? 8'b10000100 : node6455;
												assign node6455 = (inp[2]) ? 8'b10010100 : 8'b10011100;
										assign node6459 = (inp[1]) ? node6489 : node6460;
											assign node6460 = (inp[3]) ? node6474 : node6461;
												assign node6461 = (inp[2]) ? node6469 : node6462;
													assign node6462 = (inp[12]) ? node6466 : node6463;
														assign node6463 = (inp[6]) ? 8'b10111100 : 8'b10101101;
														assign node6466 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node6469 = (inp[6]) ? node6471 : 8'b10111100;
														assign node6471 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node6474 = (inp[2]) ? node6482 : node6475;
													assign node6475 = (inp[6]) ? node6479 : node6476;
														assign node6476 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node6479 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node6482 = (inp[12]) ? node6486 : node6483;
														assign node6483 = (inp[6]) ? 8'b10110001 : 8'b10100001;
														assign node6486 = (inp[6]) ? 8'b10100100 : 8'b10110001;
											assign node6489 = (inp[3]) ? node6505 : node6490;
												assign node6490 = (inp[2]) ? node6498 : node6491;
													assign node6491 = (inp[6]) ? node6495 : node6492;
														assign node6492 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node6495 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node6498 = (inp[12]) ? node6502 : node6499;
														assign node6499 = (inp[6]) ? 8'b10110000 : 8'b10100000;
														assign node6502 = (inp[6]) ? 8'b10100001 : 8'b10110000;
												assign node6505 = (inp[2]) ? node6513 : node6506;
													assign node6506 = (inp[6]) ? node6510 : node6507;
														assign node6507 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node6510 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node6513 = (inp[12]) ? node6515 : 8'b10110001;
														assign node6515 = (inp[6]) ? 8'b10100100 : 8'b10110001;
									assign node6518 = (inp[1]) ? node6554 : node6519;
										assign node6519 = (inp[3]) ? node6539 : node6520;
											assign node6520 = (inp[11]) ? node6524 : node6521;
												assign node6521 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node6524 = (inp[2]) ? node6532 : node6525;
													assign node6525 = (inp[12]) ? node6529 : node6526;
														assign node6526 = (inp[6]) ? 8'b00011010 : 8'b00001011;
														assign node6529 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node6532 = (inp[6]) ? node6536 : node6533;
														assign node6533 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node6536 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node6539 = (inp[11]) ? node6547 : node6540;
												assign node6540 = (inp[6]) ? node6544 : node6541;
													assign node6541 = (inp[2]) ? 8'b10010000 : 8'b00011010;
													assign node6544 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node6547 = (inp[12]) ? node6551 : node6548;
													assign node6548 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node6551 = (inp[6]) ? 8'b00000010 : 8'b00011010;
										assign node6554 = (inp[3]) ? node6576 : node6555;
											assign node6555 = (inp[11]) ? node6561 : node6556;
												assign node6556 = (inp[6]) ? 8'b10000001 : node6557;
													assign node6557 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node6561 = (inp[2]) ? node6569 : node6562;
													assign node6562 = (inp[6]) ? node6566 : node6563;
														assign node6563 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node6566 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node6569 = (inp[6]) ? node6573 : node6570;
														assign node6570 = (inp[12]) ? 8'b10110100 : 8'b10100100;
														assign node6573 = (inp[12]) ? 8'b10100101 : 8'b10110100;
											assign node6576 = (inp[2]) ? node6588 : node6577;
												assign node6577 = (inp[6]) ? node6583 : node6578;
													assign node6578 = (inp[12]) ? 8'b00011010 : node6579;
														assign node6579 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node6583 = (inp[12]) ? 8'b00000010 : node6584;
														assign node6584 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node6588 = (inp[11]) ? node6594 : node6589;
													assign node6589 = (inp[6]) ? node6591 : 8'b10010000;
														assign node6591 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node6594 = (inp[6]) ? node6598 : node6595;
														assign node6595 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node6598 = (inp[12]) ? 8'b00000010 : 8'b11110111;
					assign node6601 = (inp[11]) ? node6975 : node6602;
						assign node6602 = (inp[0]) ? node6902 : node6603;
							assign node6603 = (inp[9]) ? node6743 : node6604;
								assign node6604 = (inp[10]) ? node6672 : node6605;
									assign node6605 = (inp[8]) ? node6637 : node6606;
										assign node6606 = (inp[3]) ? node6618 : node6607;
											assign node6607 = (inp[1]) ? node6615 : node6608;
												assign node6608 = (inp[6]) ? node6612 : node6609;
													assign node6609 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node6612 = (inp[2]) ? 8'b00011111 : 8'b00001111;
												assign node6615 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node6618 = (inp[1]) ? node6632 : node6619;
												assign node6619 = (inp[12]) ? node6625 : node6620;
													assign node6620 = (inp[2]) ? node6622 : 8'b00011110;
														assign node6622 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node6625 = (inp[6]) ? node6629 : node6626;
														assign node6626 = (inp[2]) ? 8'b00001110 : 8'b00011110;
														assign node6629 = (inp[2]) ? 8'b00011110 : 8'b00001110;
												assign node6632 = (inp[2]) ? node6634 : 8'b00011111;
													assign node6634 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node6637 = (inp[3]) ? node6655 : node6638;
											assign node6638 = (inp[1]) ? node6646 : node6639;
												assign node6639 = (inp[2]) ? node6643 : node6640;
													assign node6640 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node6643 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node6646 = (inp[12]) ? node6648 : 8'b10000010;
													assign node6648 = (inp[2]) ? node6652 : node6649;
														assign node6649 = (inp[6]) ? 8'b00000010 : 8'b00011010;
														assign node6652 = (inp[6]) ? 8'b10010000 : 8'b00000010;
											assign node6655 = (inp[1]) ? node6665 : node6656;
												assign node6656 = (inp[2]) ? node6662 : node6657;
													assign node6657 = (inp[6]) ? node6659 : 8'b00011010;
														assign node6659 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node6662 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node6665 = (inp[2]) ? node6669 : node6666;
													assign node6666 = (inp[6]) ? 8'b10000001 : 8'b10011001;
													assign node6669 = (inp[6]) ? 8'b10010001 : 8'b10000001;
									assign node6672 = (inp[8]) ? node6710 : node6673;
										assign node6673 = (inp[1]) ? node6693 : node6674;
											assign node6674 = (inp[3]) ? node6682 : node6675;
												assign node6675 = (inp[2]) ? node6679 : node6676;
													assign node6676 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node6679 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node6682 = (inp[2]) ? node6688 : node6683;
													assign node6683 = (inp[6]) ? node6685 : 8'b00011010;
														assign node6685 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node6688 = (inp[6]) ? 8'b10010000 : node6689;
														assign node6689 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node6693 = (inp[3]) ? node6703 : node6694;
												assign node6694 = (inp[6]) ? node6700 : node6695;
													assign node6695 = (inp[2]) ? node6697 : 8'b00011010;
														assign node6697 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node6700 = (inp[2]) ? 8'b10010000 : 8'b10000010;
												assign node6703 = (inp[6]) ? node6707 : node6704;
													assign node6704 = (inp[2]) ? 8'b10000001 : 8'b10011001;
													assign node6707 = (inp[2]) ? 8'b10010001 : 8'b10000001;
										assign node6710 = (inp[1]) ? node6726 : node6711;
											assign node6711 = (inp[3]) ? node6719 : node6712;
												assign node6712 = (inp[6]) ? node6716 : node6713;
													assign node6713 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node6716 = (inp[2]) ? 8'b10011101 : 8'b10001101;
												assign node6719 = (inp[6]) ? node6723 : node6720;
													assign node6720 = (inp[2]) ? 8'b10000100 : 8'b10011100;
													assign node6723 = (inp[2]) ? 8'b10010100 : 8'b10000100;
											assign node6726 = (inp[3]) ? node6734 : node6727;
												assign node6727 = (inp[2]) ? node6731 : node6728;
													assign node6728 = (inp[6]) ? 8'b10000100 : 8'b10011100;
													assign node6731 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node6734 = (inp[12]) ? 8'b10000101 : node6735;
													assign node6735 = (inp[6]) ? node6739 : node6736;
														assign node6736 = (inp[2]) ? 8'b10000101 : 8'b10011101;
														assign node6739 = (inp[2]) ? 8'b10010101 : 8'b10000101;
								assign node6743 = (inp[1]) ? node6831 : node6744;
									assign node6744 = (inp[3]) ? node6800 : node6745;
										assign node6745 = (inp[12]) ? node6771 : node6746;
											assign node6746 = (inp[6]) ? node6756 : node6747;
												assign node6747 = (inp[2]) ? node6749 : 8'b11111101;
													assign node6749 = (inp[8]) ? node6753 : node6750;
														assign node6750 = (inp[10]) ? 8'b10101001 : 8'b10101101;
														assign node6753 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node6756 = (inp[2]) ? node6764 : node6757;
													assign node6757 = (inp[8]) ? node6761 : node6758;
														assign node6758 = (inp[10]) ? 8'b10101001 : 8'b10101101;
														assign node6761 = (inp[10]) ? 8'b10101101 : 8'b10101001;
													assign node6764 = (inp[10]) ? node6768 : node6765;
														assign node6765 = (inp[8]) ? 8'b10111001 : 8'b11111101;
														assign node6768 = (inp[8]) ? 8'b11111101 : 8'b10111001;
											assign node6771 = (inp[10]) ? node6785 : node6772;
												assign node6772 = (inp[8]) ? node6778 : node6773;
													assign node6773 = (inp[2]) ? 8'b11111101 : node6774;
														assign node6774 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node6778 = (inp[6]) ? node6782 : node6779;
														assign node6779 = (inp[2]) ? 8'b10101001 : 8'b10111001;
														assign node6782 = (inp[2]) ? 8'b10111001 : 8'b10101001;
												assign node6785 = (inp[8]) ? node6793 : node6786;
													assign node6786 = (inp[2]) ? node6790 : node6787;
														assign node6787 = (inp[6]) ? 8'b10101001 : 8'b10111001;
														assign node6790 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node6793 = (inp[6]) ? node6797 : node6794;
														assign node6794 = (inp[2]) ? 8'b10101101 : 8'b11111101;
														assign node6797 = (inp[2]) ? 8'b11111101 : 8'b10101101;
										assign node6800 = (inp[10]) ? node6816 : node6801;
											assign node6801 = (inp[8]) ? node6809 : node6802;
												assign node6802 = (inp[2]) ? node6806 : node6803;
													assign node6803 = (inp[6]) ? 8'b10101100 : 8'b10111100;
													assign node6806 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node6809 = (inp[6]) ? node6813 : node6810;
													assign node6810 = (inp[2]) ? 8'b10100000 : 8'b10111000;
													assign node6813 = (inp[2]) ? 8'b10110000 : 8'b10100000;
											assign node6816 = (inp[8]) ? node6824 : node6817;
												assign node6817 = (inp[6]) ? node6821 : node6818;
													assign node6818 = (inp[2]) ? 8'b10100000 : 8'b10111000;
													assign node6821 = (inp[2]) ? 8'b10110000 : 8'b10100000;
												assign node6824 = (inp[6]) ? node6828 : node6825;
													assign node6825 = (inp[2]) ? 8'b10100100 : 8'b10111100;
													assign node6828 = (inp[2]) ? 8'b10110100 : 8'b10100100;
									assign node6831 = (inp[3]) ? node6865 : node6832;
										assign node6832 = (inp[6]) ? node6848 : node6833;
											assign node6833 = (inp[2]) ? node6841 : node6834;
												assign node6834 = (inp[8]) ? node6838 : node6835;
													assign node6835 = (inp[10]) ? 8'b10111000 : 8'b10111100;
													assign node6838 = (inp[10]) ? 8'b10111100 : 8'b10111000;
												assign node6841 = (inp[10]) ? node6845 : node6842;
													assign node6842 = (inp[8]) ? 8'b10100000 : 8'b10101100;
													assign node6845 = (inp[8]) ? 8'b10100100 : 8'b10100000;
											assign node6848 = (inp[2]) ? node6858 : node6849;
												assign node6849 = (inp[12]) ? node6851 : 8'b10100000;
													assign node6851 = (inp[8]) ? node6855 : node6852;
														assign node6852 = (inp[10]) ? 8'b10100000 : 8'b10101100;
														assign node6855 = (inp[10]) ? 8'b10100100 : 8'b10100000;
												assign node6858 = (inp[8]) ? node6862 : node6859;
													assign node6859 = (inp[10]) ? 8'b10110000 : 8'b10111100;
													assign node6862 = (inp[10]) ? 8'b10110100 : 8'b10110000;
										assign node6865 = (inp[6]) ? node6887 : node6866;
											assign node6866 = (inp[2]) ? node6880 : node6867;
												assign node6867 = (inp[12]) ? node6873 : node6868;
													assign node6868 = (inp[8]) ? 8'b10111001 : node6869;
														assign node6869 = (inp[10]) ? 8'b10111001 : 8'b11111101;
													assign node6873 = (inp[8]) ? node6877 : node6874;
														assign node6874 = (inp[10]) ? 8'b10111001 : 8'b11111101;
														assign node6877 = (inp[10]) ? 8'b11111101 : 8'b10111001;
												assign node6880 = (inp[10]) ? node6884 : node6881;
													assign node6881 = (inp[8]) ? 8'b10100001 : 8'b10101101;
													assign node6884 = (inp[8]) ? 8'b10100101 : 8'b10100001;
											assign node6887 = (inp[2]) ? node6895 : node6888;
												assign node6888 = (inp[10]) ? node6892 : node6889;
													assign node6889 = (inp[8]) ? 8'b10100001 : 8'b10101101;
													assign node6892 = (inp[8]) ? 8'b10100101 : 8'b10100001;
												assign node6895 = (inp[8]) ? node6899 : node6896;
													assign node6896 = (inp[10]) ? 8'b10110001 : 8'b11111101;
													assign node6899 = (inp[10]) ? 8'b11110101 : 8'b10110001;
							assign node6902 = (inp[6]) ? node6932 : node6903;
								assign node6903 = (inp[8]) ? node6921 : node6904;
									assign node6904 = (inp[10]) ? node6910 : node6905;
										assign node6905 = (inp[1]) ? 8'b11111101 : node6906;
											assign node6906 = (inp[3]) ? 8'b10111100 : 8'b11111101;
										assign node6910 = (inp[2]) ? node6916 : node6911;
											assign node6911 = (inp[3]) ? node6913 : 8'b10111001;
												assign node6913 = (inp[1]) ? 8'b10111001 : 8'b10111000;
											assign node6916 = (inp[1]) ? 8'b10110001 : node6917;
												assign node6917 = (inp[3]) ? 8'b10110000 : 8'b10111001;
									assign node6921 = (inp[2]) ? node6927 : node6922;
										assign node6922 = (inp[3]) ? node6924 : 8'b11111101;
											assign node6924 = (inp[1]) ? 8'b11111101 : 8'b10111100;
										assign node6927 = (inp[1]) ? 8'b11110101 : node6928;
											assign node6928 = (inp[3]) ? 8'b10110100 : 8'b11111101;
								assign node6932 = (inp[2]) ? node6950 : node6933;
									assign node6933 = (inp[1]) ? node6945 : node6934;
										assign node6934 = (inp[3]) ? node6940 : node6935;
											assign node6935 = (inp[8]) ? 8'b10101101 : node6936;
												assign node6936 = (inp[10]) ? 8'b10101001 : 8'b10101101;
											assign node6940 = (inp[8]) ? 8'b10100100 : node6941;
												assign node6941 = (inp[10]) ? 8'b10100000 : 8'b10101100;
										assign node6945 = (inp[8]) ? 8'b10100101 : node6946;
											assign node6946 = (inp[10]) ? 8'b10100001 : 8'b10101101;
									assign node6950 = (inp[10]) ? node6964 : node6951;
										assign node6951 = (inp[3]) ? node6957 : node6952;
											assign node6952 = (inp[1]) ? node6954 : 8'b11111101;
												assign node6954 = (inp[8]) ? 8'b11110101 : 8'b11111101;
											assign node6957 = (inp[1]) ? node6961 : node6958;
												assign node6958 = (inp[8]) ? 8'b10110100 : 8'b10111100;
												assign node6961 = (inp[8]) ? 8'b11110101 : 8'b11111101;
										assign node6964 = (inp[8]) ? node6970 : node6965;
											assign node6965 = (inp[1]) ? 8'b10110001 : node6966;
												assign node6966 = (inp[3]) ? 8'b10110000 : 8'b10111001;
											assign node6970 = (inp[1]) ? 8'b11110101 : node6971;
												assign node6971 = (inp[3]) ? 8'b10110100 : 8'b11111101;
						assign node6975 = (inp[8]) ? node7259 : node6976;
							assign node6976 = (inp[10]) ? node7116 : node6977;
								assign node6977 = (inp[0]) ? node7081 : node6978;
									assign node6978 = (inp[9]) ? node7030 : node6979;
										assign node6979 = (inp[3]) ? node7005 : node6980;
											assign node6980 = (inp[1]) ? node6990 : node6981;
												assign node6981 = (inp[2]) ? node6985 : node6982;
													assign node6982 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node6985 = (inp[6]) ? node6987 : 8'b00011110;
														assign node6987 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node6990 = (inp[6]) ? node6998 : node6991;
													assign node6991 = (inp[12]) ? node6995 : node6992;
														assign node6992 = (inp[2]) ? 8'b00011011 : 8'b00001110;
														assign node6995 = (inp[2]) ? 8'b00001110 : 8'b00011110;
													assign node6998 = (inp[12]) ? node7002 : node6999;
														assign node6999 = (inp[2]) ? 8'b00001011 : 8'b00011011;
														assign node7002 = (inp[2]) ? 8'b00011011 : 8'b00001110;
											assign node7005 = (inp[1]) ? node7017 : node7006;
												assign node7006 = (inp[2]) ? node7012 : node7007;
													assign node7007 = (inp[6]) ? node7009 : 8'b00001110;
														assign node7009 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node7012 = (inp[6]) ? node7014 : 8'b00011011;
														assign node7014 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node7017 = (inp[12]) ? node7025 : node7018;
													assign node7018 = (inp[2]) ? node7022 : node7019;
														assign node7019 = (inp[6]) ? 8'b00011010 : 8'b00001011;
														assign node7022 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node7025 = (inp[6]) ? 8'b00001011 : node7026;
														assign node7026 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node7030 = (inp[1]) ? node7056 : node7031;
											assign node7031 = (inp[3]) ? node7045 : node7032;
												assign node7032 = (inp[6]) ? node7040 : node7033;
													assign node7033 = (inp[2]) ? node7037 : node7034;
														assign node7034 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node7037 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node7040 = (inp[2]) ? node7042 : 8'b10111100;
														assign node7042 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node7045 = (inp[12]) ? node7051 : node7046;
													assign node7046 = (inp[6]) ? node7048 : 8'b10111001;
														assign node7048 = (inp[2]) ? 8'b10101001 : 8'b10111001;
													assign node7051 = (inp[6]) ? 8'b10101100 : node7052;
														assign node7052 = (inp[2]) ? 8'b10101100 : 8'b10111100;
											assign node7056 = (inp[6]) ? node7070 : node7057;
												assign node7057 = (inp[3]) ? node7063 : node7058;
													assign node7058 = (inp[2]) ? node7060 : 8'b10101100;
														assign node7060 = (inp[12]) ? 8'b10101100 : 8'b10111001;
													assign node7063 = (inp[2]) ? node7067 : node7064;
														assign node7064 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node7067 = (inp[12]) ? 8'b10101001 : 8'b10111000;
												assign node7070 = (inp[3]) ? node7076 : node7071;
													assign node7071 = (inp[12]) ? 8'b10111001 : node7072;
														assign node7072 = (inp[2]) ? 8'b10101001 : 8'b10111001;
													assign node7076 = (inp[2]) ? 8'b10111000 : node7077;
														assign node7077 = (inp[12]) ? 8'b10101001 : 8'b10111000;
									assign node7081 = (inp[1]) ? node7105 : node7082;
										assign node7082 = (inp[3]) ? node7094 : node7083;
											assign node7083 = (inp[2]) ? node7091 : node7084;
												assign node7084 = (inp[6]) ? node7088 : node7085;
													assign node7085 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node7088 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node7091 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node7094 = (inp[2]) ? node7102 : node7095;
												assign node7095 = (inp[12]) ? node7099 : node7096;
													assign node7096 = (inp[6]) ? 8'b10111001 : 8'b10101100;
													assign node7099 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node7102 = (inp[12]) ? 8'b10111001 : 8'b10101001;
										assign node7105 = (inp[2]) ? node7113 : node7106;
											assign node7106 = (inp[6]) ? node7110 : node7107;
												assign node7107 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node7110 = (inp[12]) ? 8'b10101001 : 8'b10111000;
											assign node7113 = (inp[12]) ? 8'b10111000 : 8'b10101000;
								assign node7116 = (inp[1]) ? node7192 : node7117;
									assign node7117 = (inp[3]) ? node7155 : node7118;
										assign node7118 = (inp[9]) ? node7138 : node7119;
											assign node7119 = (inp[0]) ? node7129 : node7120;
												assign node7120 = (inp[12]) ? node7122 : 8'b00001010;
													assign node7122 = (inp[2]) ? node7126 : node7123;
														assign node7123 = (inp[6]) ? 8'b00001011 : 8'b00011011;
														assign node7126 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node7129 = (inp[12]) ? 8'b10111000 : node7130;
													assign node7130 = (inp[6]) ? node7134 : node7131;
														assign node7131 = (inp[2]) ? 8'b10101000 : 8'b10101001;
														assign node7134 = (inp[2]) ? 8'b10101000 : 8'b10111000;
											assign node7138 = (inp[2]) ? node7146 : node7139;
												assign node7139 = (inp[12]) ? node7143 : node7140;
													assign node7140 = (inp[6]) ? 8'b10111000 : 8'b10101001;
													assign node7143 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node7146 = (inp[0]) ? node7152 : node7147;
													assign node7147 = (inp[12]) ? node7149 : 8'b10111000;
														assign node7149 = (inp[6]) ? 8'b10111000 : 8'b10101001;
													assign node7152 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node7155 = (inp[2]) ? node7175 : node7156;
											assign node7156 = (inp[6]) ? node7164 : node7157;
												assign node7157 = (inp[9]) ? node7161 : node7158;
													assign node7158 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node7161 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node7164 = (inp[12]) ? node7170 : node7165;
													assign node7165 = (inp[0]) ? 8'b10010101 : node7166;
														assign node7166 = (inp[9]) ? 8'b10010101 : 8'b11110111;
													assign node7170 = (inp[9]) ? 8'b10100000 : node7171;
														assign node7171 = (inp[0]) ? 8'b10100000 : 8'b00000010;
											assign node7175 = (inp[0]) ? node7189 : node7176;
												assign node7176 = (inp[12]) ? node7184 : node7177;
													assign node7177 = (inp[9]) ? node7181 : node7178;
														assign node7178 = (inp[6]) ? 8'b10100101 : 8'b11110111;
														assign node7181 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node7184 = (inp[6]) ? 8'b11110101 : node7185;
														assign node7185 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node7189 = (inp[12]) ? 8'b10010101 : 8'b10000101;
									assign node7192 = (inp[2]) ? node7230 : node7193;
										assign node7193 = (inp[6]) ? node7211 : node7194;
											assign node7194 = (inp[12]) ? node7204 : node7195;
												assign node7195 = (inp[0]) ? 8'b10001101 : node7196;
													assign node7196 = (inp[3]) ? node7200 : node7197;
														assign node7197 = (inp[9]) ? 8'b10101000 : 8'b00001010;
														assign node7200 = (inp[9]) ? 8'b10001101 : 8'b10101101;
												assign node7204 = (inp[0]) ? 8'b10011101 : node7205;
													assign node7205 = (inp[3]) ? node7207 : 8'b00011010;
														assign node7207 = (inp[9]) ? 8'b10011101 : 8'b11111101;
											assign node7211 = (inp[12]) ? node7221 : node7212;
												assign node7212 = (inp[0]) ? 8'b10010100 : node7213;
													assign node7213 = (inp[9]) ? node7217 : node7214;
														assign node7214 = (inp[3]) ? 8'b10110100 : 8'b11110111;
														assign node7217 = (inp[3]) ? 8'b10010100 : 8'b10010101;
												assign node7221 = (inp[0]) ? 8'b10000101 : node7222;
													assign node7222 = (inp[3]) ? node7226 : node7223;
														assign node7223 = (inp[9]) ? 8'b10100000 : 8'b00000010;
														assign node7226 = (inp[9]) ? 8'b10000101 : 8'b10100101;
										assign node7230 = (inp[0]) ? node7256 : node7231;
											assign node7231 = (inp[9]) ? node7245 : node7232;
												assign node7232 = (inp[3]) ? node7238 : node7233;
													assign node7233 = (inp[6]) ? node7235 : 8'b00000010;
														assign node7235 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node7238 = (inp[12]) ? node7242 : node7239;
														assign node7239 = (inp[6]) ? 8'b10100100 : 8'b10110100;
														assign node7242 = (inp[6]) ? 8'b10110100 : 8'b10100101;
												assign node7245 = (inp[12]) ? node7251 : node7246;
													assign node7246 = (inp[3]) ? 8'b10000100 : node7247;
														assign node7247 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node7251 = (inp[3]) ? node7253 : 8'b10100000;
														assign node7253 = (inp[6]) ? 8'b10010100 : 8'b10000101;
											assign node7256 = (inp[12]) ? 8'b10010100 : 8'b10000100;
							assign node7259 = (inp[1]) ? node7399 : node7260;
								assign node7260 = (inp[3]) ? node7332 : node7261;
									assign node7261 = (inp[0]) ? node7321 : node7262;
										assign node7262 = (inp[10]) ? node7290 : node7263;
											assign node7263 = (inp[9]) ? node7277 : node7264;
												assign node7264 = (inp[2]) ? node7272 : node7265;
													assign node7265 = (inp[12]) ? node7269 : node7266;
														assign node7266 = (inp[6]) ? 8'b00011010 : 8'b00001011;
														assign node7269 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node7272 = (inp[6]) ? node7274 : 8'b00011010;
														assign node7274 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node7277 = (inp[6]) ? node7285 : node7278;
													assign node7278 = (inp[2]) ? node7282 : node7279;
														assign node7279 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node7282 = (inp[12]) ? 8'b10101001 : 8'b10111000;
													assign node7285 = (inp[12]) ? 8'b10111000 : node7286;
														assign node7286 = (inp[2]) ? 8'b10101000 : 8'b10111000;
											assign node7290 = (inp[9]) ? node7306 : node7291;
												assign node7291 = (inp[12]) ? node7299 : node7292;
													assign node7292 = (inp[2]) ? node7296 : node7293;
														assign node7293 = (inp[6]) ? 8'b10111100 : 8'b10101101;
														assign node7296 = (inp[6]) ? 8'b10101100 : 8'b10111100;
													assign node7299 = (inp[6]) ? node7303 : node7300;
														assign node7300 = (inp[2]) ? 8'b10101101 : 8'b11111101;
														assign node7303 = (inp[2]) ? 8'b10111100 : 8'b10101101;
												assign node7306 = (inp[6]) ? node7314 : node7307;
													assign node7307 = (inp[12]) ? node7311 : node7308;
														assign node7308 = (inp[2]) ? 8'b10011100 : 8'b10001101;
														assign node7311 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node7314 = (inp[12]) ? node7318 : node7315;
														assign node7315 = (inp[2]) ? 8'b10001100 : 8'b10011100;
														assign node7318 = (inp[2]) ? 8'b10011100 : 8'b10001101;
										assign node7321 = (inp[2]) ? node7329 : node7322;
											assign node7322 = (inp[6]) ? node7326 : node7323;
												assign node7323 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node7326 = (inp[12]) ? 8'b10001101 : 8'b10011100;
											assign node7329 = (inp[12]) ? 8'b10011100 : 8'b10001100;
									assign node7332 = (inp[2]) ? node7364 : node7333;
										assign node7333 = (inp[6]) ? node7351 : node7334;
											assign node7334 = (inp[12]) ? node7344 : node7335;
												assign node7335 = (inp[0]) ? 8'b10001100 : node7336;
													assign node7336 = (inp[10]) ? node7340 : node7337;
														assign node7337 = (inp[9]) ? 8'b10101000 : 8'b00001010;
														assign node7340 = (inp[9]) ? 8'b10001100 : 8'b10101100;
												assign node7344 = (inp[0]) ? 8'b10011100 : node7345;
													assign node7345 = (inp[10]) ? node7347 : 8'b00011010;
														assign node7347 = (inp[9]) ? 8'b10011100 : 8'b10111100;
											assign node7351 = (inp[12]) ? node7357 : node7352;
												assign node7352 = (inp[10]) ? 8'b10010001 : node7353;
													assign node7353 = (inp[9]) ? 8'b10010101 : 8'b11110111;
												assign node7357 = (inp[0]) ? 8'b10000100 : node7358;
													assign node7358 = (inp[10]) ? node7360 : 8'b10100000;
														assign node7360 = (inp[9]) ? 8'b10000100 : 8'b10100100;
										assign node7364 = (inp[0]) ? node7396 : node7365;
											assign node7365 = (inp[9]) ? node7381 : node7366;
												assign node7366 = (inp[10]) ? node7374 : node7367;
													assign node7367 = (inp[6]) ? node7371 : node7368;
														assign node7368 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node7371 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node7374 = (inp[12]) ? node7378 : node7375;
														assign node7375 = (inp[6]) ? 8'b10100001 : 8'b10110001;
														assign node7378 = (inp[6]) ? 8'b10110001 : 8'b10100100;
												assign node7381 = (inp[10]) ? node7389 : node7382;
													assign node7382 = (inp[12]) ? node7386 : node7383;
														assign node7383 = (inp[6]) ? 8'b10000101 : 8'b10010101;
														assign node7386 = (inp[6]) ? 8'b10010101 : 8'b10100000;
													assign node7389 = (inp[12]) ? node7393 : node7390;
														assign node7390 = (inp[6]) ? 8'b10000001 : 8'b10010001;
														assign node7393 = (inp[6]) ? 8'b10010001 : 8'b10000100;
											assign node7396 = (inp[12]) ? 8'b10010001 : 8'b10000001;
								assign node7399 = (inp[0]) ? node7507 : node7400;
									assign node7400 = (inp[9]) ? node7454 : node7401;
										assign node7401 = (inp[10]) ? node7427 : node7402;
											assign node7402 = (inp[3]) ? node7414 : node7403;
												assign node7403 = (inp[6]) ? node7409 : node7404;
													assign node7404 = (inp[2]) ? 8'b00000010 : node7405;
														assign node7405 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node7409 = (inp[2]) ? 8'b11110101 : node7410;
														assign node7410 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node7414 = (inp[6]) ? node7420 : node7415;
													assign node7415 = (inp[2]) ? 8'b10100101 : node7416;
														assign node7416 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node7420 = (inp[2]) ? node7424 : node7421;
														assign node7421 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node7424 = (inp[12]) ? 8'b10110100 : 8'b10100100;
											assign node7427 = (inp[6]) ? node7441 : node7428;
												assign node7428 = (inp[2]) ? node7436 : node7429;
													assign node7429 = (inp[3]) ? node7433 : node7430;
														assign node7430 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node7433 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node7436 = (inp[12]) ? 8'b10100100 : node7437;
														assign node7437 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node7441 = (inp[3]) ? node7449 : node7442;
													assign node7442 = (inp[2]) ? node7446 : node7443;
														assign node7443 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node7446 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node7449 = (inp[2]) ? node7451 : 8'b10110000;
														assign node7451 = (inp[12]) ? 8'b10110000 : 8'b10100000;
										assign node7454 = (inp[6]) ? node7482 : node7455;
											assign node7455 = (inp[2]) ? node7469 : node7456;
												assign node7456 = (inp[3]) ? node7464 : node7457;
													assign node7457 = (inp[10]) ? node7461 : node7458;
														assign node7458 = (inp[12]) ? 8'b10111000 : 8'b10101000;
														assign node7461 = (inp[12]) ? 8'b10011100 : 8'b10001100;
													assign node7464 = (inp[10]) ? node7466 : 8'b10001101;
														assign node7466 = (inp[12]) ? 8'b10011001 : 8'b10001001;
												assign node7469 = (inp[12]) ? node7475 : node7470;
													assign node7470 = (inp[3]) ? 8'b10010100 : node7471;
														assign node7471 = (inp[10]) ? 8'b10010001 : 8'b10010101;
													assign node7475 = (inp[3]) ? node7479 : node7476;
														assign node7476 = (inp[10]) ? 8'b10000100 : 8'b10100000;
														assign node7479 = (inp[10]) ? 8'b10000001 : 8'b10000101;
											assign node7482 = (inp[10]) ? node7492 : node7483;
												assign node7483 = (inp[3]) ? 8'b10010100 : node7484;
													assign node7484 = (inp[2]) ? node7488 : node7485;
														assign node7485 = (inp[12]) ? 8'b10100000 : 8'b10010101;
														assign node7488 = (inp[12]) ? 8'b10010101 : 8'b10000101;
												assign node7492 = (inp[3]) ? node7500 : node7493;
													assign node7493 = (inp[2]) ? node7497 : node7494;
														assign node7494 = (inp[12]) ? 8'b10000100 : 8'b10010001;
														assign node7497 = (inp[12]) ? 8'b10010001 : 8'b10000001;
													assign node7500 = (inp[12]) ? node7504 : node7501;
														assign node7501 = (inp[2]) ? 8'b10000000 : 8'b10010000;
														assign node7504 = (inp[2]) ? 8'b10010000 : 8'b10000001;
									assign node7507 = (inp[2]) ? node7515 : node7508;
										assign node7508 = (inp[6]) ? node7512 : node7509;
											assign node7509 = (inp[12]) ? 8'b10011001 : 8'b10001001;
											assign node7512 = (inp[12]) ? 8'b10000001 : 8'b10010000;
										assign node7515 = (inp[12]) ? 8'b10010000 : 8'b10000000;
			assign node7518 = (inp[11]) ? node7938 : node7519;
				assign node7519 = (inp[0]) ? node7717 : node7520;
					assign node7520 = (inp[5]) ? node7524 : node7521;
						assign node7521 = (inp[12]) ? 8'b00000010 : 8'b10000010;
						assign node7524 = (inp[8]) ? node7600 : node7525;
							assign node7525 = (inp[3]) ? node7555 : node7526;
								assign node7526 = (inp[6]) ? node7538 : node7527;
									assign node7527 = (inp[12]) ? node7533 : node7528;
										assign node7528 = (inp[9]) ? node7530 : 8'b10000010;
											assign node7530 = (inp[13]) ? 8'b10100000 : 8'b10000010;
										assign node7533 = (inp[9]) ? node7535 : 8'b00000010;
											assign node7535 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node7538 = (inp[2]) ? node7550 : node7539;
										assign node7539 = (inp[12]) ? node7545 : node7540;
											assign node7540 = (inp[13]) ? node7542 : 8'b10000010;
												assign node7542 = (inp[9]) ? 8'b10100000 : 8'b10000010;
											assign node7545 = (inp[9]) ? node7547 : 8'b00000010;
												assign node7547 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node7550 = (inp[9]) ? node7552 : 8'b10010000;
											assign node7552 = (inp[13]) ? 8'b10110000 : 8'b10010000;
								assign node7555 = (inp[1]) ? node7583 : node7556;
									assign node7556 = (inp[9]) ? node7568 : node7557;
										assign node7557 = (inp[12]) ? node7563 : node7558;
											assign node7558 = (inp[2]) ? node7560 : 8'b10000010;
												assign node7560 = (inp[6]) ? 8'b10010000 : 8'b10000010;
											assign node7563 = (inp[2]) ? node7565 : 8'b00000010;
												assign node7565 = (inp[6]) ? 8'b10010000 : 8'b00000010;
										assign node7568 = (inp[13]) ? node7578 : node7569;
											assign node7569 = (inp[6]) ? node7573 : node7570;
												assign node7570 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7573 = (inp[2]) ? 8'b10010000 : node7574;
													assign node7574 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7578 = (inp[2]) ? node7580 : 8'b10100000;
												assign node7580 = (inp[6]) ? 8'b10110000 : 8'b10100000;
									assign node7583 = (inp[9]) ? node7589 : node7584;
										assign node7584 = (inp[2]) ? node7586 : 8'b10000001;
											assign node7586 = (inp[6]) ? 8'b10010001 : 8'b10000001;
										assign node7589 = (inp[13]) ? node7595 : node7590;
											assign node7590 = (inp[6]) ? node7592 : 8'b10000001;
												assign node7592 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node7595 = (inp[6]) ? node7597 : 8'b10100001;
												assign node7597 = (inp[2]) ? 8'b10110001 : 8'b10100001;
							assign node7600 = (inp[10]) ? node7668 : node7601;
								assign node7601 = (inp[2]) ? node7629 : node7602;
									assign node7602 = (inp[1]) ? node7614 : node7603;
										assign node7603 = (inp[12]) ? node7609 : node7604;
											assign node7604 = (inp[9]) ? node7606 : 8'b10000010;
												assign node7606 = (inp[13]) ? 8'b10100000 : 8'b10000010;
											assign node7609 = (inp[9]) ? node7611 : 8'b00000010;
												assign node7611 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node7614 = (inp[3]) ? node7624 : node7615;
											assign node7615 = (inp[9]) ? node7619 : node7616;
												assign node7616 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7619 = (inp[13]) ? 8'b10100000 : node7620;
													assign node7620 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7624 = (inp[13]) ? node7626 : 8'b10000001;
												assign node7626 = (inp[9]) ? 8'b10100001 : 8'b10000001;
									assign node7629 = (inp[6]) ? node7651 : node7630;
										assign node7630 = (inp[13]) ? node7638 : node7631;
											assign node7631 = (inp[12]) ? 8'b00000010 : node7632;
												assign node7632 = (inp[1]) ? node7634 : 8'b10000010;
													assign node7634 = (inp[3]) ? 8'b10000001 : 8'b10000010;
											assign node7638 = (inp[9]) ? node7648 : node7639;
												assign node7639 = (inp[1]) ? node7643 : node7640;
													assign node7640 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node7643 = (inp[3]) ? 8'b10000001 : node7644;
														assign node7644 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7648 = (inp[1]) ? 8'b10100001 : 8'b10100000;
										assign node7651 = (inp[3]) ? node7657 : node7652;
											assign node7652 = (inp[13]) ? node7654 : 8'b10010000;
												assign node7654 = (inp[9]) ? 8'b10110000 : 8'b10010000;
											assign node7657 = (inp[1]) ? node7663 : node7658;
												assign node7658 = (inp[9]) ? node7660 : 8'b10010000;
													assign node7660 = (inp[13]) ? 8'b10110000 : 8'b10010000;
												assign node7663 = (inp[9]) ? node7665 : 8'b10010001;
													assign node7665 = (inp[13]) ? 8'b10110001 : 8'b10010001;
								assign node7668 = (inp[9]) ? node7686 : node7669;
									assign node7669 = (inp[6]) ? node7675 : node7670;
										assign node7670 = (inp[3]) ? node7672 : 8'b10000100;
											assign node7672 = (inp[1]) ? 8'b10000101 : 8'b10000100;
										assign node7675 = (inp[2]) ? node7681 : node7676;
											assign node7676 = (inp[3]) ? node7678 : 8'b10000100;
												assign node7678 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node7681 = (inp[1]) ? node7683 : 8'b10010100;
												assign node7683 = (inp[3]) ? 8'b10010101 : 8'b10010100;
									assign node7686 = (inp[13]) ? node7700 : node7687;
										assign node7687 = (inp[3]) ? node7693 : node7688;
											assign node7688 = (inp[6]) ? node7690 : 8'b10000100;
												assign node7690 = (inp[2]) ? 8'b10010100 : 8'b10000100;
											assign node7693 = (inp[1]) ? node7695 : 8'b10000100;
												assign node7695 = (inp[6]) ? node7697 : 8'b10000101;
													assign node7697 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node7700 = (inp[2]) ? node7706 : node7701;
											assign node7701 = (inp[1]) ? node7703 : 8'b10100100;
												assign node7703 = (inp[3]) ? 8'b10100101 : 8'b10100100;
											assign node7706 = (inp[6]) ? node7712 : node7707;
												assign node7707 = (inp[3]) ? node7709 : 8'b10100100;
													assign node7709 = (inp[1]) ? 8'b10100101 : 8'b10100100;
												assign node7712 = (inp[1]) ? node7714 : 8'b10110100;
													assign node7714 = (inp[3]) ? 8'b11110101 : 8'b10110100;
					assign node7717 = (inp[2]) ? node7801 : node7718;
						assign node7718 = (inp[13]) ? node7750 : node7719;
							assign node7719 = (inp[1]) ? node7731 : node7720;
								assign node7720 = (inp[8]) ? node7724 : node7721;
									assign node7721 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7724 = (inp[10]) ? node7726 : 8'b10000100;
										assign node7726 = (inp[5]) ? 8'b10000100 : node7727;
											assign node7727 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node7731 = (inp[8]) ? node7739 : node7732;
									assign node7732 = (inp[5]) ? 8'b10000001 : node7733;
										assign node7733 = (inp[3]) ? node7735 : 8'b10000001;
											assign node7735 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7739 = (inp[5]) ? 8'b10000101 : node7740;
										assign node7740 = (inp[10]) ? node7744 : node7741;
											assign node7741 = (inp[3]) ? 8'b10000100 : 8'b10000101;
											assign node7744 = (inp[3]) ? node7746 : 8'b10000001;
												assign node7746 = (inp[12]) ? 8'b00000010 : 8'b10000010;
							assign node7750 = (inp[1]) ? node7770 : node7751;
								assign node7751 = (inp[8]) ? node7759 : node7752;
									assign node7752 = (inp[9]) ? node7754 : 8'b10100000;
										assign node7754 = (inp[5]) ? 8'b10100000 : node7755;
											assign node7755 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7759 = (inp[5]) ? 8'b10100100 : node7760;
										assign node7760 = (inp[10]) ? node7764 : node7761;
											assign node7761 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node7764 = (inp[9]) ? node7766 : 8'b10100000;
												assign node7766 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node7770 = (inp[5]) ? node7798 : node7771;
									assign node7771 = (inp[9]) ? node7783 : node7772;
										assign node7772 = (inp[3]) ? node7778 : node7773;
											assign node7773 = (inp[8]) ? node7775 : 8'b10100001;
												assign node7775 = (inp[10]) ? 8'b10100001 : 8'b10100101;
											assign node7778 = (inp[8]) ? node7780 : 8'b10100000;
												assign node7780 = (inp[10]) ? 8'b10100000 : 8'b10100100;
										assign node7783 = (inp[3]) ? node7789 : node7784;
											assign node7784 = (inp[8]) ? node7786 : 8'b10000001;
												assign node7786 = (inp[10]) ? 8'b10000001 : 8'b10000101;
											assign node7789 = (inp[8]) ? node7793 : node7790;
												assign node7790 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7793 = (inp[10]) ? node7795 : 8'b10000100;
													assign node7795 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7798 = (inp[8]) ? 8'b10100101 : 8'b10100001;
						assign node7801 = (inp[1]) ? node7853 : node7802;
							assign node7802 = (inp[8]) ? node7822 : node7803;
								assign node7803 = (inp[13]) ? node7811 : node7804;
									assign node7804 = (inp[5]) ? 8'b10010000 : node7805;
										assign node7805 = (inp[6]) ? node7807 : 8'b10010000;
											assign node7807 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7811 = (inp[5]) ? 8'b10110000 : node7812;
										assign node7812 = (inp[6]) ? node7816 : node7813;
											assign node7813 = (inp[9]) ? 8'b10010000 : 8'b10110000;
											assign node7816 = (inp[9]) ? node7818 : 8'b10100000;
												assign node7818 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node7822 = (inp[5]) ? node7850 : node7823;
									assign node7823 = (inp[6]) ? node7835 : node7824;
										assign node7824 = (inp[10]) ? node7830 : node7825;
											assign node7825 = (inp[9]) ? 8'b10010100 : node7826;
												assign node7826 = (inp[13]) ? 8'b10110100 : 8'b10010100;
											assign node7830 = (inp[13]) ? node7832 : 8'b10010000;
												assign node7832 = (inp[9]) ? 8'b10010000 : 8'b10110000;
										assign node7835 = (inp[10]) ? node7841 : node7836;
											assign node7836 = (inp[13]) ? node7838 : 8'b10000100;
												assign node7838 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node7841 = (inp[9]) ? node7847 : node7842;
												assign node7842 = (inp[13]) ? 8'b10100000 : node7843;
													assign node7843 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7847 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7850 = (inp[13]) ? 8'b10110100 : 8'b10010100;
							assign node7853 = (inp[5]) ? node7931 : node7854;
								assign node7854 = (inp[3]) ? node7890 : node7855;
									assign node7855 = (inp[6]) ? node7873 : node7856;
										assign node7856 = (inp[8]) ? node7862 : node7857;
											assign node7857 = (inp[9]) ? 8'b10010001 : node7858;
												assign node7858 = (inp[13]) ? 8'b10110001 : 8'b10010001;
											assign node7862 = (inp[10]) ? node7868 : node7863;
												assign node7863 = (inp[13]) ? node7865 : 8'b10010101;
													assign node7865 = (inp[9]) ? 8'b10010101 : 8'b11110101;
												assign node7868 = (inp[13]) ? node7870 : 8'b10010001;
													assign node7870 = (inp[9]) ? 8'b10010001 : 8'b10110001;
										assign node7873 = (inp[10]) ? node7885 : node7874;
											assign node7874 = (inp[8]) ? node7880 : node7875;
												assign node7875 = (inp[13]) ? node7877 : 8'b10000001;
													assign node7877 = (inp[9]) ? 8'b10000001 : 8'b10100001;
												assign node7880 = (inp[13]) ? node7882 : 8'b10000101;
													assign node7882 = (inp[9]) ? 8'b10000101 : 8'b10100101;
											assign node7885 = (inp[9]) ? 8'b10000001 : node7886;
												assign node7886 = (inp[13]) ? 8'b10100001 : 8'b10000001;
									assign node7890 = (inp[6]) ? node7906 : node7891;
										assign node7891 = (inp[13]) ? node7897 : node7892;
											assign node7892 = (inp[8]) ? node7894 : 8'b10010000;
												assign node7894 = (inp[10]) ? 8'b10010000 : 8'b10010100;
											assign node7897 = (inp[9]) ? node7903 : node7898;
												assign node7898 = (inp[8]) ? node7900 : 8'b10110000;
													assign node7900 = (inp[10]) ? 8'b10110000 : 8'b10110100;
												assign node7903 = (inp[10]) ? 8'b10010000 : 8'b10010100;
										assign node7906 = (inp[13]) ? node7918 : node7907;
											assign node7907 = (inp[12]) ? node7913 : node7908;
												assign node7908 = (inp[10]) ? 8'b10000010 : node7909;
													assign node7909 = (inp[8]) ? 8'b10000100 : 8'b10000010;
												assign node7913 = (inp[10]) ? 8'b00000010 : node7914;
													assign node7914 = (inp[8]) ? 8'b10000100 : 8'b00000010;
											assign node7918 = (inp[9]) ? node7924 : node7919;
												assign node7919 = (inp[10]) ? 8'b10100000 : node7920;
													assign node7920 = (inp[8]) ? 8'b10100100 : 8'b10100000;
												assign node7924 = (inp[10]) ? node7928 : node7925;
													assign node7925 = (inp[8]) ? 8'b10000100 : 8'b10000010;
													assign node7928 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node7931 = (inp[8]) ? node7935 : node7932;
									assign node7932 = (inp[13]) ? 8'b10110001 : 8'b10010001;
									assign node7935 = (inp[13]) ? 8'b11110101 : 8'b10010101;
				assign node7938 = (inp[12]) ? node8276 : node7939;
					assign node7939 = (inp[5]) ? node8101 : node7940;
						assign node7940 = (inp[0]) ? node7942 : 8'b11110111;
							assign node7942 = (inp[8]) ? node7996 : node7943;
								assign node7943 = (inp[1]) ? node7961 : node7944;
									assign node7944 = (inp[6]) ? node7956 : node7945;
										assign node7945 = (inp[2]) ? node7951 : node7946;
											assign node7946 = (inp[9]) ? 8'b11110111 : node7947;
												assign node7947 = (inp[13]) ? 8'b10010101 : 8'b11110111;
											assign node7951 = (inp[9]) ? 8'b10100101 : node7952;
												assign node7952 = (inp[13]) ? 8'b10000101 : 8'b10100101;
										assign node7956 = (inp[13]) ? node7958 : 8'b11110111;
											assign node7958 = (inp[9]) ? 8'b11110111 : 8'b10010101;
									assign node7961 = (inp[3]) ? node7979 : node7962;
										assign node7962 = (inp[2]) ? node7968 : node7963;
											assign node7963 = (inp[9]) ? 8'b10110100 : node7964;
												assign node7964 = (inp[13]) ? 8'b10010100 : 8'b10110100;
											assign node7968 = (inp[6]) ? node7974 : node7969;
												assign node7969 = (inp[13]) ? node7971 : 8'b10100100;
													assign node7971 = (inp[9]) ? 8'b10100100 : 8'b10000100;
												assign node7974 = (inp[13]) ? node7976 : 8'b10110100;
													assign node7976 = (inp[9]) ? 8'b10110100 : 8'b10010100;
										assign node7979 = (inp[9]) ? node7991 : node7980;
											assign node7980 = (inp[13]) ? node7986 : node7981;
												assign node7981 = (inp[6]) ? 8'b11110111 : node7982;
													assign node7982 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node7986 = (inp[2]) ? node7988 : 8'b10010101;
													assign node7988 = (inp[6]) ? 8'b10010101 : 8'b10000101;
											assign node7991 = (inp[6]) ? 8'b11110111 : node7992;
												assign node7992 = (inp[2]) ? 8'b10100101 : 8'b11110111;
								assign node7996 = (inp[10]) ? node8048 : node7997;
									assign node7997 = (inp[13]) ? node8015 : node7998;
										assign node7998 = (inp[6]) ? node8010 : node7999;
											assign node7999 = (inp[2]) ? node8005 : node8000;
												assign node8000 = (inp[1]) ? node8002 : 8'b10110001;
													assign node8002 = (inp[3]) ? 8'b10110001 : 8'b10110000;
												assign node8005 = (inp[3]) ? 8'b10100001 : node8006;
													assign node8006 = (inp[1]) ? 8'b10100000 : 8'b10100001;
											assign node8010 = (inp[3]) ? 8'b10110001 : node8011;
												assign node8011 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node8015 = (inp[9]) ? node8033 : node8016;
											assign node8016 = (inp[2]) ? node8022 : node8017;
												assign node8017 = (inp[1]) ? node8019 : 8'b10010001;
													assign node8019 = (inp[3]) ? 8'b10010001 : 8'b10010000;
												assign node8022 = (inp[6]) ? node8028 : node8023;
													assign node8023 = (inp[1]) ? node8025 : 8'b10000001;
														assign node8025 = (inp[3]) ? 8'b10000001 : 8'b10000000;
													assign node8028 = (inp[3]) ? 8'b10010001 : node8029;
														assign node8029 = (inp[1]) ? 8'b10010000 : 8'b10010001;
											assign node8033 = (inp[3]) ? node8043 : node8034;
												assign node8034 = (inp[1]) ? node8038 : node8035;
													assign node8035 = (inp[2]) ? 8'b10100001 : 8'b10110001;
													assign node8038 = (inp[2]) ? node8040 : 8'b10110000;
														assign node8040 = (inp[6]) ? 8'b10110000 : 8'b10100000;
												assign node8043 = (inp[2]) ? node8045 : 8'b10110001;
													assign node8045 = (inp[6]) ? 8'b10110001 : 8'b10100001;
									assign node8048 = (inp[9]) ? node8084 : node8049;
										assign node8049 = (inp[13]) ? node8067 : node8050;
											assign node8050 = (inp[1]) ? node8056 : node8051;
												assign node8051 = (inp[6]) ? 8'b11110111 : node8052;
													assign node8052 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node8056 = (inp[3]) ? node8062 : node8057;
													assign node8057 = (inp[2]) ? node8059 : 8'b10110100;
														assign node8059 = (inp[6]) ? 8'b10110100 : 8'b10100100;
													assign node8062 = (inp[2]) ? node8064 : 8'b11110111;
														assign node8064 = (inp[6]) ? 8'b11110111 : 8'b10100101;
											assign node8067 = (inp[6]) ? node8079 : node8068;
												assign node8068 = (inp[2]) ? node8074 : node8069;
													assign node8069 = (inp[1]) ? node8071 : 8'b10010101;
														assign node8071 = (inp[3]) ? 8'b10010101 : 8'b10010100;
													assign node8074 = (inp[3]) ? 8'b10000101 : node8075;
														assign node8075 = (inp[1]) ? 8'b10000100 : 8'b10000101;
												assign node8079 = (inp[1]) ? node8081 : 8'b10010101;
													assign node8081 = (inp[3]) ? 8'b10010101 : 8'b10010100;
										assign node8084 = (inp[2]) ? node8090 : node8085;
											assign node8085 = (inp[1]) ? node8087 : 8'b11110111;
												assign node8087 = (inp[3]) ? 8'b11110111 : 8'b10110100;
											assign node8090 = (inp[6]) ? node8096 : node8091;
												assign node8091 = (inp[1]) ? node8093 : 8'b10100101;
													assign node8093 = (inp[3]) ? 8'b10100101 : 8'b10100100;
												assign node8096 = (inp[1]) ? node8098 : 8'b11110111;
													assign node8098 = (inp[3]) ? 8'b11110111 : 8'b10110100;
						assign node8101 = (inp[13]) ? node8167 : node8102;
							assign node8102 = (inp[1]) ? node8128 : node8103;
								assign node8103 = (inp[2]) ? node8111 : node8104;
									assign node8104 = (inp[8]) ? node8106 : 8'b11110111;
										assign node8106 = (inp[0]) ? 8'b10110001 : node8107;
											assign node8107 = (inp[10]) ? 8'b10110001 : 8'b11110111;
									assign node8111 = (inp[6]) ? node8121 : node8112;
										assign node8112 = (inp[0]) ? node8118 : node8113;
											assign node8113 = (inp[8]) ? node8115 : 8'b11110111;
												assign node8115 = (inp[10]) ? 8'b10110001 : 8'b11110111;
											assign node8118 = (inp[8]) ? 8'b10100001 : 8'b10100101;
										assign node8121 = (inp[8]) ? node8123 : 8'b10100101;
											assign node8123 = (inp[0]) ? 8'b10100001 : node8124;
												assign node8124 = (inp[10]) ? 8'b10100001 : 8'b10100101;
								assign node8128 = (inp[8]) ? node8144 : node8129;
									assign node8129 = (inp[0]) ? node8141 : node8130;
										assign node8130 = (inp[3]) ? node8136 : node8131;
											assign node8131 = (inp[6]) ? node8133 : 8'b11110111;
												assign node8133 = (inp[2]) ? 8'b10100101 : 8'b11110111;
											assign node8136 = (inp[2]) ? node8138 : 8'b10110100;
												assign node8138 = (inp[6]) ? 8'b10100100 : 8'b10110100;
										assign node8141 = (inp[2]) ? 8'b10100100 : 8'b10110100;
									assign node8144 = (inp[0]) ? node8164 : node8145;
										assign node8145 = (inp[10]) ? node8153 : node8146;
											assign node8146 = (inp[3]) ? 8'b10110100 : node8147;
												assign node8147 = (inp[2]) ? node8149 : 8'b11110111;
													assign node8149 = (inp[6]) ? 8'b10100101 : 8'b11110111;
											assign node8153 = (inp[3]) ? node8159 : node8154;
												assign node8154 = (inp[6]) ? node8156 : 8'b10110001;
													assign node8156 = (inp[2]) ? 8'b10100001 : 8'b10110001;
												assign node8159 = (inp[2]) ? node8161 : 8'b10110000;
													assign node8161 = (inp[6]) ? 8'b10100000 : 8'b10110000;
										assign node8164 = (inp[2]) ? 8'b10100000 : 8'b10110000;
							assign node8167 = (inp[8]) ? node8213 : node8168;
								assign node8168 = (inp[2]) ? node8186 : node8169;
									assign node8169 = (inp[9]) ? node8179 : node8170;
										assign node8170 = (inp[0]) ? node8176 : node8171;
											assign node8171 = (inp[3]) ? node8173 : 8'b11110111;
												assign node8173 = (inp[1]) ? 8'b10110100 : 8'b11110111;
											assign node8176 = (inp[1]) ? 8'b10010100 : 8'b10010101;
										assign node8179 = (inp[1]) ? node8181 : 8'b10010101;
											assign node8181 = (inp[3]) ? 8'b10010100 : node8182;
												assign node8182 = (inp[0]) ? 8'b10010100 : 8'b10010101;
									assign node8186 = (inp[0]) ? node8210 : node8187;
										assign node8187 = (inp[9]) ? node8199 : node8188;
											assign node8188 = (inp[6]) ? node8194 : node8189;
												assign node8189 = (inp[3]) ? node8191 : 8'b11110111;
													assign node8191 = (inp[1]) ? 8'b10110100 : 8'b11110111;
												assign node8194 = (inp[3]) ? node8196 : 8'b10100101;
													assign node8196 = (inp[1]) ? 8'b10100100 : 8'b10100101;
											assign node8199 = (inp[6]) ? node8205 : node8200;
												assign node8200 = (inp[3]) ? node8202 : 8'b10010101;
													assign node8202 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node8205 = (inp[1]) ? node8207 : 8'b10000101;
													assign node8207 = (inp[3]) ? 8'b10000100 : 8'b10000101;
										assign node8210 = (inp[1]) ? 8'b10000100 : 8'b10000101;
								assign node8213 = (inp[1]) ? node8241 : node8214;
									assign node8214 = (inp[0]) ? node8238 : node8215;
										assign node8215 = (inp[10]) ? node8227 : node8216;
											assign node8216 = (inp[9]) ? node8222 : node8217;
												assign node8217 = (inp[6]) ? node8219 : 8'b11110111;
													assign node8219 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node8222 = (inp[6]) ? node8224 : 8'b10010101;
													assign node8224 = (inp[2]) ? 8'b10000101 : 8'b10010101;
											assign node8227 = (inp[9]) ? node8233 : node8228;
												assign node8228 = (inp[2]) ? node8230 : 8'b10110001;
													assign node8230 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node8233 = (inp[6]) ? node8235 : 8'b10010001;
													assign node8235 = (inp[2]) ? 8'b10000001 : 8'b10010001;
										assign node8238 = (inp[2]) ? 8'b10000001 : 8'b10010001;
									assign node8241 = (inp[0]) ? node8273 : node8242;
										assign node8242 = (inp[10]) ? node8260 : node8243;
											assign node8243 = (inp[3]) ? node8249 : node8244;
												assign node8244 = (inp[9]) ? node8246 : 8'b11110111;
													assign node8246 = (inp[6]) ? 8'b10000101 : 8'b10010101;
												assign node8249 = (inp[9]) ? node8255 : node8250;
													assign node8250 = (inp[6]) ? node8252 : 8'b10110100;
														assign node8252 = (inp[2]) ? 8'b10100100 : 8'b10110100;
													assign node8255 = (inp[2]) ? node8257 : 8'b10010100;
														assign node8257 = (inp[6]) ? 8'b10000100 : 8'b10010100;
											assign node8260 = (inp[3]) ? node8266 : node8261;
												assign node8261 = (inp[9]) ? 8'b10010001 : node8262;
													assign node8262 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node8266 = (inp[9]) ? node8268 : 8'b10110000;
													assign node8268 = (inp[2]) ? node8270 : 8'b10010000;
														assign node8270 = (inp[6]) ? 8'b10000000 : 8'b10010000;
										assign node8273 = (inp[2]) ? 8'b10000000 : 8'b10010000;
					assign node8276 = (inp[0]) ? node8434 : node8277;
						assign node8277 = (inp[5]) ? node8279 : 8'b00000010;
							assign node8279 = (inp[6]) ? node8333 : node8280;
								assign node8280 = (inp[1]) ? node8298 : node8281;
									assign node8281 = (inp[10]) ? node8287 : node8282;
										assign node8282 = (inp[13]) ? node8284 : 8'b00000010;
											assign node8284 = (inp[9]) ? 8'b10100000 : 8'b00000010;
										assign node8287 = (inp[8]) ? node8293 : node8288;
											assign node8288 = (inp[13]) ? node8290 : 8'b00000010;
												assign node8290 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node8293 = (inp[9]) ? node8295 : 8'b10100100;
												assign node8295 = (inp[13]) ? 8'b10000100 : 8'b10100100;
									assign node8298 = (inp[3]) ? node8316 : node8299;
										assign node8299 = (inp[13]) ? node8305 : node8300;
											assign node8300 = (inp[10]) ? node8302 : 8'b00000010;
												assign node8302 = (inp[8]) ? 8'b10100100 : 8'b00000010;
											assign node8305 = (inp[9]) ? node8311 : node8306;
												assign node8306 = (inp[10]) ? node8308 : 8'b00000010;
													assign node8308 = (inp[8]) ? 8'b10100100 : 8'b00000010;
												assign node8311 = (inp[8]) ? node8313 : 8'b10100000;
													assign node8313 = (inp[10]) ? 8'b10000100 : 8'b10100000;
										assign node8316 = (inp[10]) ? node8322 : node8317;
											assign node8317 = (inp[9]) ? node8319 : 8'b10100101;
												assign node8319 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node8322 = (inp[8]) ? node8328 : node8323;
												assign node8323 = (inp[9]) ? node8325 : 8'b10100101;
													assign node8325 = (inp[13]) ? 8'b10000101 : 8'b10100101;
												assign node8328 = (inp[13]) ? node8330 : 8'b10100001;
													assign node8330 = (inp[9]) ? 8'b10000001 : 8'b10100001;
								assign node8333 = (inp[2]) ? node8385 : node8334;
									assign node8334 = (inp[3]) ? node8352 : node8335;
										assign node8335 = (inp[10]) ? node8341 : node8336;
											assign node8336 = (inp[13]) ? node8338 : 8'b00000010;
												assign node8338 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node8341 = (inp[8]) ? node8347 : node8342;
												assign node8342 = (inp[13]) ? node8344 : 8'b00000010;
													assign node8344 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node8347 = (inp[13]) ? node8349 : 8'b10100100;
													assign node8349 = (inp[9]) ? 8'b10000100 : 8'b10100100;
										assign node8352 = (inp[1]) ? node8368 : node8353;
											assign node8353 = (inp[8]) ? node8359 : node8354;
												assign node8354 = (inp[13]) ? node8356 : 8'b00000010;
													assign node8356 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node8359 = (inp[10]) ? node8363 : node8360;
													assign node8360 = (inp[13]) ? 8'b10100000 : 8'b00000010;
													assign node8363 = (inp[13]) ? node8365 : 8'b10100100;
														assign node8365 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node8368 = (inp[13]) ? node8374 : node8369;
												assign node8369 = (inp[8]) ? node8371 : 8'b10100101;
													assign node8371 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node8374 = (inp[9]) ? node8380 : node8375;
													assign node8375 = (inp[8]) ? node8377 : 8'b10100101;
														assign node8377 = (inp[10]) ? 8'b10100001 : 8'b10100101;
													assign node8380 = (inp[8]) ? node8382 : 8'b10000101;
														assign node8382 = (inp[10]) ? 8'b10000001 : 8'b10000101;
									assign node8385 = (inp[13]) ? node8403 : node8386;
										assign node8386 = (inp[1]) ? node8392 : node8387;
											assign node8387 = (inp[10]) ? node8389 : 8'b11110101;
												assign node8389 = (inp[8]) ? 8'b10110001 : 8'b11110101;
											assign node8392 = (inp[3]) ? node8398 : node8393;
												assign node8393 = (inp[10]) ? node8395 : 8'b11110101;
													assign node8395 = (inp[8]) ? 8'b10110001 : 8'b11110101;
												assign node8398 = (inp[8]) ? node8400 : 8'b10110100;
													assign node8400 = (inp[10]) ? 8'b10110000 : 8'b10110100;
										assign node8403 = (inp[9]) ? node8421 : node8404;
											assign node8404 = (inp[8]) ? node8410 : node8405;
												assign node8405 = (inp[1]) ? node8407 : 8'b11110101;
													assign node8407 = (inp[3]) ? 8'b10110100 : 8'b11110101;
												assign node8410 = (inp[10]) ? node8416 : node8411;
													assign node8411 = (inp[3]) ? node8413 : 8'b11110101;
														assign node8413 = (inp[1]) ? 8'b10110100 : 8'b11110101;
													assign node8416 = (inp[3]) ? node8418 : 8'b10110001;
														assign node8418 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node8421 = (inp[3]) ? node8427 : node8422;
												assign node8422 = (inp[8]) ? node8424 : 8'b10010101;
													assign node8424 = (inp[10]) ? 8'b10010001 : 8'b10010101;
												assign node8427 = (inp[1]) ? node8429 : 8'b10010101;
													assign node8429 = (inp[10]) ? node8431 : 8'b10010100;
														assign node8431 = (inp[8]) ? 8'b10010000 : 8'b10010100;
						assign node8434 = (inp[2]) ? node8510 : node8435;
							assign node8435 = (inp[1]) ? node8461 : node8436;
								assign node8436 = (inp[8]) ? node8444 : node8437;
									assign node8437 = (inp[13]) ? node8439 : 8'b00000010;
										assign node8439 = (inp[9]) ? node8441 : 8'b10100000;
											assign node8441 = (inp[5]) ? 8'b10100000 : 8'b00000010;
									assign node8444 = (inp[10]) ? node8452 : node8445;
										assign node8445 = (inp[13]) ? node8447 : 8'b10100100;
											assign node8447 = (inp[9]) ? node8449 : 8'b10000100;
												assign node8449 = (inp[5]) ? 8'b10000100 : 8'b10100100;
										assign node8452 = (inp[5]) ? node8458 : node8453;
											assign node8453 = (inp[13]) ? node8455 : 8'b00000010;
												assign node8455 = (inp[9]) ? 8'b00000010 : 8'b10100000;
											assign node8458 = (inp[13]) ? 8'b10000100 : 8'b10100100;
								assign node8461 = (inp[3]) ? node8485 : node8462;
									assign node8462 = (inp[13]) ? node8470 : node8463;
										assign node8463 = (inp[8]) ? node8465 : 8'b10100101;
											assign node8465 = (inp[5]) ? 8'b10100001 : node8466;
												assign node8466 = (inp[10]) ? 8'b10100101 : 8'b10100001;
										assign node8470 = (inp[8]) ? node8476 : node8471;
											assign node8471 = (inp[9]) ? node8473 : 8'b10000101;
												assign node8473 = (inp[5]) ? 8'b10000101 : 8'b10100101;
											assign node8476 = (inp[5]) ? 8'b10000001 : node8477;
												assign node8477 = (inp[9]) ? node8481 : node8478;
													assign node8478 = (inp[10]) ? 8'b10000101 : 8'b10000001;
													assign node8481 = (inp[10]) ? 8'b10100101 : 8'b10100001;
									assign node8485 = (inp[5]) ? node8503 : node8486;
										assign node8486 = (inp[8]) ? node8492 : node8487;
											assign node8487 = (inp[9]) ? 8'b00000010 : node8488;
												assign node8488 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node8492 = (inp[10]) ? node8498 : node8493;
												assign node8493 = (inp[9]) ? 8'b10100100 : node8494;
													assign node8494 = (inp[13]) ? 8'b10000100 : 8'b10100100;
												assign node8498 = (inp[13]) ? node8500 : 8'b00000010;
													assign node8500 = (inp[9]) ? 8'b00000010 : 8'b10100000;
										assign node8503 = (inp[8]) ? node8507 : node8504;
											assign node8504 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node8507 = (inp[13]) ? 8'b10000001 : 8'b10100001;
							assign node8510 = (inp[6]) ? node8574 : node8511;
								assign node8511 = (inp[13]) ? node8531 : node8512;
									assign node8512 = (inp[8]) ? node8520 : node8513;
										assign node8513 = (inp[1]) ? node8515 : 8'b11110101;
											assign node8515 = (inp[3]) ? node8517 : 8'b10110100;
												assign node8517 = (inp[5]) ? 8'b10110100 : 8'b11110101;
										assign node8520 = (inp[5]) ? node8528 : node8521;
											assign node8521 = (inp[10]) ? node8523 : 8'b10110001;
												assign node8523 = (inp[3]) ? 8'b11110101 : node8524;
													assign node8524 = (inp[1]) ? 8'b10110100 : 8'b11110101;
											assign node8528 = (inp[1]) ? 8'b10110000 : 8'b10110001;
									assign node8531 = (inp[8]) ? node8547 : node8532;
										assign node8532 = (inp[1]) ? node8538 : node8533;
											assign node8533 = (inp[9]) ? node8535 : 8'b10010101;
												assign node8535 = (inp[5]) ? 8'b10010101 : 8'b11110101;
											assign node8538 = (inp[5]) ? 8'b10010100 : node8539;
												assign node8539 = (inp[9]) ? node8543 : node8540;
													assign node8540 = (inp[3]) ? 8'b10010101 : 8'b10010100;
													assign node8543 = (inp[3]) ? 8'b11110101 : 8'b10110100;
										assign node8547 = (inp[5]) ? node8571 : node8548;
											assign node8548 = (inp[9]) ? node8560 : node8549;
												assign node8549 = (inp[10]) ? node8555 : node8550;
													assign node8550 = (inp[1]) ? node8552 : 8'b10010001;
														assign node8552 = (inp[3]) ? 8'b10010001 : 8'b10010000;
													assign node8555 = (inp[1]) ? node8557 : 8'b10010101;
														assign node8557 = (inp[3]) ? 8'b10010101 : 8'b10010100;
												assign node8560 = (inp[10]) ? node8566 : node8561;
													assign node8561 = (inp[3]) ? 8'b10110001 : node8562;
														assign node8562 = (inp[1]) ? 8'b10110000 : 8'b10110001;
													assign node8566 = (inp[1]) ? node8568 : 8'b11110101;
														assign node8568 = (inp[3]) ? 8'b11110101 : 8'b10110100;
											assign node8571 = (inp[1]) ? 8'b10010000 : 8'b10010001;
								assign node8574 = (inp[5]) ? node8622 : node8575;
									assign node8575 = (inp[1]) ? node8593 : node8576;
										assign node8576 = (inp[8]) ? node8582 : node8577;
											assign node8577 = (inp[9]) ? 8'b00000010 : node8578;
												assign node8578 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node8582 = (inp[10]) ? node8588 : node8583;
												assign node8583 = (inp[9]) ? 8'b10100100 : node8584;
													assign node8584 = (inp[13]) ? 8'b10000100 : 8'b10100100;
												assign node8588 = (inp[13]) ? node8590 : 8'b00000010;
													assign node8590 = (inp[9]) ? 8'b00000010 : 8'b10100000;
										assign node8593 = (inp[3]) ? node8607 : node8594;
											assign node8594 = (inp[8]) ? node8600 : node8595;
												assign node8595 = (inp[13]) ? node8597 : 8'b10100101;
													assign node8597 = (inp[9]) ? 8'b10100101 : 8'b10000101;
												assign node8600 = (inp[10]) ? 8'b10100101 : node8601;
													assign node8601 = (inp[13]) ? node8603 : 8'b10100001;
														assign node8603 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node8607 = (inp[10]) ? node8617 : node8608;
												assign node8608 = (inp[8]) ? node8614 : node8609;
													assign node8609 = (inp[9]) ? 8'b00000010 : node8610;
														assign node8610 = (inp[13]) ? 8'b10100000 : 8'b00000010;
													assign node8614 = (inp[9]) ? 8'b10100100 : 8'b10000100;
												assign node8617 = (inp[9]) ? 8'b00000010 : node8618;
													assign node8618 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node8622 = (inp[13]) ? node8630 : node8623;
										assign node8623 = (inp[8]) ? node8627 : node8624;
											assign node8624 = (inp[1]) ? 8'b10110100 : 8'b11110101;
											assign node8627 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node8630 = (inp[8]) ? node8634 : node8631;
											assign node8631 = (inp[1]) ? 8'b10010100 : 8'b10010101;
											assign node8634 = (inp[1]) ? 8'b10010000 : 8'b10010001;

endmodule