module dtc_split125_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node10;
	wire [15-1:0] node11;
	wire [15-1:0] node12;
	wire [15-1:0] node17;
	wire [15-1:0] node19;
	wire [15-1:0] node21;
	wire [15-1:0] node22;
	wire [15-1:0] node26;
	wire [15-1:0] node27;
	wire [15-1:0] node28;
	wire [15-1:0] node29;
	wire [15-1:0] node30;
	wire [15-1:0] node35;
	wire [15-1:0] node36;
	wire [15-1:0] node37;
	wire [15-1:0] node42;
	wire [15-1:0] node44;
	wire [15-1:0] node47;
	wire [15-1:0] node48;
	wire [15-1:0] node50;
	wire [15-1:0] node51;
	wire [15-1:0] node54;
	wire [15-1:0] node57;
	wire [15-1:0] node59;
	wire [15-1:0] node61;
	wire [15-1:0] node62;
	wire [15-1:0] node66;
	wire [15-1:0] node67;
	wire [15-1:0] node68;
	wire [15-1:0] node70;
	wire [15-1:0] node73;
	wire [15-1:0] node74;
	wire [15-1:0] node77;
	wire [15-1:0] node79;
	wire [15-1:0] node82;
	wire [15-1:0] node83;
	wire [15-1:0] node84;
	wire [15-1:0] node85;
	wire [15-1:0] node86;
	wire [15-1:0] node90;
	wire [15-1:0] node93;
	wire [15-1:0] node95;
	wire [15-1:0] node98;
	wire [15-1:0] node99;
	wire [15-1:0] node100;
	wire [15-1:0] node104;
	wire [15-1:0] node105;
	wire [15-1:0] node107;
	wire [15-1:0] node111;
	wire [15-1:0] node112;
	wire [15-1:0] node113;
	wire [15-1:0] node114;
	wire [15-1:0] node115;
	wire [15-1:0] node116;
	wire [15-1:0] node118;
	wire [15-1:0] node122;
	wire [15-1:0] node124;
	wire [15-1:0] node125;
	wire [15-1:0] node129;
	wire [15-1:0] node130;
	wire [15-1:0] node132;
	wire [15-1:0] node133;
	wire [15-1:0] node136;
	wire [15-1:0] node139;
	wire [15-1:0] node140;
	wire [15-1:0] node143;
	wire [15-1:0] node146;
	wire [15-1:0] node147;
	wire [15-1:0] node148;
	wire [15-1:0] node150;
	wire [15-1:0] node153;
	wire [15-1:0] node155;
	wire [15-1:0] node158;
	wire [15-1:0] node159;
	wire [15-1:0] node162;
	wire [15-1:0] node163;
	wire [15-1:0] node165;
	wire [15-1:0] node168;
	wire [15-1:0] node171;
	wire [15-1:0] node172;
	wire [15-1:0] node173;
	wire [15-1:0] node174;
	wire [15-1:0] node176;
	wire [15-1:0] node179;
	wire [15-1:0] node180;
	wire [15-1:0] node184;
	wire [15-1:0] node185;
	wire [15-1:0] node187;
	wire [15-1:0] node191;
	wire [15-1:0] node192;
	wire [15-1:0] node193;
	wire [15-1:0] node197;
	wire [15-1:0] node198;
	wire [15-1:0] node201;
	wire [15-1:0] node202;
	wire [15-1:0] node206;
	wire [15-1:0] node207;
	wire [15-1:0] node208;
	wire [15-1:0] node209;
	wire [15-1:0] node210;
	wire [15-1:0] node211;
	wire [15-1:0] node212;
	wire [15-1:0] node217;
	wire [15-1:0] node218;
	wire [15-1:0] node219;
	wire [15-1:0] node222;
	wire [15-1:0] node223;
	wire [15-1:0] node228;
	wire [15-1:0] node229;
	wire [15-1:0] node230;
	wire [15-1:0] node233;
	wire [15-1:0] node234;
	wire [15-1:0] node235;
	wire [15-1:0] node239;
	wire [15-1:0] node242;
	wire [15-1:0] node243;
	wire [15-1:0] node246;
	wire [15-1:0] node248;
	wire [15-1:0] node250;
	wire [15-1:0] node253;
	wire [15-1:0] node254;
	wire [15-1:0] node255;
	wire [15-1:0] node256;
	wire [15-1:0] node258;
	wire [15-1:0] node262;
	wire [15-1:0] node264;
	wire [15-1:0] node265;
	wire [15-1:0] node267;
	wire [15-1:0] node268;
	wire [15-1:0] node272;
	wire [15-1:0] node275;
	wire [15-1:0] node276;
	wire [15-1:0] node277;
	wire [15-1:0] node280;
	wire [15-1:0] node283;
	wire [15-1:0] node284;
	wire [15-1:0] node285;
	wire [15-1:0] node286;
	wire [15-1:0] node291;
	wire [15-1:0] node293;
	wire [15-1:0] node296;
	wire [15-1:0] node297;
	wire [15-1:0] node298;
	wire [15-1:0] node299;
	wire [15-1:0] node300;
	wire [15-1:0] node302;
	wire [15-1:0] node303;
	wire [15-1:0] node307;
	wire [15-1:0] node308;
	wire [15-1:0] node310;
	wire [15-1:0] node313;
	wire [15-1:0] node314;
	wire [15-1:0] node315;
	wire [15-1:0] node320;
	wire [15-1:0] node321;
	wire [15-1:0] node322;
	wire [15-1:0] node326;
	wire [15-1:0] node329;
	wire [15-1:0] node330;
	wire [15-1:0] node331;
	wire [15-1:0] node334;
	wire [15-1:0] node337;
	wire [15-1:0] node338;
	wire [15-1:0] node339;
	wire [15-1:0] node342;
	wire [15-1:0] node344;
	wire [15-1:0] node347;
	wire [15-1:0] node350;
	wire [15-1:0] node351;
	wire [15-1:0] node352;
	wire [15-1:0] node354;
	wire [15-1:0] node357;
	wire [15-1:0] node358;
	wire [15-1:0] node359;
	wire [15-1:0] node363;
	wire [15-1:0] node365;
	wire [15-1:0] node366;
	wire [15-1:0] node370;
	wire [15-1:0] node371;
	wire [15-1:0] node372;
	wire [15-1:0] node375;
	wire [15-1:0] node378;
	wire [15-1:0] node379;
	wire [15-1:0] node382;
	wire [15-1:0] node385;
	wire [15-1:0] node386;
	wire [15-1:0] node387;
	wire [15-1:0] node388;
	wire [15-1:0] node389;
	wire [15-1:0] node390;
	wire [15-1:0] node391;
	wire [15-1:0] node395;
	wire [15-1:0] node396;
	wire [15-1:0] node400;
	wire [15-1:0] node401;
	wire [15-1:0] node402;
	wire [15-1:0] node403;
	wire [15-1:0] node404;
	wire [15-1:0] node408;
	wire [15-1:0] node411;
	wire [15-1:0] node414;
	wire [15-1:0] node415;
	wire [15-1:0] node416;
	wire [15-1:0] node417;
	wire [15-1:0] node419;
	wire [15-1:0] node423;
	wire [15-1:0] node424;
	wire [15-1:0] node428;
	wire [15-1:0] node431;
	wire [15-1:0] node432;
	wire [15-1:0] node433;
	wire [15-1:0] node434;
	wire [15-1:0] node437;
	wire [15-1:0] node439;
	wire [15-1:0] node442;
	wire [15-1:0] node443;
	wire [15-1:0] node445;
	wire [15-1:0] node446;
	wire [15-1:0] node450;
	wire [15-1:0] node451;
	wire [15-1:0] node455;
	wire [15-1:0] node457;
	wire [15-1:0] node459;
	wire [15-1:0] node460;
	wire [15-1:0] node464;
	wire [15-1:0] node465;
	wire [15-1:0] node466;
	wire [15-1:0] node467;
	wire [15-1:0] node468;
	wire [15-1:0] node470;
	wire [15-1:0] node473;
	wire [15-1:0] node474;
	wire [15-1:0] node476;
	wire [15-1:0] node480;
	wire [15-1:0] node481;
	wire [15-1:0] node482;
	wire [15-1:0] node487;
	wire [15-1:0] node488;
	wire [15-1:0] node489;
	wire [15-1:0] node490;
	wire [15-1:0] node491;
	wire [15-1:0] node493;
	wire [15-1:0] node498;
	wire [15-1:0] node501;
	wire [15-1:0] node502;
	wire [15-1:0] node503;
	wire [15-1:0] node507;
	wire [15-1:0] node509;
	wire [15-1:0] node511;
	wire [15-1:0] node514;
	wire [15-1:0] node515;
	wire [15-1:0] node516;
	wire [15-1:0] node517;
	wire [15-1:0] node518;
	wire [15-1:0] node521;
	wire [15-1:0] node524;
	wire [15-1:0] node527;
	wire [15-1:0] node528;
	wire [15-1:0] node530;
	wire [15-1:0] node531;
	wire [15-1:0] node532;
	wire [15-1:0] node537;
	wire [15-1:0] node538;
	wire [15-1:0] node541;
	wire [15-1:0] node544;
	wire [15-1:0] node545;
	wire [15-1:0] node547;
	wire [15-1:0] node550;
	wire [15-1:0] node551;
	wire [15-1:0] node554;
	wire [15-1:0] node557;
	wire [15-1:0] node558;
	wire [15-1:0] node559;
	wire [15-1:0] node560;
	wire [15-1:0] node561;
	wire [15-1:0] node562;
	wire [15-1:0] node564;
	wire [15-1:0] node568;
	wire [15-1:0] node569;
	wire [15-1:0] node570;
	wire [15-1:0] node574;
	wire [15-1:0] node576;
	wire [15-1:0] node579;
	wire [15-1:0] node580;
	wire [15-1:0] node581;
	wire [15-1:0] node585;
	wire [15-1:0] node586;
	wire [15-1:0] node589;
	wire [15-1:0] node590;
	wire [15-1:0] node594;
	wire [15-1:0] node595;
	wire [15-1:0] node596;
	wire [15-1:0] node597;
	wire [15-1:0] node598;
	wire [15-1:0] node601;
	wire [15-1:0] node603;
	wire [15-1:0] node606;
	wire [15-1:0] node607;
	wire [15-1:0] node609;
	wire [15-1:0] node613;
	wire [15-1:0] node614;
	wire [15-1:0] node615;
	wire [15-1:0] node617;
	wire [15-1:0] node618;
	wire [15-1:0] node623;
	wire [15-1:0] node626;
	wire [15-1:0] node627;
	wire [15-1:0] node628;
	wire [15-1:0] node629;
	wire [15-1:0] node633;
	wire [15-1:0] node636;
	wire [15-1:0] node637;
	wire [15-1:0] node640;
	wire [15-1:0] node641;
	wire [15-1:0] node644;
	wire [15-1:0] node647;
	wire [15-1:0] node648;
	wire [15-1:0] node649;
	wire [15-1:0] node650;
	wire [15-1:0] node651;
	wire [15-1:0] node652;
	wire [15-1:0] node654;
	wire [15-1:0] node657;
	wire [15-1:0] node659;
	wire [15-1:0] node661;
	wire [15-1:0] node665;
	wire [15-1:0] node666;
	wire [15-1:0] node667;
	wire [15-1:0] node670;
	wire [15-1:0] node672;
	wire [15-1:0] node675;
	wire [15-1:0] node676;
	wire [15-1:0] node680;
	wire [15-1:0] node681;
	wire [15-1:0] node682;
	wire [15-1:0] node683;
	wire [15-1:0] node684;
	wire [15-1:0] node686;
	wire [15-1:0] node690;
	wire [15-1:0] node693;
	wire [15-1:0] node695;
	wire [15-1:0] node698;
	wire [15-1:0] node699;
	wire [15-1:0] node701;
	wire [15-1:0] node704;
	wire [15-1:0] node706;
	wire [15-1:0] node709;
	wire [15-1:0] node710;
	wire [15-1:0] node711;
	wire [15-1:0] node712;
	wire [15-1:0] node713;
	wire [15-1:0] node714;
	wire [15-1:0] node717;
	wire [15-1:0] node721;
	wire [15-1:0] node722;
	wire [15-1:0] node724;
	wire [15-1:0] node728;
	wire [15-1:0] node729;
	wire [15-1:0] node730;
	wire [15-1:0] node731;
	wire [15-1:0] node736;
	wire [15-1:0] node737;
	wire [15-1:0] node740;
	wire [15-1:0] node741;
	wire [15-1:0] node743;
	wire [15-1:0] node747;
	wire [15-1:0] node748;
	wire [15-1:0] node749;
	wire [15-1:0] node750;
	wire [15-1:0] node752;
	wire [15-1:0] node755;
	wire [15-1:0] node757;
	wire [15-1:0] node760;
	wire [15-1:0] node762;
	wire [15-1:0] node763;
	wire [15-1:0] node767;
	wire [15-1:0] node768;
	wire [15-1:0] node769;
	wire [15-1:0] node771;
	wire [15-1:0] node775;
	wire [15-1:0] node776;
	wire [15-1:0] node780;
	wire [15-1:0] node781;
	wire [15-1:0] node782;
	wire [15-1:0] node783;
	wire [15-1:0] node784;
	wire [15-1:0] node785;
	wire [15-1:0] node786;
	wire [15-1:0] node787;
	wire [15-1:0] node788;
	wire [15-1:0] node789;
	wire [15-1:0] node793;
	wire [15-1:0] node794;
	wire [15-1:0] node798;
	wire [15-1:0] node800;
	wire [15-1:0] node803;
	wire [15-1:0] node805;
	wire [15-1:0] node807;
	wire [15-1:0] node810;
	wire [15-1:0] node811;
	wire [15-1:0] node813;
	wire [15-1:0] node816;
	wire [15-1:0] node817;
	wire [15-1:0] node818;
	wire [15-1:0] node819;
	wire [15-1:0] node825;
	wire [15-1:0] node826;
	wire [15-1:0] node827;
	wire [15-1:0] node828;
	wire [15-1:0] node830;
	wire [15-1:0] node834;
	wire [15-1:0] node836;
	wire [15-1:0] node838;
	wire [15-1:0] node841;
	wire [15-1:0] node842;
	wire [15-1:0] node843;
	wire [15-1:0] node845;
	wire [15-1:0] node846;
	wire [15-1:0] node848;
	wire [15-1:0] node849;
	wire [15-1:0] node854;
	wire [15-1:0] node856;
	wire [15-1:0] node859;
	wire [15-1:0] node860;
	wire [15-1:0] node863;
	wire [15-1:0] node865;
	wire [15-1:0] node867;
	wire [15-1:0] node870;
	wire [15-1:0] node871;
	wire [15-1:0] node872;
	wire [15-1:0] node873;
	wire [15-1:0] node874;
	wire [15-1:0] node875;
	wire [15-1:0] node877;
	wire [15-1:0] node881;
	wire [15-1:0] node883;
	wire [15-1:0] node886;
	wire [15-1:0] node887;
	wire [15-1:0] node890;
	wire [15-1:0] node893;
	wire [15-1:0] node894;
	wire [15-1:0] node895;
	wire [15-1:0] node898;
	wire [15-1:0] node899;
	wire [15-1:0] node900;
	wire [15-1:0] node904;
	wire [15-1:0] node905;
	wire [15-1:0] node908;
	wire [15-1:0] node911;
	wire [15-1:0] node912;
	wire [15-1:0] node915;
	wire [15-1:0] node918;
	wire [15-1:0] node919;
	wire [15-1:0] node920;
	wire [15-1:0] node921;
	wire [15-1:0] node922;
	wire [15-1:0] node923;
	wire [15-1:0] node928;
	wire [15-1:0] node931;
	wire [15-1:0] node933;
	wire [15-1:0] node935;
	wire [15-1:0] node938;
	wire [15-1:0] node939;
	wire [15-1:0] node941;
	wire [15-1:0] node943;
	wire [15-1:0] node944;
	wire [15-1:0] node947;
	wire [15-1:0] node950;
	wire [15-1:0] node951;
	wire [15-1:0] node952;
	wire [15-1:0] node956;
	wire [15-1:0] node959;
	wire [15-1:0] node960;
	wire [15-1:0] node961;
	wire [15-1:0] node962;
	wire [15-1:0] node963;
	wire [15-1:0] node964;
	wire [15-1:0] node965;
	wire [15-1:0] node970;
	wire [15-1:0] node971;
	wire [15-1:0] node972;
	wire [15-1:0] node976;
	wire [15-1:0] node977;
	wire [15-1:0] node978;
	wire [15-1:0] node982;
	wire [15-1:0] node985;
	wire [15-1:0] node986;
	wire [15-1:0] node987;
	wire [15-1:0] node988;
	wire [15-1:0] node989;
	wire [15-1:0] node993;
	wire [15-1:0] node994;
	wire [15-1:0] node999;
	wire [15-1:0] node1000;
	wire [15-1:0] node1002;
	wire [15-1:0] node1006;
	wire [15-1:0] node1007;
	wire [15-1:0] node1008;
	wire [15-1:0] node1009;
	wire [15-1:0] node1013;
	wire [15-1:0] node1014;
	wire [15-1:0] node1015;
	wire [15-1:0] node1017;
	wire [15-1:0] node1018;
	wire [15-1:0] node1022;
	wire [15-1:0] node1025;
	wire [15-1:0] node1028;
	wire [15-1:0] node1029;
	wire [15-1:0] node1030;
	wire [15-1:0] node1034;
	wire [15-1:0] node1035;
	wire [15-1:0] node1037;
	wire [15-1:0] node1038;
	wire [15-1:0] node1042;
	wire [15-1:0] node1045;
	wire [15-1:0] node1046;
	wire [15-1:0] node1047;
	wire [15-1:0] node1048;
	wire [15-1:0] node1049;
	wire [15-1:0] node1050;
	wire [15-1:0] node1053;
	wire [15-1:0] node1056;
	wire [15-1:0] node1058;
	wire [15-1:0] node1061;
	wire [15-1:0] node1062;
	wire [15-1:0] node1065;
	wire [15-1:0] node1068;
	wire [15-1:0] node1069;
	wire [15-1:0] node1070;
	wire [15-1:0] node1072;
	wire [15-1:0] node1076;
	wire [15-1:0] node1077;
	wire [15-1:0] node1078;
	wire [15-1:0] node1082;
	wire [15-1:0] node1083;
	wire [15-1:0] node1084;
	wire [15-1:0] node1088;
	wire [15-1:0] node1091;
	wire [15-1:0] node1092;
	wire [15-1:0] node1093;
	wire [15-1:0] node1095;
	wire [15-1:0] node1098;
	wire [15-1:0] node1099;
	wire [15-1:0] node1101;
	wire [15-1:0] node1104;
	wire [15-1:0] node1107;
	wire [15-1:0] node1108;
	wire [15-1:0] node1109;
	wire [15-1:0] node1111;
	wire [15-1:0] node1112;
	wire [15-1:0] node1116;
	wire [15-1:0] node1117;
	wire [15-1:0] node1120;
	wire [15-1:0] node1123;
	wire [15-1:0] node1124;
	wire [15-1:0] node1126;
	wire [15-1:0] node1129;
	wire [15-1:0] node1132;
	wire [15-1:0] node1133;
	wire [15-1:0] node1134;
	wire [15-1:0] node1135;
	wire [15-1:0] node1136;
	wire [15-1:0] node1137;
	wire [15-1:0] node1138;
	wire [15-1:0] node1139;
	wire [15-1:0] node1141;
	wire [15-1:0] node1144;
	wire [15-1:0] node1147;
	wire [15-1:0] node1149;
	wire [15-1:0] node1150;
	wire [15-1:0] node1154;
	wire [15-1:0] node1155;
	wire [15-1:0] node1157;
	wire [15-1:0] node1161;
	wire [15-1:0] node1162;
	wire [15-1:0] node1163;
	wire [15-1:0] node1165;
	wire [15-1:0] node1166;
	wire [15-1:0] node1171;
	wire [15-1:0] node1172;
	wire [15-1:0] node1174;
	wire [15-1:0] node1176;
	wire [15-1:0] node1177;
	wire [15-1:0] node1181;
	wire [15-1:0] node1184;
	wire [15-1:0] node1185;
	wire [15-1:0] node1186;
	wire [15-1:0] node1187;
	wire [15-1:0] node1188;
	wire [15-1:0] node1192;
	wire [15-1:0] node1194;
	wire [15-1:0] node1197;
	wire [15-1:0] node1198;
	wire [15-1:0] node1201;
	wire [15-1:0] node1204;
	wire [15-1:0] node1205;
	wire [15-1:0] node1206;
	wire [15-1:0] node1209;
	wire [15-1:0] node1211;
	wire [15-1:0] node1212;
	wire [15-1:0] node1216;
	wire [15-1:0] node1217;
	wire [15-1:0] node1218;
	wire [15-1:0] node1219;
	wire [15-1:0] node1223;
	wire [15-1:0] node1225;
	wire [15-1:0] node1229;
	wire [15-1:0] node1230;
	wire [15-1:0] node1231;
	wire [15-1:0] node1232;
	wire [15-1:0] node1234;
	wire [15-1:0] node1236;
	wire [15-1:0] node1237;
	wire [15-1:0] node1239;
	wire [15-1:0] node1243;
	wire [15-1:0] node1244;
	wire [15-1:0] node1248;
	wire [15-1:0] node1249;
	wire [15-1:0] node1250;
	wire [15-1:0] node1253;
	wire [15-1:0] node1255;
	wire [15-1:0] node1256;
	wire [15-1:0] node1258;
	wire [15-1:0] node1262;
	wire [15-1:0] node1263;
	wire [15-1:0] node1264;
	wire [15-1:0] node1267;
	wire [15-1:0] node1269;
	wire [15-1:0] node1272;
	wire [15-1:0] node1273;
	wire [15-1:0] node1275;
	wire [15-1:0] node1276;
	wire [15-1:0] node1280;
	wire [15-1:0] node1283;
	wire [15-1:0] node1284;
	wire [15-1:0] node1285;
	wire [15-1:0] node1286;
	wire [15-1:0] node1290;
	wire [15-1:0] node1291;
	wire [15-1:0] node1292;
	wire [15-1:0] node1296;
	wire [15-1:0] node1298;
	wire [15-1:0] node1301;
	wire [15-1:0] node1302;
	wire [15-1:0] node1304;
	wire [15-1:0] node1307;
	wire [15-1:0] node1308;
	wire [15-1:0] node1309;
	wire [15-1:0] node1313;
	wire [15-1:0] node1314;
	wire [15-1:0] node1318;
	wire [15-1:0] node1319;
	wire [15-1:0] node1320;
	wire [15-1:0] node1321;
	wire [15-1:0] node1322;
	wire [15-1:0] node1323;
	wire [15-1:0] node1324;
	wire [15-1:0] node1328;
	wire [15-1:0] node1329;
	wire [15-1:0] node1330;
	wire [15-1:0] node1334;
	wire [15-1:0] node1335;
	wire [15-1:0] node1339;
	wire [15-1:0] node1340;
	wire [15-1:0] node1341;
	wire [15-1:0] node1346;
	wire [15-1:0] node1347;
	wire [15-1:0] node1348;
	wire [15-1:0] node1349;
	wire [15-1:0] node1351;
	wire [15-1:0] node1355;
	wire [15-1:0] node1358;
	wire [15-1:0] node1360;
	wire [15-1:0] node1363;
	wire [15-1:0] node1364;
	wire [15-1:0] node1365;
	wire [15-1:0] node1368;
	wire [15-1:0] node1369;
	wire [15-1:0] node1370;
	wire [15-1:0] node1374;
	wire [15-1:0] node1375;
	wire [15-1:0] node1379;
	wire [15-1:0] node1380;
	wire [15-1:0] node1381;
	wire [15-1:0] node1384;
	wire [15-1:0] node1385;
	wire [15-1:0] node1389;
	wire [15-1:0] node1390;
	wire [15-1:0] node1394;
	wire [15-1:0] node1395;
	wire [15-1:0] node1396;
	wire [15-1:0] node1397;
	wire [15-1:0] node1398;
	wire [15-1:0] node1402;
	wire [15-1:0] node1403;
	wire [15-1:0] node1404;
	wire [15-1:0] node1406;
	wire [15-1:0] node1409;
	wire [15-1:0] node1411;
	wire [15-1:0] node1414;
	wire [15-1:0] node1416;
	wire [15-1:0] node1419;
	wire [15-1:0] node1420;
	wire [15-1:0] node1421;
	wire [15-1:0] node1422;
	wire [15-1:0] node1423;
	wire [15-1:0] node1425;
	wire [15-1:0] node1431;
	wire [15-1:0] node1433;
	wire [15-1:0] node1434;
	wire [15-1:0] node1437;
	wire [15-1:0] node1440;
	wire [15-1:0] node1441;
	wire [15-1:0] node1442;
	wire [15-1:0] node1443;
	wire [15-1:0] node1446;
	wire [15-1:0] node1449;
	wire [15-1:0] node1451;
	wire [15-1:0] node1453;
	wire [15-1:0] node1456;
	wire [15-1:0] node1457;
	wire [15-1:0] node1458;
	wire [15-1:0] node1461;
	wire [15-1:0] node1462;
	wire [15-1:0] node1466;
	wire [15-1:0] node1468;
	wire [15-1:0] node1469;
	wire [15-1:0] node1473;
	wire [15-1:0] node1474;
	wire [15-1:0] node1475;
	wire [15-1:0] node1476;
	wire [15-1:0] node1477;
	wire [15-1:0] node1478;
	wire [15-1:0] node1479;
	wire [15-1:0] node1480;
	wire [15-1:0] node1481;
	wire [15-1:0] node1483;
	wire [15-1:0] node1486;
	wire [15-1:0] node1487;
	wire [15-1:0] node1491;
	wire [15-1:0] node1494;
	wire [15-1:0] node1495;
	wire [15-1:0] node1496;
	wire [15-1:0] node1500;
	wire [15-1:0] node1501;
	wire [15-1:0] node1502;
	wire [15-1:0] node1504;
	wire [15-1:0] node1509;
	wire [15-1:0] node1510;
	wire [15-1:0] node1511;
	wire [15-1:0] node1512;
	wire [15-1:0] node1513;
	wire [15-1:0] node1516;
	wire [15-1:0] node1518;
	wire [15-1:0] node1522;
	wire [15-1:0] node1523;
	wire [15-1:0] node1525;
	wire [15-1:0] node1526;
	wire [15-1:0] node1530;
	wire [15-1:0] node1532;
	wire [15-1:0] node1533;
	wire [15-1:0] node1534;
	wire [15-1:0] node1539;
	wire [15-1:0] node1540;
	wire [15-1:0] node1541;
	wire [15-1:0] node1545;
	wire [15-1:0] node1546;
	wire [15-1:0] node1547;
	wire [15-1:0] node1552;
	wire [15-1:0] node1553;
	wire [15-1:0] node1554;
	wire [15-1:0] node1555;
	wire [15-1:0] node1556;
	wire [15-1:0] node1557;
	wire [15-1:0] node1558;
	wire [15-1:0] node1560;
	wire [15-1:0] node1565;
	wire [15-1:0] node1566;
	wire [15-1:0] node1568;
	wire [15-1:0] node1570;
	wire [15-1:0] node1574;
	wire [15-1:0] node1575;
	wire [15-1:0] node1579;
	wire [15-1:0] node1580;
	wire [15-1:0] node1581;
	wire [15-1:0] node1582;
	wire [15-1:0] node1586;
	wire [15-1:0] node1589;
	wire [15-1:0] node1590;
	wire [15-1:0] node1592;
	wire [15-1:0] node1595;
	wire [15-1:0] node1596;
	wire [15-1:0] node1600;
	wire [15-1:0] node1601;
	wire [15-1:0] node1602;
	wire [15-1:0] node1604;
	wire [15-1:0] node1607;
	wire [15-1:0] node1608;
	wire [15-1:0] node1609;
	wire [15-1:0] node1613;
	wire [15-1:0] node1616;
	wire [15-1:0] node1617;
	wire [15-1:0] node1619;
	wire [15-1:0] node1622;
	wire [15-1:0] node1623;
	wire [15-1:0] node1625;
	wire [15-1:0] node1626;
	wire [15-1:0] node1630;
	wire [15-1:0] node1631;
	wire [15-1:0] node1633;
	wire [15-1:0] node1637;
	wire [15-1:0] node1638;
	wire [15-1:0] node1639;
	wire [15-1:0] node1640;
	wire [15-1:0] node1641;
	wire [15-1:0] node1643;
	wire [15-1:0] node1644;
	wire [15-1:0] node1646;
	wire [15-1:0] node1649;
	wire [15-1:0] node1650;
	wire [15-1:0] node1651;
	wire [15-1:0] node1652;
	wire [15-1:0] node1658;
	wire [15-1:0] node1659;
	wire [15-1:0] node1660;
	wire [15-1:0] node1664;
	wire [15-1:0] node1665;
	wire [15-1:0] node1666;
	wire [15-1:0] node1670;
	wire [15-1:0] node1672;
	wire [15-1:0] node1675;
	wire [15-1:0] node1676;
	wire [15-1:0] node1677;
	wire [15-1:0] node1679;
	wire [15-1:0] node1682;
	wire [15-1:0] node1685;
	wire [15-1:0] node1686;
	wire [15-1:0] node1689;
	wire [15-1:0] node1690;
	wire [15-1:0] node1692;
	wire [15-1:0] node1696;
	wire [15-1:0] node1697;
	wire [15-1:0] node1698;
	wire [15-1:0] node1700;
	wire [15-1:0] node1703;
	wire [15-1:0] node1704;
	wire [15-1:0] node1707;
	wire [15-1:0] node1708;
	wire [15-1:0] node1711;
	wire [15-1:0] node1712;
	wire [15-1:0] node1716;
	wire [15-1:0] node1717;
	wire [15-1:0] node1718;
	wire [15-1:0] node1720;
	wire [15-1:0] node1721;
	wire [15-1:0] node1726;
	wire [15-1:0] node1727;
	wire [15-1:0] node1728;
	wire [15-1:0] node1732;
	wire [15-1:0] node1734;
	wire [15-1:0] node1735;
	wire [15-1:0] node1739;
	wire [15-1:0] node1740;
	wire [15-1:0] node1741;
	wire [15-1:0] node1742;
	wire [15-1:0] node1744;
	wire [15-1:0] node1747;
	wire [15-1:0] node1749;
	wire [15-1:0] node1752;
	wire [15-1:0] node1753;
	wire [15-1:0] node1754;
	wire [15-1:0] node1757;
	wire [15-1:0] node1758;
	wire [15-1:0] node1762;
	wire [15-1:0] node1763;
	wire [15-1:0] node1767;
	wire [15-1:0] node1768;
	wire [15-1:0] node1769;
	wire [15-1:0] node1770;
	wire [15-1:0] node1773;
	wire [15-1:0] node1775;
	wire [15-1:0] node1776;
	wire [15-1:0] node1780;
	wire [15-1:0] node1781;
	wire [15-1:0] node1783;
	wire [15-1:0] node1785;
	wire [15-1:0] node1788;
	wire [15-1:0] node1791;
	wire [15-1:0] node1792;
	wire [15-1:0] node1793;
	wire [15-1:0] node1796;
	wire [15-1:0] node1797;
	wire [15-1:0] node1801;
	wire [15-1:0] node1803;
	wire [15-1:0] node1806;
	wire [15-1:0] node1807;
	wire [15-1:0] node1808;
	wire [15-1:0] node1809;
	wire [15-1:0] node1810;
	wire [15-1:0] node1811;
	wire [15-1:0] node1812;
	wire [15-1:0] node1813;
	wire [15-1:0] node1817;
	wire [15-1:0] node1818;
	wire [15-1:0] node1821;
	wire [15-1:0] node1824;
	wire [15-1:0] node1825;
	wire [15-1:0] node1826;
	wire [15-1:0] node1831;
	wire [15-1:0] node1832;
	wire [15-1:0] node1833;
	wire [15-1:0] node1836;
	wire [15-1:0] node1837;
	wire [15-1:0] node1838;
	wire [15-1:0] node1842;
	wire [15-1:0] node1843;
	wire [15-1:0] node1847;
	wire [15-1:0] node1848;
	wire [15-1:0] node1850;
	wire [15-1:0] node1853;
	wire [15-1:0] node1854;
	wire [15-1:0] node1858;
	wire [15-1:0] node1859;
	wire [15-1:0] node1860;
	wire [15-1:0] node1861;
	wire [15-1:0] node1862;
	wire [15-1:0] node1863;
	wire [15-1:0] node1867;
	wire [15-1:0] node1870;
	wire [15-1:0] node1873;
	wire [15-1:0] node1874;
	wire [15-1:0] node1875;
	wire [15-1:0] node1877;
	wire [15-1:0] node1881;
	wire [15-1:0] node1883;
	wire [15-1:0] node1886;
	wire [15-1:0] node1887;
	wire [15-1:0] node1888;
	wire [15-1:0] node1889;
	wire [15-1:0] node1892;
	wire [15-1:0] node1893;
	wire [15-1:0] node1897;
	wire [15-1:0] node1898;
	wire [15-1:0] node1902;
	wire [15-1:0] node1904;
	wire [15-1:0] node1906;
	wire [15-1:0] node1909;
	wire [15-1:0] node1910;
	wire [15-1:0] node1911;
	wire [15-1:0] node1912;
	wire [15-1:0] node1913;
	wire [15-1:0] node1914;
	wire [15-1:0] node1915;
	wire [15-1:0] node1920;
	wire [15-1:0] node1923;
	wire [15-1:0] node1924;
	wire [15-1:0] node1926;
	wire [15-1:0] node1927;
	wire [15-1:0] node1931;
	wire [15-1:0] node1932;
	wire [15-1:0] node1934;
	wire [15-1:0] node1938;
	wire [15-1:0] node1939;
	wire [15-1:0] node1940;
	wire [15-1:0] node1942;
	wire [15-1:0] node1944;
	wire [15-1:0] node1945;
	wire [15-1:0] node1949;
	wire [15-1:0] node1950;
	wire [15-1:0] node1953;
	wire [15-1:0] node1954;
	wire [15-1:0] node1958;
	wire [15-1:0] node1960;
	wire [15-1:0] node1961;
	wire [15-1:0] node1962;
	wire [15-1:0] node1966;
	wire [15-1:0] node1967;
	wire [15-1:0] node1971;
	wire [15-1:0] node1972;
	wire [15-1:0] node1973;
	wire [15-1:0] node1974;
	wire [15-1:0] node1975;
	wire [15-1:0] node1979;
	wire [15-1:0] node1982;
	wire [15-1:0] node1983;
	wire [15-1:0] node1984;
	wire [15-1:0] node1988;
	wire [15-1:0] node1991;
	wire [15-1:0] node1992;
	wire [15-1:0] node1993;
	wire [15-1:0] node1994;
	wire [15-1:0] node1997;
	wire [15-1:0] node2001;
	wire [15-1:0] node2002;
	wire [15-1:0] node2005;
	wire [15-1:0] node2008;
	wire [15-1:0] node2009;
	wire [15-1:0] node2010;
	wire [15-1:0] node2011;
	wire [15-1:0] node2012;
	wire [15-1:0] node2013;
	wire [15-1:0] node2016;
	wire [15-1:0] node2019;
	wire [15-1:0] node2020;
	wire [15-1:0] node2024;
	wire [15-1:0] node2025;
	wire [15-1:0] node2026;
	wire [15-1:0] node2029;
	wire [15-1:0] node2030;
	wire [15-1:0] node2033;
	wire [15-1:0] node2034;
	wire [15-1:0] node2039;
	wire [15-1:0] node2040;
	wire [15-1:0] node2041;
	wire [15-1:0] node2042;
	wire [15-1:0] node2045;
	wire [15-1:0] node2046;
	wire [15-1:0] node2050;
	wire [15-1:0] node2051;
	wire [15-1:0] node2052;
	wire [15-1:0] node2053;
	wire [15-1:0] node2058;
	wire [15-1:0] node2061;
	wire [15-1:0] node2062;
	wire [15-1:0] node2063;
	wire [15-1:0] node2065;
	wire [15-1:0] node2066;
	wire [15-1:0] node2071;
	wire [15-1:0] node2072;
	wire [15-1:0] node2074;
	wire [15-1:0] node2077;
	wire [15-1:0] node2079;
	wire [15-1:0] node2081;
	wire [15-1:0] node2083;
	wire [15-1:0] node2086;
	wire [15-1:0] node2087;
	wire [15-1:0] node2088;
	wire [15-1:0] node2089;
	wire [15-1:0] node2091;
	wire [15-1:0] node2094;
	wire [15-1:0] node2095;
	wire [15-1:0] node2098;
	wire [15-1:0] node2100;
	wire [15-1:0] node2102;
	wire [15-1:0] node2105;
	wire [15-1:0] node2106;
	wire [15-1:0] node2107;
	wire [15-1:0] node2108;
	wire [15-1:0] node2109;
	wire [15-1:0] node2113;
	wire [15-1:0] node2114;
	wire [15-1:0] node2118;
	wire [15-1:0] node2119;
	wire [15-1:0] node2123;
	wire [15-1:0] node2124;
	wire [15-1:0] node2127;
	wire [15-1:0] node2128;
	wire [15-1:0] node2130;
	wire [15-1:0] node2131;
	wire [15-1:0] node2136;
	wire [15-1:0] node2137;
	wire [15-1:0] node2138;
	wire [15-1:0] node2139;
	wire [15-1:0] node2142;
	wire [15-1:0] node2144;
	wire [15-1:0] node2147;
	wire [15-1:0] node2148;
	wire [15-1:0] node2149;
	wire [15-1:0] node2153;
	wire [15-1:0] node2156;
	wire [15-1:0] node2157;
	wire [15-1:0] node2158;
	wire [15-1:0] node2159;
	wire [15-1:0] node2160;
	wire [15-1:0] node2164;
	wire [15-1:0] node2165;
	wire [15-1:0] node2168;
	wire [15-1:0] node2172;
	wire [15-1:0] node2173;
	wire [15-1:0] node2174;
	wire [15-1:0] node2176;
	wire [15-1:0] node2179;
	wire [15-1:0] node2182;
	wire [15-1:0] node2185;
	wire [15-1:0] node2186;
	wire [15-1:0] node2187;
	wire [15-1:0] node2188;
	wire [15-1:0] node2189;
	wire [15-1:0] node2190;
	wire [15-1:0] node2191;
	wire [15-1:0] node2192;
	wire [15-1:0] node2193;
	wire [15-1:0] node2196;
	wire [15-1:0] node2199;
	wire [15-1:0] node2201;
	wire [15-1:0] node2202;
	wire [15-1:0] node2206;
	wire [15-1:0] node2207;
	wire [15-1:0] node2210;
	wire [15-1:0] node2213;
	wire [15-1:0] node2214;
	wire [15-1:0] node2215;
	wire [15-1:0] node2217;
	wire [15-1:0] node2220;
	wire [15-1:0] node2221;
	wire [15-1:0] node2225;
	wire [15-1:0] node2226;
	wire [15-1:0] node2228;
	wire [15-1:0] node2229;
	wire [15-1:0] node2233;
	wire [15-1:0] node2236;
	wire [15-1:0] node2237;
	wire [15-1:0] node2238;
	wire [15-1:0] node2239;
	wire [15-1:0] node2242;
	wire [15-1:0] node2243;
	wire [15-1:0] node2247;
	wire [15-1:0] node2249;
	wire [15-1:0] node2252;
	wire [15-1:0] node2253;
	wire [15-1:0] node2254;
	wire [15-1:0] node2258;
	wire [15-1:0] node2259;
	wire [15-1:0] node2260;
	wire [15-1:0] node2261;
	wire [15-1:0] node2265;
	wire [15-1:0] node2268;
	wire [15-1:0] node2270;
	wire [15-1:0] node2273;
	wire [15-1:0] node2274;
	wire [15-1:0] node2275;
	wire [15-1:0] node2276;
	wire [15-1:0] node2278;
	wire [15-1:0] node2279;
	wire [15-1:0] node2283;
	wire [15-1:0] node2284;
	wire [15-1:0] node2285;
	wire [15-1:0] node2290;
	wire [15-1:0] node2291;
	wire [15-1:0] node2292;
	wire [15-1:0] node2294;
	wire [15-1:0] node2295;
	wire [15-1:0] node2299;
	wire [15-1:0] node2300;
	wire [15-1:0] node2302;
	wire [15-1:0] node2306;
	wire [15-1:0] node2307;
	wire [15-1:0] node2310;
	wire [15-1:0] node2311;
	wire [15-1:0] node2314;
	wire [15-1:0] node2317;
	wire [15-1:0] node2318;
	wire [15-1:0] node2319;
	wire [15-1:0] node2320;
	wire [15-1:0] node2322;
	wire [15-1:0] node2325;
	wire [15-1:0] node2326;
	wire [15-1:0] node2330;
	wire [15-1:0] node2331;
	wire [15-1:0] node2333;
	wire [15-1:0] node2336;
	wire [15-1:0] node2337;
	wire [15-1:0] node2341;
	wire [15-1:0] node2342;
	wire [15-1:0] node2344;
	wire [15-1:0] node2347;
	wire [15-1:0] node2348;
	wire [15-1:0] node2350;
	wire [15-1:0] node2353;
	wire [15-1:0] node2355;
	wire [15-1:0] node2356;
	wire [15-1:0] node2360;
	wire [15-1:0] node2361;
	wire [15-1:0] node2362;
	wire [15-1:0] node2363;
	wire [15-1:0] node2364;
	wire [15-1:0] node2365;
	wire [15-1:0] node2366;
	wire [15-1:0] node2367;
	wire [15-1:0] node2371;
	wire [15-1:0] node2372;
	wire [15-1:0] node2376;
	wire [15-1:0] node2379;
	wire [15-1:0] node2380;
	wire [15-1:0] node2383;
	wire [15-1:0] node2386;
	wire [15-1:0] node2387;
	wire [15-1:0] node2388;
	wire [15-1:0] node2390;
	wire [15-1:0] node2393;
	wire [15-1:0] node2396;
	wire [15-1:0] node2397;
	wire [15-1:0] node2398;
	wire [15-1:0] node2400;
	wire [15-1:0] node2405;
	wire [15-1:0] node2406;
	wire [15-1:0] node2407;
	wire [15-1:0] node2408;
	wire [15-1:0] node2411;
	wire [15-1:0] node2413;
	wire [15-1:0] node2416;
	wire [15-1:0] node2417;
	wire [15-1:0] node2418;
	wire [15-1:0] node2420;
	wire [15-1:0] node2423;
	wire [15-1:0] node2425;
	wire [15-1:0] node2428;
	wire [15-1:0] node2429;
	wire [15-1:0] node2431;
	wire [15-1:0] node2435;
	wire [15-1:0] node2436;
	wire [15-1:0] node2438;
	wire [15-1:0] node2439;
	wire [15-1:0] node2441;
	wire [15-1:0] node2445;
	wire [15-1:0] node2446;
	wire [15-1:0] node2449;
	wire [15-1:0] node2450;
	wire [15-1:0] node2452;
	wire [15-1:0] node2454;
	wire [15-1:0] node2458;
	wire [15-1:0] node2459;
	wire [15-1:0] node2460;
	wire [15-1:0] node2461;
	wire [15-1:0] node2462;
	wire [15-1:0] node2466;
	wire [15-1:0] node2467;
	wire [15-1:0] node2468;
	wire [15-1:0] node2471;
	wire [15-1:0] node2474;
	wire [15-1:0] node2475;
	wire [15-1:0] node2478;
	wire [15-1:0] node2479;
	wire [15-1:0] node2483;
	wire [15-1:0] node2484;
	wire [15-1:0] node2485;
	wire [15-1:0] node2486;
	wire [15-1:0] node2490;
	wire [15-1:0] node2491;
	wire [15-1:0] node2494;
	wire [15-1:0] node2497;
	wire [15-1:0] node2498;
	wire [15-1:0] node2500;
	wire [15-1:0] node2502;
	wire [15-1:0] node2505;
	wire [15-1:0] node2506;
	wire [15-1:0] node2508;
	wire [15-1:0] node2512;
	wire [15-1:0] node2513;
	wire [15-1:0] node2514;
	wire [15-1:0] node2516;
	wire [15-1:0] node2517;
	wire [15-1:0] node2521;
	wire [15-1:0] node2522;
	wire [15-1:0] node2523;
	wire [15-1:0] node2525;
	wire [15-1:0] node2529;
	wire [15-1:0] node2530;
	wire [15-1:0] node2534;
	wire [15-1:0] node2535;
	wire [15-1:0] node2536;
	wire [15-1:0] node2539;
	wire [15-1:0] node2541;
	wire [15-1:0] node2544;
	wire [15-1:0] node2545;
	wire [15-1:0] node2547;
	wire [15-1:0] node2551;
	wire [15-1:0] node2552;
	wire [15-1:0] node2553;
	wire [15-1:0] node2554;
	wire [15-1:0] node2555;
	wire [15-1:0] node2556;
	wire [15-1:0] node2557;
	wire [15-1:0] node2559;
	wire [15-1:0] node2562;
	wire [15-1:0] node2563;
	wire [15-1:0] node2564;
	wire [15-1:0] node2568;
	wire [15-1:0] node2569;
	wire [15-1:0] node2573;
	wire [15-1:0] node2574;
	wire [15-1:0] node2575;
	wire [15-1:0] node2576;
	wire [15-1:0] node2577;
	wire [15-1:0] node2583;
	wire [15-1:0] node2586;
	wire [15-1:0] node2587;
	wire [15-1:0] node2588;
	wire [15-1:0] node2591;
	wire [15-1:0] node2592;
	wire [15-1:0] node2593;
	wire [15-1:0] node2598;
	wire [15-1:0] node2600;
	wire [15-1:0] node2601;
	wire [15-1:0] node2604;
	wire [15-1:0] node2605;
	wire [15-1:0] node2607;
	wire [15-1:0] node2611;
	wire [15-1:0] node2612;
	wire [15-1:0] node2613;
	wire [15-1:0] node2614;
	wire [15-1:0] node2618;
	wire [15-1:0] node2619;
	wire [15-1:0] node2622;
	wire [15-1:0] node2625;
	wire [15-1:0] node2626;
	wire [15-1:0] node2627;
	wire [15-1:0] node2631;
	wire [15-1:0] node2632;
	wire [15-1:0] node2634;
	wire [15-1:0] node2637;
	wire [15-1:0] node2638;
	wire [15-1:0] node2642;
	wire [15-1:0] node2643;
	wire [15-1:0] node2644;
	wire [15-1:0] node2645;
	wire [15-1:0] node2646;
	wire [15-1:0] node2649;
	wire [15-1:0] node2652;
	wire [15-1:0] node2653;
	wire [15-1:0] node2656;
	wire [15-1:0] node2657;
	wire [15-1:0] node2659;
	wire [15-1:0] node2661;
	wire [15-1:0] node2665;
	wire [15-1:0] node2666;
	wire [15-1:0] node2667;
	wire [15-1:0] node2668;
	wire [15-1:0] node2669;
	wire [15-1:0] node2675;
	wire [15-1:0] node2676;
	wire [15-1:0] node2679;
	wire [15-1:0] node2682;
	wire [15-1:0] node2683;
	wire [15-1:0] node2684;
	wire [15-1:0] node2685;
	wire [15-1:0] node2687;
	wire [15-1:0] node2690;
	wire [15-1:0] node2693;
	wire [15-1:0] node2694;
	wire [15-1:0] node2698;
	wire [15-1:0] node2699;
	wire [15-1:0] node2700;
	wire [15-1:0] node2703;
	wire [15-1:0] node2705;
	wire [15-1:0] node2708;
	wire [15-1:0] node2709;
	wire [15-1:0] node2710;
	wire [15-1:0] node2711;
	wire [15-1:0] node2716;
	wire [15-1:0] node2719;
	wire [15-1:0] node2720;
	wire [15-1:0] node2721;
	wire [15-1:0] node2722;
	wire [15-1:0] node2723;
	wire [15-1:0] node2724;
	wire [15-1:0] node2727;
	wire [15-1:0] node2729;
	wire [15-1:0] node2732;
	wire [15-1:0] node2733;
	wire [15-1:0] node2735;
	wire [15-1:0] node2737;
	wire [15-1:0] node2738;
	wire [15-1:0] node2742;
	wire [15-1:0] node2744;
	wire [15-1:0] node2747;
	wire [15-1:0] node2748;
	wire [15-1:0] node2749;
	wire [15-1:0] node2750;
	wire [15-1:0] node2753;
	wire [15-1:0] node2755;
	wire [15-1:0] node2757;
	wire [15-1:0] node2761;
	wire [15-1:0] node2762;
	wire [15-1:0] node2763;
	wire [15-1:0] node2767;
	wire [15-1:0] node2769;
	wire [15-1:0] node2770;
	wire [15-1:0] node2771;
	wire [15-1:0] node2775;
	wire [15-1:0] node2778;
	wire [15-1:0] node2779;
	wire [15-1:0] node2780;
	wire [15-1:0] node2781;
	wire [15-1:0] node2783;
	wire [15-1:0] node2786;
	wire [15-1:0] node2789;
	wire [15-1:0] node2791;
	wire [15-1:0] node2792;
	wire [15-1:0] node2793;
	wire [15-1:0] node2798;
	wire [15-1:0] node2799;
	wire [15-1:0] node2802;
	wire [15-1:0] node2803;
	wire [15-1:0] node2806;
	wire [15-1:0] node2807;
	wire [15-1:0] node2811;
	wire [15-1:0] node2812;
	wire [15-1:0] node2813;
	wire [15-1:0] node2814;
	wire [15-1:0] node2815;
	wire [15-1:0] node2816;
	wire [15-1:0] node2818;
	wire [15-1:0] node2822;
	wire [15-1:0] node2823;
	wire [15-1:0] node2824;
	wire [15-1:0] node2828;
	wire [15-1:0] node2829;
	wire [15-1:0] node2833;
	wire [15-1:0] node2834;
	wire [15-1:0] node2835;
	wire [15-1:0] node2836;
	wire [15-1:0] node2839;
	wire [15-1:0] node2842;
	wire [15-1:0] node2843;
	wire [15-1:0] node2847;
	wire [15-1:0] node2850;
	wire [15-1:0] node2851;
	wire [15-1:0] node2852;
	wire [15-1:0] node2856;
	wire [15-1:0] node2857;
	wire [15-1:0] node2858;
	wire [15-1:0] node2862;
	wire [15-1:0] node2863;
	wire [15-1:0] node2864;
	wire [15-1:0] node2867;
	wire [15-1:0] node2871;
	wire [15-1:0] node2872;
	wire [15-1:0] node2873;
	wire [15-1:0] node2874;
	wire [15-1:0] node2875;
	wire [15-1:0] node2876;
	wire [15-1:0] node2882;
	wire [15-1:0] node2884;
	wire [15-1:0] node2885;
	wire [15-1:0] node2889;
	wire [15-1:0] node2890;
	wire [15-1:0] node2891;
	wire [15-1:0] node2892;
	wire [15-1:0] node2896;
	wire [15-1:0] node2897;
	wire [15-1:0] node2900;
	wire [15-1:0] node2903;
	wire [15-1:0] node2904;
	wire [15-1:0] node2907;
	wire [15-1:0] node2908;
	wire [15-1:0] node2911;
	wire [15-1:0] node2912;
	wire [15-1:0] node2916;
	wire [15-1:0] node2917;
	wire [15-1:0] node2918;
	wire [15-1:0] node2919;
	wire [15-1:0] node2920;
	wire [15-1:0] node2921;
	wire [15-1:0] node2922;
	wire [15-1:0] node2923;
	wire [15-1:0] node2924;
	wire [15-1:0] node2925;
	wire [15-1:0] node2927;
	wire [15-1:0] node2928;
	wire [15-1:0] node2933;
	wire [15-1:0] node2934;
	wire [15-1:0] node2935;
	wire [15-1:0] node2938;
	wire [15-1:0] node2941;
	wire [15-1:0] node2942;
	wire [15-1:0] node2945;
	wire [15-1:0] node2948;
	wire [15-1:0] node2949;
	wire [15-1:0] node2950;
	wire [15-1:0] node2951;
	wire [15-1:0] node2953;
	wire [15-1:0] node2955;
	wire [15-1:0] node2959;
	wire [15-1:0] node2961;
	wire [15-1:0] node2964;
	wire [15-1:0] node2967;
	wire [15-1:0] node2968;
	wire [15-1:0] node2969;
	wire [15-1:0] node2970;
	wire [15-1:0] node2972;
	wire [15-1:0] node2973;
	wire [15-1:0] node2977;
	wire [15-1:0] node2979;
	wire [15-1:0] node2982;
	wire [15-1:0] node2983;
	wire [15-1:0] node2985;
	wire [15-1:0] node2987;
	wire [15-1:0] node2988;
	wire [15-1:0] node2992;
	wire [15-1:0] node2993;
	wire [15-1:0] node2997;
	wire [15-1:0] node2998;
	wire [15-1:0] node2999;
	wire [15-1:0] node3000;
	wire [15-1:0] node3004;
	wire [15-1:0] node3006;
	wire [15-1:0] node3007;
	wire [15-1:0] node3011;
	wire [15-1:0] node3012;
	wire [15-1:0] node3013;
	wire [15-1:0] node3015;
	wire [15-1:0] node3016;
	wire [15-1:0] node3022;
	wire [15-1:0] node3023;
	wire [15-1:0] node3024;
	wire [15-1:0] node3025;
	wire [15-1:0] node3027;
	wire [15-1:0] node3030;
	wire [15-1:0] node3031;
	wire [15-1:0] node3033;
	wire [15-1:0] node3035;
	wire [15-1:0] node3036;
	wire [15-1:0] node3037;
	wire [15-1:0] node3043;
	wire [15-1:0] node3044;
	wire [15-1:0] node3045;
	wire [15-1:0] node3047;
	wire [15-1:0] node3050;
	wire [15-1:0] node3053;
	wire [15-1:0] node3054;
	wire [15-1:0] node3056;
	wire [15-1:0] node3060;
	wire [15-1:0] node3061;
	wire [15-1:0] node3062;
	wire [15-1:0] node3063;
	wire [15-1:0] node3065;
	wire [15-1:0] node3066;
	wire [15-1:0] node3070;
	wire [15-1:0] node3071;
	wire [15-1:0] node3073;
	wire [15-1:0] node3076;
	wire [15-1:0] node3078;
	wire [15-1:0] node3081;
	wire [15-1:0] node3082;
	wire [15-1:0] node3085;
	wire [15-1:0] node3087;
	wire [15-1:0] node3090;
	wire [15-1:0] node3091;
	wire [15-1:0] node3092;
	wire [15-1:0] node3094;
	wire [15-1:0] node3098;
	wire [15-1:0] node3099;
	wire [15-1:0] node3102;
	wire [15-1:0] node3104;
	wire [15-1:0] node3106;
	wire [15-1:0] node3109;
	wire [15-1:0] node3110;
	wire [15-1:0] node3111;
	wire [15-1:0] node3112;
	wire [15-1:0] node3113;
	wire [15-1:0] node3114;
	wire [15-1:0] node3115;
	wire [15-1:0] node3116;
	wire [15-1:0] node3121;
	wire [15-1:0] node3122;
	wire [15-1:0] node3124;
	wire [15-1:0] node3128;
	wire [15-1:0] node3129;
	wire [15-1:0] node3130;
	wire [15-1:0] node3132;
	wire [15-1:0] node3136;
	wire [15-1:0] node3139;
	wire [15-1:0] node3140;
	wire [15-1:0] node3141;
	wire [15-1:0] node3144;
	wire [15-1:0] node3147;
	wire [15-1:0] node3148;
	wire [15-1:0] node3150;
	wire [15-1:0] node3153;
	wire [15-1:0] node3154;
	wire [15-1:0] node3155;
	wire [15-1:0] node3159;
	wire [15-1:0] node3162;
	wire [15-1:0] node3163;
	wire [15-1:0] node3164;
	wire [15-1:0] node3166;
	wire [15-1:0] node3168;
	wire [15-1:0] node3171;
	wire [15-1:0] node3172;
	wire [15-1:0] node3174;
	wire [15-1:0] node3177;
	wire [15-1:0] node3178;
	wire [15-1:0] node3182;
	wire [15-1:0] node3183;
	wire [15-1:0] node3184;
	wire [15-1:0] node3187;
	wire [15-1:0] node3190;
	wire [15-1:0] node3191;
	wire [15-1:0] node3193;
	wire [15-1:0] node3195;
	wire [15-1:0] node3199;
	wire [15-1:0] node3200;
	wire [15-1:0] node3201;
	wire [15-1:0] node3202;
	wire [15-1:0] node3203;
	wire [15-1:0] node3205;
	wire [15-1:0] node3208;
	wire [15-1:0] node3209;
	wire [15-1:0] node3211;
	wire [15-1:0] node3212;
	wire [15-1:0] node3217;
	wire [15-1:0] node3218;
	wire [15-1:0] node3219;
	wire [15-1:0] node3223;
	wire [15-1:0] node3224;
	wire [15-1:0] node3228;
	wire [15-1:0] node3229;
	wire [15-1:0] node3230;
	wire [15-1:0] node3233;
	wire [15-1:0] node3235;
	wire [15-1:0] node3236;
	wire [15-1:0] node3240;
	wire [15-1:0] node3241;
	wire [15-1:0] node3243;
	wire [15-1:0] node3244;
	wire [15-1:0] node3247;
	wire [15-1:0] node3250;
	wire [15-1:0] node3252;
	wire [15-1:0] node3254;
	wire [15-1:0] node3257;
	wire [15-1:0] node3258;
	wire [15-1:0] node3259;
	wire [15-1:0] node3260;
	wire [15-1:0] node3263;
	wire [15-1:0] node3266;
	wire [15-1:0] node3267;
	wire [15-1:0] node3268;
	wire [15-1:0] node3272;
	wire [15-1:0] node3273;
	wire [15-1:0] node3275;
	wire [15-1:0] node3279;
	wire [15-1:0] node3280;
	wire [15-1:0] node3281;
	wire [15-1:0] node3282;
	wire [15-1:0] node3283;
	wire [15-1:0] node3285;
	wire [15-1:0] node3289;
	wire [15-1:0] node3292;
	wire [15-1:0] node3294;
	wire [15-1:0] node3297;
	wire [15-1:0] node3298;
	wire [15-1:0] node3300;
	wire [15-1:0] node3301;
	wire [15-1:0] node3305;
	wire [15-1:0] node3308;
	wire [15-1:0] node3309;
	wire [15-1:0] node3310;
	wire [15-1:0] node3311;
	wire [15-1:0] node3312;
	wire [15-1:0] node3313;
	wire [15-1:0] node3315;
	wire [15-1:0] node3318;
	wire [15-1:0] node3319;
	wire [15-1:0] node3320;
	wire [15-1:0] node3322;
	wire [15-1:0] node3325;
	wire [15-1:0] node3326;
	wire [15-1:0] node3329;
	wire [15-1:0] node3333;
	wire [15-1:0] node3334;
	wire [15-1:0] node3335;
	wire [15-1:0] node3338;
	wire [15-1:0] node3341;
	wire [15-1:0] node3343;
	wire [15-1:0] node3344;
	wire [15-1:0] node3345;
	wire [15-1:0] node3350;
	wire [15-1:0] node3351;
	wire [15-1:0] node3352;
	wire [15-1:0] node3353;
	wire [15-1:0] node3357;
	wire [15-1:0] node3358;
	wire [15-1:0] node3360;
	wire [15-1:0] node3364;
	wire [15-1:0] node3365;
	wire [15-1:0] node3366;
	wire [15-1:0] node3369;
	wire [15-1:0] node3371;
	wire [15-1:0] node3374;
	wire [15-1:0] node3375;
	wire [15-1:0] node3376;
	wire [15-1:0] node3381;
	wire [15-1:0] node3382;
	wire [15-1:0] node3383;
	wire [15-1:0] node3384;
	wire [15-1:0] node3385;
	wire [15-1:0] node3387;
	wire [15-1:0] node3388;
	wire [15-1:0] node3393;
	wire [15-1:0] node3394;
	wire [15-1:0] node3395;
	wire [15-1:0] node3400;
	wire [15-1:0] node3401;
	wire [15-1:0] node3403;
	wire [15-1:0] node3405;
	wire [15-1:0] node3406;
	wire [15-1:0] node3410;
	wire [15-1:0] node3411;
	wire [15-1:0] node3412;
	wire [15-1:0] node3416;
	wire [15-1:0] node3418;
	wire [15-1:0] node3421;
	wire [15-1:0] node3422;
	wire [15-1:0] node3423;
	wire [15-1:0] node3424;
	wire [15-1:0] node3426;
	wire [15-1:0] node3427;
	wire [15-1:0] node3431;
	wire [15-1:0] node3433;
	wire [15-1:0] node3436;
	wire [15-1:0] node3437;
	wire [15-1:0] node3440;
	wire [15-1:0] node3442;
	wire [15-1:0] node3445;
	wire [15-1:0] node3446;
	wire [15-1:0] node3447;
	wire [15-1:0] node3450;
	wire [15-1:0] node3451;
	wire [15-1:0] node3452;
	wire [15-1:0] node3453;
	wire [15-1:0] node3458;
	wire [15-1:0] node3459;
	wire [15-1:0] node3463;
	wire [15-1:0] node3464;
	wire [15-1:0] node3465;
	wire [15-1:0] node3469;
	wire [15-1:0] node3470;
	wire [15-1:0] node3471;
	wire [15-1:0] node3475;
	wire [15-1:0] node3478;
	wire [15-1:0] node3479;
	wire [15-1:0] node3480;
	wire [15-1:0] node3481;
	wire [15-1:0] node3482;
	wire [15-1:0] node3483;
	wire [15-1:0] node3485;
	wire [15-1:0] node3488;
	wire [15-1:0] node3492;
	wire [15-1:0] node3493;
	wire [15-1:0] node3494;
	wire [15-1:0] node3495;
	wire [15-1:0] node3496;
	wire [15-1:0] node3498;
	wire [15-1:0] node3500;
	wire [15-1:0] node3505;
	wire [15-1:0] node3508;
	wire [15-1:0] node3509;
	wire [15-1:0] node3511;
	wire [15-1:0] node3514;
	wire [15-1:0] node3517;
	wire [15-1:0] node3518;
	wire [15-1:0] node3519;
	wire [15-1:0] node3520;
	wire [15-1:0] node3521;
	wire [15-1:0] node3525;
	wire [15-1:0] node3527;
	wire [15-1:0] node3530;
	wire [15-1:0] node3531;
	wire [15-1:0] node3534;
	wire [15-1:0] node3535;
	wire [15-1:0] node3538;
	wire [15-1:0] node3539;
	wire [15-1:0] node3543;
	wire [15-1:0] node3544;
	wire [15-1:0] node3545;
	wire [15-1:0] node3548;
	wire [15-1:0] node3550;
	wire [15-1:0] node3551;
	wire [15-1:0] node3553;
	wire [15-1:0] node3554;
	wire [15-1:0] node3559;
	wire [15-1:0] node3560;
	wire [15-1:0] node3563;
	wire [15-1:0] node3565;
	wire [15-1:0] node3566;
	wire [15-1:0] node3569;
	wire [15-1:0] node3572;
	wire [15-1:0] node3573;
	wire [15-1:0] node3574;
	wire [15-1:0] node3575;
	wire [15-1:0] node3576;
	wire [15-1:0] node3577;
	wire [15-1:0] node3580;
	wire [15-1:0] node3582;
	wire [15-1:0] node3585;
	wire [15-1:0] node3586;
	wire [15-1:0] node3590;
	wire [15-1:0] node3591;
	wire [15-1:0] node3592;
	wire [15-1:0] node3593;
	wire [15-1:0] node3597;
	wire [15-1:0] node3599;
	wire [15-1:0] node3600;
	wire [15-1:0] node3604;
	wire [15-1:0] node3605;
	wire [15-1:0] node3609;
	wire [15-1:0] node3610;
	wire [15-1:0] node3611;
	wire [15-1:0] node3613;
	wire [15-1:0] node3616;
	wire [15-1:0] node3617;
	wire [15-1:0] node3621;
	wire [15-1:0] node3622;
	wire [15-1:0] node3623;
	wire [15-1:0] node3627;
	wire [15-1:0] node3628;
	wire [15-1:0] node3632;
	wire [15-1:0] node3633;
	wire [15-1:0] node3634;
	wire [15-1:0] node3636;
	wire [15-1:0] node3639;
	wire [15-1:0] node3642;
	wire [15-1:0] node3643;
	wire [15-1:0] node3644;
	wire [15-1:0] node3646;
	wire [15-1:0] node3650;
	wire [15-1:0] node3651;
	wire [15-1:0] node3652;
	wire [15-1:0] node3654;
	wire [15-1:0] node3658;
	wire [15-1:0] node3659;
	wire [15-1:0] node3662;
	wire [15-1:0] node3664;
	wire [15-1:0] node3667;
	wire [15-1:0] node3668;
	wire [15-1:0] node3669;
	wire [15-1:0] node3670;
	wire [15-1:0] node3671;
	wire [15-1:0] node3672;
	wire [15-1:0] node3673;
	wire [15-1:0] node3674;
	wire [15-1:0] node3678;
	wire [15-1:0] node3679;
	wire [15-1:0] node3680;
	wire [15-1:0] node3682;
	wire [15-1:0] node3686;
	wire [15-1:0] node3687;
	wire [15-1:0] node3690;
	wire [15-1:0] node3692;
	wire [15-1:0] node3695;
	wire [15-1:0] node3697;
	wire [15-1:0] node3698;
	wire [15-1:0] node3702;
	wire [15-1:0] node3703;
	wire [15-1:0] node3704;
	wire [15-1:0] node3706;
	wire [15-1:0] node3709;
	wire [15-1:0] node3710;
	wire [15-1:0] node3712;
	wire [15-1:0] node3715;
	wire [15-1:0] node3716;
	wire [15-1:0] node3717;
	wire [15-1:0] node3720;
	wire [15-1:0] node3724;
	wire [15-1:0] node3725;
	wire [15-1:0] node3726;
	wire [15-1:0] node3728;
	wire [15-1:0] node3731;
	wire [15-1:0] node3732;
	wire [15-1:0] node3734;
	wire [15-1:0] node3737;
	wire [15-1:0] node3740;
	wire [15-1:0] node3741;
	wire [15-1:0] node3744;
	wire [15-1:0] node3745;
	wire [15-1:0] node3749;
	wire [15-1:0] node3750;
	wire [15-1:0] node3751;
	wire [15-1:0] node3752;
	wire [15-1:0] node3753;
	wire [15-1:0] node3754;
	wire [15-1:0] node3756;
	wire [15-1:0] node3761;
	wire [15-1:0] node3762;
	wire [15-1:0] node3765;
	wire [15-1:0] node3766;
	wire [15-1:0] node3767;
	wire [15-1:0] node3771;
	wire [15-1:0] node3774;
	wire [15-1:0] node3775;
	wire [15-1:0] node3776;
	wire [15-1:0] node3779;
	wire [15-1:0] node3781;
	wire [15-1:0] node3784;
	wire [15-1:0] node3785;
	wire [15-1:0] node3786;
	wire [15-1:0] node3790;
	wire [15-1:0] node3793;
	wire [15-1:0] node3794;
	wire [15-1:0] node3795;
	wire [15-1:0] node3796;
	wire [15-1:0] node3798;
	wire [15-1:0] node3802;
	wire [15-1:0] node3803;
	wire [15-1:0] node3807;
	wire [15-1:0] node3808;
	wire [15-1:0] node3809;
	wire [15-1:0] node3811;
	wire [15-1:0] node3812;
	wire [15-1:0] node3815;
	wire [15-1:0] node3818;
	wire [15-1:0] node3821;
	wire [15-1:0] node3822;
	wire [15-1:0] node3825;
	wire [15-1:0] node3827;
	wire [15-1:0] node3829;
	wire [15-1:0] node3832;
	wire [15-1:0] node3833;
	wire [15-1:0] node3834;
	wire [15-1:0] node3835;
	wire [15-1:0] node3836;
	wire [15-1:0] node3837;
	wire [15-1:0] node3840;
	wire [15-1:0] node3842;
	wire [15-1:0] node3843;
	wire [15-1:0] node3844;
	wire [15-1:0] node3849;
	wire [15-1:0] node3850;
	wire [15-1:0] node3851;
	wire [15-1:0] node3856;
	wire [15-1:0] node3857;
	wire [15-1:0] node3858;
	wire [15-1:0] node3861;
	wire [15-1:0] node3863;
	wire [15-1:0] node3866;
	wire [15-1:0] node3867;
	wire [15-1:0] node3868;
	wire [15-1:0] node3872;
	wire [15-1:0] node3875;
	wire [15-1:0] node3876;
	wire [15-1:0] node3877;
	wire [15-1:0] node3878;
	wire [15-1:0] node3880;
	wire [15-1:0] node3883;
	wire [15-1:0] node3886;
	wire [15-1:0] node3887;
	wire [15-1:0] node3890;
	wire [15-1:0] node3893;
	wire [15-1:0] node3894;
	wire [15-1:0] node3895;
	wire [15-1:0] node3898;
	wire [15-1:0] node3899;
	wire [15-1:0] node3902;
	wire [15-1:0] node3903;
	wire [15-1:0] node3905;
	wire [15-1:0] node3909;
	wire [15-1:0] node3910;
	wire [15-1:0] node3912;
	wire [15-1:0] node3915;
	wire [15-1:0] node3917;
	wire [15-1:0] node3920;
	wire [15-1:0] node3921;
	wire [15-1:0] node3922;
	wire [15-1:0] node3923;
	wire [15-1:0] node3924;
	wire [15-1:0] node3925;
	wire [15-1:0] node3929;
	wire [15-1:0] node3930;
	wire [15-1:0] node3932;
	wire [15-1:0] node3936;
	wire [15-1:0] node3937;
	wire [15-1:0] node3938;
	wire [15-1:0] node3942;
	wire [15-1:0] node3943;
	wire [15-1:0] node3947;
	wire [15-1:0] node3948;
	wire [15-1:0] node3950;
	wire [15-1:0] node3953;
	wire [15-1:0] node3956;
	wire [15-1:0] node3957;
	wire [15-1:0] node3958;
	wire [15-1:0] node3959;
	wire [15-1:0] node3962;
	wire [15-1:0] node3964;
	wire [15-1:0] node3965;
	wire [15-1:0] node3969;
	wire [15-1:0] node3970;
	wire [15-1:0] node3973;
	wire [15-1:0] node3975;
	wire [15-1:0] node3977;
	wire [15-1:0] node3980;
	wire [15-1:0] node3981;
	wire [15-1:0] node3982;
	wire [15-1:0] node3983;
	wire [15-1:0] node3987;
	wire [15-1:0] node3990;
	wire [15-1:0] node3991;
	wire [15-1:0] node3994;
	wire [15-1:0] node3997;
	wire [15-1:0] node3998;
	wire [15-1:0] node3999;
	wire [15-1:0] node4000;
	wire [15-1:0] node4001;
	wire [15-1:0] node4002;
	wire [15-1:0] node4004;
	wire [15-1:0] node4005;
	wire [15-1:0] node4006;
	wire [15-1:0] node4010;
	wire [15-1:0] node4012;
	wire [15-1:0] node4015;
	wire [15-1:0] node4016;
	wire [15-1:0] node4018;
	wire [15-1:0] node4022;
	wire [15-1:0] node4023;
	wire [15-1:0] node4024;
	wire [15-1:0] node4025;
	wire [15-1:0] node4029;
	wire [15-1:0] node4031;
	wire [15-1:0] node4032;
	wire [15-1:0] node4036;
	wire [15-1:0] node4037;
	wire [15-1:0] node4039;
	wire [15-1:0] node4042;
	wire [15-1:0] node4043;
	wire [15-1:0] node4044;
	wire [15-1:0] node4048;
	wire [15-1:0] node4049;
	wire [15-1:0] node4053;
	wire [15-1:0] node4054;
	wire [15-1:0] node4055;
	wire [15-1:0] node4056;
	wire [15-1:0] node4057;
	wire [15-1:0] node4061;
	wire [15-1:0] node4062;
	wire [15-1:0] node4064;
	wire [15-1:0] node4068;
	wire [15-1:0] node4069;
	wire [15-1:0] node4071;
	wire [15-1:0] node4073;
	wire [15-1:0] node4076;
	wire [15-1:0] node4079;
	wire [15-1:0] node4080;
	wire [15-1:0] node4081;
	wire [15-1:0] node4084;
	wire [15-1:0] node4085;
	wire [15-1:0] node4086;
	wire [15-1:0] node4089;
	wire [15-1:0] node4093;
	wire [15-1:0] node4094;
	wire [15-1:0] node4095;
	wire [15-1:0] node4098;
	wire [15-1:0] node4099;
	wire [15-1:0] node4103;
	wire [15-1:0] node4105;
	wire [15-1:0] node4106;
	wire [15-1:0] node4110;
	wire [15-1:0] node4111;
	wire [15-1:0] node4112;
	wire [15-1:0] node4113;
	wire [15-1:0] node4115;
	wire [15-1:0] node4118;
	wire [15-1:0] node4119;
	wire [15-1:0] node4120;
	wire [15-1:0] node4122;
	wire [15-1:0] node4127;
	wire [15-1:0] node4128;
	wire [15-1:0] node4129;
	wire [15-1:0] node4131;
	wire [15-1:0] node4134;
	wire [15-1:0] node4137;
	wire [15-1:0] node4138;
	wire [15-1:0] node4141;
	wire [15-1:0] node4144;
	wire [15-1:0] node4145;
	wire [15-1:0] node4146;
	wire [15-1:0] node4149;
	wire [15-1:0] node4150;
	wire [15-1:0] node4151;
	wire [15-1:0] node4153;
	wire [15-1:0] node4157;
	wire [15-1:0] node4160;
	wire [15-1:0] node4161;
	wire [15-1:0] node4162;
	wire [15-1:0] node4165;
	wire [15-1:0] node4168;
	wire [15-1:0] node4169;
	wire [15-1:0] node4170;
	wire [15-1:0] node4172;
	wire [15-1:0] node4175;
	wire [15-1:0] node4177;
	wire [15-1:0] node4180;
	wire [15-1:0] node4182;
	wire [15-1:0] node4183;
	wire [15-1:0] node4187;
	wire [15-1:0] node4188;
	wire [15-1:0] node4189;
	wire [15-1:0] node4190;
	wire [15-1:0] node4191;
	wire [15-1:0] node4193;
	wire [15-1:0] node4194;
	wire [15-1:0] node4198;
	wire [15-1:0] node4199;
	wire [15-1:0] node4200;
	wire [15-1:0] node4204;
	wire [15-1:0] node4206;
	wire [15-1:0] node4209;
	wire [15-1:0] node4210;
	wire [15-1:0] node4211;
	wire [15-1:0] node4212;
	wire [15-1:0] node4215;
	wire [15-1:0] node4216;
	wire [15-1:0] node4219;
	wire [15-1:0] node4222;
	wire [15-1:0] node4225;
	wire [15-1:0] node4226;
	wire [15-1:0] node4229;
	wire [15-1:0] node4231;
	wire [15-1:0] node4234;
	wire [15-1:0] node4235;
	wire [15-1:0] node4236;
	wire [15-1:0] node4238;
	wire [15-1:0] node4241;
	wire [15-1:0] node4242;
	wire [15-1:0] node4243;
	wire [15-1:0] node4245;
	wire [15-1:0] node4246;
	wire [15-1:0] node4251;
	wire [15-1:0] node4252;
	wire [15-1:0] node4253;
	wire [15-1:0] node4256;
	wire [15-1:0] node4259;
	wire [15-1:0] node4262;
	wire [15-1:0] node4263;
	wire [15-1:0] node4264;
	wire [15-1:0] node4267;
	wire [15-1:0] node4268;
	wire [15-1:0] node4272;
	wire [15-1:0] node4274;
	wire [15-1:0] node4277;
	wire [15-1:0] node4278;
	wire [15-1:0] node4279;
	wire [15-1:0] node4280;
	wire [15-1:0] node4281;
	wire [15-1:0] node4285;
	wire [15-1:0] node4286;
	wire [15-1:0] node4287;
	wire [15-1:0] node4291;
	wire [15-1:0] node4294;
	wire [15-1:0] node4295;
	wire [15-1:0] node4296;
	wire [15-1:0] node4298;
	wire [15-1:0] node4302;
	wire [15-1:0] node4303;
	wire [15-1:0] node4306;
	wire [15-1:0] node4309;
	wire [15-1:0] node4310;
	wire [15-1:0] node4311;
	wire [15-1:0] node4312;
	wire [15-1:0] node4315;
	wire [15-1:0] node4316;
	wire [15-1:0] node4317;
	wire [15-1:0] node4319;
	wire [15-1:0] node4324;
	wire [15-1:0] node4325;
	wire [15-1:0] node4326;
	wire [15-1:0] node4328;
	wire [15-1:0] node4329;
	wire [15-1:0] node4334;
	wire [15-1:0] node4336;
	wire [15-1:0] node4337;
	wire [15-1:0] node4341;
	wire [15-1:0] node4342;
	wire [15-1:0] node4344;
	wire [15-1:0] node4345;
	wire [15-1:0] node4349;
	wire [15-1:0] node4350;
	wire [15-1:0] node4352;
	wire [15-1:0] node4353;
	wire [15-1:0] node4354;
	wire [15-1:0] node4359;
	wire [15-1:0] node4360;
	wire [15-1:0] node4362;
	wire [15-1:0] node4365;
	wire [15-1:0] node4368;
	wire [15-1:0] node4369;
	wire [15-1:0] node4370;
	wire [15-1:0] node4371;
	wire [15-1:0] node4372;
	wire [15-1:0] node4373;
	wire [15-1:0] node4374;
	wire [15-1:0] node4375;
	wire [15-1:0] node4376;
	wire [15-1:0] node4377;
	wire [15-1:0] node4378;
	wire [15-1:0] node4380;
	wire [15-1:0] node4381;
	wire [15-1:0] node4387;
	wire [15-1:0] node4388;
	wire [15-1:0] node4392;
	wire [15-1:0] node4393;
	wire [15-1:0] node4394;
	wire [15-1:0] node4396;
	wire [15-1:0] node4399;
	wire [15-1:0] node4400;
	wire [15-1:0] node4404;
	wire [15-1:0] node4407;
	wire [15-1:0] node4408;
	wire [15-1:0] node4409;
	wire [15-1:0] node4411;
	wire [15-1:0] node4414;
	wire [15-1:0] node4415;
	wire [15-1:0] node4416;
	wire [15-1:0] node4420;
	wire [15-1:0] node4422;
	wire [15-1:0] node4425;
	wire [15-1:0] node4426;
	wire [15-1:0] node4427;
	wire [15-1:0] node4431;
	wire [15-1:0] node4434;
	wire [15-1:0] node4435;
	wire [15-1:0] node4436;
	wire [15-1:0] node4437;
	wire [15-1:0] node4439;
	wire [15-1:0] node4442;
	wire [15-1:0] node4445;
	wire [15-1:0] node4448;
	wire [15-1:0] node4449;
	wire [15-1:0] node4451;
	wire [15-1:0] node4452;
	wire [15-1:0] node4453;
	wire [15-1:0] node4458;
	wire [15-1:0] node4459;
	wire [15-1:0] node4463;
	wire [15-1:0] node4464;
	wire [15-1:0] node4465;
	wire [15-1:0] node4466;
	wire [15-1:0] node4467;
	wire [15-1:0] node4468;
	wire [15-1:0] node4472;
	wire [15-1:0] node4473;
	wire [15-1:0] node4475;
	wire [15-1:0] node4479;
	wire [15-1:0] node4480;
	wire [15-1:0] node4482;
	wire [15-1:0] node4483;
	wire [15-1:0] node4488;
	wire [15-1:0] node4489;
	wire [15-1:0] node4490;
	wire [15-1:0] node4493;
	wire [15-1:0] node4495;
	wire [15-1:0] node4498;
	wire [15-1:0] node4499;
	wire [15-1:0] node4500;
	wire [15-1:0] node4502;
	wire [15-1:0] node4505;
	wire [15-1:0] node4509;
	wire [15-1:0] node4510;
	wire [15-1:0] node4511;
	wire [15-1:0] node4512;
	wire [15-1:0] node4515;
	wire [15-1:0] node4518;
	wire [15-1:0] node4519;
	wire [15-1:0] node4520;
	wire [15-1:0] node4522;
	wire [15-1:0] node4527;
	wire [15-1:0] node4528;
	wire [15-1:0] node4530;
	wire [15-1:0] node4533;
	wire [15-1:0] node4534;
	wire [15-1:0] node4537;
	wire [15-1:0] node4538;
	wire [15-1:0] node4542;
	wire [15-1:0] node4543;
	wire [15-1:0] node4544;
	wire [15-1:0] node4545;
	wire [15-1:0] node4546;
	wire [15-1:0] node4547;
	wire [15-1:0] node4548;
	wire [15-1:0] node4550;
	wire [15-1:0] node4553;
	wire [15-1:0] node4556;
	wire [15-1:0] node4557;
	wire [15-1:0] node4559;
	wire [15-1:0] node4563;
	wire [15-1:0] node4564;
	wire [15-1:0] node4565;
	wire [15-1:0] node4567;
	wire [15-1:0] node4572;
	wire [15-1:0] node4573;
	wire [15-1:0] node4574;
	wire [15-1:0] node4577;
	wire [15-1:0] node4580;
	wire [15-1:0] node4581;
	wire [15-1:0] node4582;
	wire [15-1:0] node4583;
	wire [15-1:0] node4585;
	wire [15-1:0] node4591;
	wire [15-1:0] node4592;
	wire [15-1:0] node4593;
	wire [15-1:0] node4595;
	wire [15-1:0] node4597;
	wire [15-1:0] node4600;
	wire [15-1:0] node4602;
	wire [15-1:0] node4603;
	wire [15-1:0] node4607;
	wire [15-1:0] node4608;
	wire [15-1:0] node4609;
	wire [15-1:0] node4610;
	wire [15-1:0] node4612;
	wire [15-1:0] node4616;
	wire [15-1:0] node4619;
	wire [15-1:0] node4620;
	wire [15-1:0] node4621;
	wire [15-1:0] node4625;
	wire [15-1:0] node4627;
	wire [15-1:0] node4629;
	wire [15-1:0] node4632;
	wire [15-1:0] node4633;
	wire [15-1:0] node4634;
	wire [15-1:0] node4635;
	wire [15-1:0] node4636;
	wire [15-1:0] node4637;
	wire [15-1:0] node4641;
	wire [15-1:0] node4642;
	wire [15-1:0] node4645;
	wire [15-1:0] node4646;
	wire [15-1:0] node4650;
	wire [15-1:0] node4652;
	wire [15-1:0] node4655;
	wire [15-1:0] node4656;
	wire [15-1:0] node4657;
	wire [15-1:0] node4658;
	wire [15-1:0] node4661;
	wire [15-1:0] node4664;
	wire [15-1:0] node4665;
	wire [15-1:0] node4666;
	wire [15-1:0] node4671;
	wire [15-1:0] node4673;
	wire [15-1:0] node4674;
	wire [15-1:0] node4678;
	wire [15-1:0] node4679;
	wire [15-1:0] node4680;
	wire [15-1:0] node4683;
	wire [15-1:0] node4684;
	wire [15-1:0] node4685;
	wire [15-1:0] node4689;
	wire [15-1:0] node4692;
	wire [15-1:0] node4693;
	wire [15-1:0] node4694;
	wire [15-1:0] node4698;
	wire [15-1:0] node4700;
	wire [15-1:0] node4701;
	wire [15-1:0] node4704;
	wire [15-1:0] node4705;
	wire [15-1:0] node4709;
	wire [15-1:0] node4710;
	wire [15-1:0] node4711;
	wire [15-1:0] node4712;
	wire [15-1:0] node4713;
	wire [15-1:0] node4714;
	wire [15-1:0] node4715;
	wire [15-1:0] node4717;
	wire [15-1:0] node4721;
	wire [15-1:0] node4722;
	wire [15-1:0] node4723;
	wire [15-1:0] node4724;
	wire [15-1:0] node4728;
	wire [15-1:0] node4731;
	wire [15-1:0] node4733;
	wire [15-1:0] node4736;
	wire [15-1:0] node4737;
	wire [15-1:0] node4738;
	wire [15-1:0] node4739;
	wire [15-1:0] node4743;
	wire [15-1:0] node4746;
	wire [15-1:0] node4747;
	wire [15-1:0] node4750;
	wire [15-1:0] node4753;
	wire [15-1:0] node4754;
	wire [15-1:0] node4755;
	wire [15-1:0] node4756;
	wire [15-1:0] node4759;
	wire [15-1:0] node4761;
	wire [15-1:0] node4762;
	wire [15-1:0] node4766;
	wire [15-1:0] node4767;
	wire [15-1:0] node4768;
	wire [15-1:0] node4773;
	wire [15-1:0] node4774;
	wire [15-1:0] node4775;
	wire [15-1:0] node4776;
	wire [15-1:0] node4778;
	wire [15-1:0] node4780;
	wire [15-1:0] node4785;
	wire [15-1:0] node4786;
	wire [15-1:0] node4787;
	wire [15-1:0] node4791;
	wire [15-1:0] node4794;
	wire [15-1:0] node4795;
	wire [15-1:0] node4796;
	wire [15-1:0] node4797;
	wire [15-1:0] node4798;
	wire [15-1:0] node4801;
	wire [15-1:0] node4803;
	wire [15-1:0] node4806;
	wire [15-1:0] node4807;
	wire [15-1:0] node4808;
	wire [15-1:0] node4812;
	wire [15-1:0] node4814;
	wire [15-1:0] node4817;
	wire [15-1:0] node4818;
	wire [15-1:0] node4819;
	wire [15-1:0] node4821;
	wire [15-1:0] node4825;
	wire [15-1:0] node4827;
	wire [15-1:0] node4828;
	wire [15-1:0] node4831;
	wire [15-1:0] node4833;
	wire [15-1:0] node4836;
	wire [15-1:0] node4837;
	wire [15-1:0] node4838;
	wire [15-1:0] node4839;
	wire [15-1:0] node4842;
	wire [15-1:0] node4845;
	wire [15-1:0] node4846;
	wire [15-1:0] node4848;
	wire [15-1:0] node4851;
	wire [15-1:0] node4853;
	wire [15-1:0] node4855;
	wire [15-1:0] node4858;
	wire [15-1:0] node4859;
	wire [15-1:0] node4860;
	wire [15-1:0] node4861;
	wire [15-1:0] node4863;
	wire [15-1:0] node4866;
	wire [15-1:0] node4869;
	wire [15-1:0] node4870;
	wire [15-1:0] node4872;
	wire [15-1:0] node4876;
	wire [15-1:0] node4877;
	wire [15-1:0] node4879;
	wire [15-1:0] node4880;
	wire [15-1:0] node4884;
	wire [15-1:0] node4885;
	wire [15-1:0] node4887;
	wire [15-1:0] node4891;
	wire [15-1:0] node4892;
	wire [15-1:0] node4893;
	wire [15-1:0] node4894;
	wire [15-1:0] node4895;
	wire [15-1:0] node4896;
	wire [15-1:0] node4899;
	wire [15-1:0] node4902;
	wire [15-1:0] node4903;
	wire [15-1:0] node4904;
	wire [15-1:0] node4908;
	wire [15-1:0] node4911;
	wire [15-1:0] node4912;
	wire [15-1:0] node4913;
	wire [15-1:0] node4915;
	wire [15-1:0] node4918;
	wire [15-1:0] node4920;
	wire [15-1:0] node4923;
	wire [15-1:0] node4924;
	wire [15-1:0] node4925;
	wire [15-1:0] node4930;
	wire [15-1:0] node4931;
	wire [15-1:0] node4932;
	wire [15-1:0] node4934;
	wire [15-1:0] node4935;
	wire [15-1:0] node4939;
	wire [15-1:0] node4940;
	wire [15-1:0] node4942;
	wire [15-1:0] node4945;
	wire [15-1:0] node4948;
	wire [15-1:0] node4949;
	wire [15-1:0] node4950;
	wire [15-1:0] node4951;
	wire [15-1:0] node4953;
	wire [15-1:0] node4957;
	wire [15-1:0] node4958;
	wire [15-1:0] node4960;
	wire [15-1:0] node4963;
	wire [15-1:0] node4964;
	wire [15-1:0] node4968;
	wire [15-1:0] node4969;
	wire [15-1:0] node4971;
	wire [15-1:0] node4974;
	wire [15-1:0] node4976;
	wire [15-1:0] node4977;
	wire [15-1:0] node4981;
	wire [15-1:0] node4982;
	wire [15-1:0] node4983;
	wire [15-1:0] node4984;
	wire [15-1:0] node4985;
	wire [15-1:0] node4986;
	wire [15-1:0] node4990;
	wire [15-1:0] node4991;
	wire [15-1:0] node4994;
	wire [15-1:0] node4996;
	wire [15-1:0] node4999;
	wire [15-1:0] node5000;
	wire [15-1:0] node5003;
	wire [15-1:0] node5006;
	wire [15-1:0] node5007;
	wire [15-1:0] node5008;
	wire [15-1:0] node5011;
	wire [15-1:0] node5014;
	wire [15-1:0] node5015;
	wire [15-1:0] node5016;
	wire [15-1:0] node5020;
	wire [15-1:0] node5023;
	wire [15-1:0] node5024;
	wire [15-1:0] node5025;
	wire [15-1:0] node5026;
	wire [15-1:0] node5029;
	wire [15-1:0] node5030;
	wire [15-1:0] node5032;
	wire [15-1:0] node5036;
	wire [15-1:0] node5037;
	wire [15-1:0] node5041;
	wire [15-1:0] node5042;
	wire [15-1:0] node5043;
	wire [15-1:0] node5045;
	wire [15-1:0] node5048;
	wire [15-1:0] node5050;
	wire [15-1:0] node5051;
	wire [15-1:0] node5053;
	wire [15-1:0] node5057;
	wire [15-1:0] node5058;
	wire [15-1:0] node5060;
	wire [15-1:0] node5061;
	wire [15-1:0] node5065;
	wire [15-1:0] node5066;
	wire [15-1:0] node5068;
	wire [15-1:0] node5072;
	wire [15-1:0] node5073;
	wire [15-1:0] node5074;
	wire [15-1:0] node5075;
	wire [15-1:0] node5076;
	wire [15-1:0] node5077;
	wire [15-1:0] node5078;
	wire [15-1:0] node5079;
	wire [15-1:0] node5080;
	wire [15-1:0] node5081;
	wire [15-1:0] node5085;
	wire [15-1:0] node5089;
	wire [15-1:0] node5090;
	wire [15-1:0] node5091;
	wire [15-1:0] node5095;
	wire [15-1:0] node5097;
	wire [15-1:0] node5098;
	wire [15-1:0] node5102;
	wire [15-1:0] node5103;
	wire [15-1:0] node5104;
	wire [15-1:0] node5106;
	wire [15-1:0] node5109;
	wire [15-1:0] node5110;
	wire [15-1:0] node5111;
	wire [15-1:0] node5116;
	wire [15-1:0] node5117;
	wire [15-1:0] node5120;
	wire [15-1:0] node5121;
	wire [15-1:0] node5123;
	wire [15-1:0] node5127;
	wire [15-1:0] node5128;
	wire [15-1:0] node5129;
	wire [15-1:0] node5130;
	wire [15-1:0] node5133;
	wire [15-1:0] node5135;
	wire [15-1:0] node5138;
	wire [15-1:0] node5139;
	wire [15-1:0] node5140;
	wire [15-1:0] node5144;
	wire [15-1:0] node5146;
	wire [15-1:0] node5148;
	wire [15-1:0] node5151;
	wire [15-1:0] node5152;
	wire [15-1:0] node5153;
	wire [15-1:0] node5156;
	wire [15-1:0] node5157;
	wire [15-1:0] node5159;
	wire [15-1:0] node5163;
	wire [15-1:0] node5164;
	wire [15-1:0] node5167;
	wire [15-1:0] node5170;
	wire [15-1:0] node5171;
	wire [15-1:0] node5172;
	wire [15-1:0] node5173;
	wire [15-1:0] node5174;
	wire [15-1:0] node5175;
	wire [15-1:0] node5179;
	wire [15-1:0] node5182;
	wire [15-1:0] node5183;
	wire [15-1:0] node5186;
	wire [15-1:0] node5187;
	wire [15-1:0] node5189;
	wire [15-1:0] node5193;
	wire [15-1:0] node5195;
	wire [15-1:0] node5196;
	wire [15-1:0] node5197;
	wire [15-1:0] node5198;
	wire [15-1:0] node5202;
	wire [15-1:0] node5205;
	wire [15-1:0] node5206;
	wire [15-1:0] node5210;
	wire [15-1:0] node5211;
	wire [15-1:0] node5212;
	wire [15-1:0] node5213;
	wire [15-1:0] node5214;
	wire [15-1:0] node5216;
	wire [15-1:0] node5220;
	wire [15-1:0] node5222;
	wire [15-1:0] node5223;
	wire [15-1:0] node5227;
	wire [15-1:0] node5228;
	wire [15-1:0] node5229;
	wire [15-1:0] node5230;
	wire [15-1:0] node5234;
	wire [15-1:0] node5236;
	wire [15-1:0] node5239;
	wire [15-1:0] node5240;
	wire [15-1:0] node5244;
	wire [15-1:0] node5245;
	wire [15-1:0] node5246;
	wire [15-1:0] node5248;
	wire [15-1:0] node5251;
	wire [15-1:0] node5253;
	wire [15-1:0] node5256;
	wire [15-1:0] node5257;
	wire [15-1:0] node5258;
	wire [15-1:0] node5262;
	wire [15-1:0] node5263;
	wire [15-1:0] node5265;
	wire [15-1:0] node5268;
	wire [15-1:0] node5269;
	wire [15-1:0] node5270;
	wire [15-1:0] node5272;
	wire [15-1:0] node5277;
	wire [15-1:0] node5278;
	wire [15-1:0] node5279;
	wire [15-1:0] node5280;
	wire [15-1:0] node5281;
	wire [15-1:0] node5283;
	wire [15-1:0] node5284;
	wire [15-1:0] node5288;
	wire [15-1:0] node5289;
	wire [15-1:0] node5292;
	wire [15-1:0] node5295;
	wire [15-1:0] node5296;
	wire [15-1:0] node5297;
	wire [15-1:0] node5298;
	wire [15-1:0] node5301;
	wire [15-1:0] node5304;
	wire [15-1:0] node5307;
	wire [15-1:0] node5308;
	wire [15-1:0] node5311;
	wire [15-1:0] node5312;
	wire [15-1:0] node5315;
	wire [15-1:0] node5317;
	wire [15-1:0] node5320;
	wire [15-1:0] node5321;
	wire [15-1:0] node5323;
	wire [15-1:0] node5324;
	wire [15-1:0] node5325;
	wire [15-1:0] node5326;
	wire [15-1:0] node5329;
	wire [15-1:0] node5331;
	wire [15-1:0] node5335;
	wire [15-1:0] node5338;
	wire [15-1:0] node5339;
	wire [15-1:0] node5340;
	wire [15-1:0] node5344;
	wire [15-1:0] node5346;
	wire [15-1:0] node5349;
	wire [15-1:0] node5350;
	wire [15-1:0] node5351;
	wire [15-1:0] node5352;
	wire [15-1:0] node5353;
	wire [15-1:0] node5356;
	wire [15-1:0] node5358;
	wire [15-1:0] node5359;
	wire [15-1:0] node5363;
	wire [15-1:0] node5364;
	wire [15-1:0] node5365;
	wire [15-1:0] node5369;
	wire [15-1:0] node5371;
	wire [15-1:0] node5373;
	wire [15-1:0] node5376;
	wire [15-1:0] node5377;
	wire [15-1:0] node5378;
	wire [15-1:0] node5381;
	wire [15-1:0] node5382;
	wire [15-1:0] node5384;
	wire [15-1:0] node5387;
	wire [15-1:0] node5389;
	wire [15-1:0] node5392;
	wire [15-1:0] node5394;
	wire [15-1:0] node5397;
	wire [15-1:0] node5398;
	wire [15-1:0] node5399;
	wire [15-1:0] node5400;
	wire [15-1:0] node5401;
	wire [15-1:0] node5405;
	wire [15-1:0] node5407;
	wire [15-1:0] node5410;
	wire [15-1:0] node5411;
	wire [15-1:0] node5414;
	wire [15-1:0] node5417;
	wire [15-1:0] node5418;
	wire [15-1:0] node5420;
	wire [15-1:0] node5422;
	wire [15-1:0] node5425;
	wire [15-1:0] node5426;
	wire [15-1:0] node5429;
	wire [15-1:0] node5430;
	wire [15-1:0] node5432;
	wire [15-1:0] node5436;
	wire [15-1:0] node5437;
	wire [15-1:0] node5438;
	wire [15-1:0] node5439;
	wire [15-1:0] node5440;
	wire [15-1:0] node5441;
	wire [15-1:0] node5442;
	wire [15-1:0] node5444;
	wire [15-1:0] node5448;
	wire [15-1:0] node5449;
	wire [15-1:0] node5450;
	wire [15-1:0] node5452;
	wire [15-1:0] node5456;
	wire [15-1:0] node5458;
	wire [15-1:0] node5461;
	wire [15-1:0] node5462;
	wire [15-1:0] node5463;
	wire [15-1:0] node5466;
	wire [15-1:0] node5468;
	wire [15-1:0] node5471;
	wire [15-1:0] node5473;
	wire [15-1:0] node5476;
	wire [15-1:0] node5477;
	wire [15-1:0] node5478;
	wire [15-1:0] node5480;
	wire [15-1:0] node5483;
	wire [15-1:0] node5485;
	wire [15-1:0] node5488;
	wire [15-1:0] node5489;
	wire [15-1:0] node5490;
	wire [15-1:0] node5491;
	wire [15-1:0] node5494;
	wire [15-1:0] node5497;
	wire [15-1:0] node5498;
	wire [15-1:0] node5500;
	wire [15-1:0] node5503;
	wire [15-1:0] node5504;
	wire [15-1:0] node5505;
	wire [15-1:0] node5510;
	wire [15-1:0] node5511;
	wire [15-1:0] node5512;
	wire [15-1:0] node5514;
	wire [15-1:0] node5516;
	wire [15-1:0] node5520;
	wire [15-1:0] node5521;
	wire [15-1:0] node5525;
	wire [15-1:0] node5526;
	wire [15-1:0] node5527;
	wire [15-1:0] node5528;
	wire [15-1:0] node5530;
	wire [15-1:0] node5531;
	wire [15-1:0] node5533;
	wire [15-1:0] node5536;
	wire [15-1:0] node5537;
	wire [15-1:0] node5538;
	wire [15-1:0] node5543;
	wire [15-1:0] node5544;
	wire [15-1:0] node5548;
	wire [15-1:0] node5549;
	wire [15-1:0] node5550;
	wire [15-1:0] node5553;
	wire [15-1:0] node5555;
	wire [15-1:0] node5558;
	wire [15-1:0] node5559;
	wire [15-1:0] node5562;
	wire [15-1:0] node5563;
	wire [15-1:0] node5564;
	wire [15-1:0] node5569;
	wire [15-1:0] node5570;
	wire [15-1:0] node5571;
	wire [15-1:0] node5572;
	wire [15-1:0] node5575;
	wire [15-1:0] node5577;
	wire [15-1:0] node5578;
	wire [15-1:0] node5582;
	wire [15-1:0] node5583;
	wire [15-1:0] node5586;
	wire [15-1:0] node5587;
	wire [15-1:0] node5588;
	wire [15-1:0] node5593;
	wire [15-1:0] node5594;
	wire [15-1:0] node5595;
	wire [15-1:0] node5597;
	wire [15-1:0] node5599;
	wire [15-1:0] node5602;
	wire [15-1:0] node5603;
	wire [15-1:0] node5605;
	wire [15-1:0] node5608;
	wire [15-1:0] node5611;
	wire [15-1:0] node5613;
	wire [15-1:0] node5615;
	wire [15-1:0] node5618;
	wire [15-1:0] node5619;
	wire [15-1:0] node5620;
	wire [15-1:0] node5621;
	wire [15-1:0] node5622;
	wire [15-1:0] node5623;
	wire [15-1:0] node5625;
	wire [15-1:0] node5626;
	wire [15-1:0] node5627;
	wire [15-1:0] node5632;
	wire [15-1:0] node5635;
	wire [15-1:0] node5636;
	wire [15-1:0] node5639;
	wire [15-1:0] node5640;
	wire [15-1:0] node5642;
	wire [15-1:0] node5646;
	wire [15-1:0] node5647;
	wire [15-1:0] node5649;
	wire [15-1:0] node5652;
	wire [15-1:0] node5653;
	wire [15-1:0] node5655;
	wire [15-1:0] node5658;
	wire [15-1:0] node5659;
	wire [15-1:0] node5662;
	wire [15-1:0] node5665;
	wire [15-1:0] node5666;
	wire [15-1:0] node5667;
	wire [15-1:0] node5668;
	wire [15-1:0] node5669;
	wire [15-1:0] node5670;
	wire [15-1:0] node5672;
	wire [15-1:0] node5677;
	wire [15-1:0] node5679;
	wire [15-1:0] node5680;
	wire [15-1:0] node5684;
	wire [15-1:0] node5685;
	wire [15-1:0] node5687;
	wire [15-1:0] node5689;
	wire [15-1:0] node5690;
	wire [15-1:0] node5691;
	wire [15-1:0] node5696;
	wire [15-1:0] node5698;
	wire [15-1:0] node5700;
	wire [15-1:0] node5703;
	wire [15-1:0] node5704;
	wire [15-1:0] node5705;
	wire [15-1:0] node5706;
	wire [15-1:0] node5708;
	wire [15-1:0] node5712;
	wire [15-1:0] node5713;
	wire [15-1:0] node5715;
	wire [15-1:0] node5719;
	wire [15-1:0] node5720;
	wire [15-1:0] node5721;
	wire [15-1:0] node5725;
	wire [15-1:0] node5728;
	wire [15-1:0] node5729;
	wire [15-1:0] node5730;
	wire [15-1:0] node5731;
	wire [15-1:0] node5733;
	wire [15-1:0] node5736;
	wire [15-1:0] node5737;
	wire [15-1:0] node5738;
	wire [15-1:0] node5740;
	wire [15-1:0] node5744;
	wire [15-1:0] node5746;
	wire [15-1:0] node5749;
	wire [15-1:0] node5750;
	wire [15-1:0] node5751;
	wire [15-1:0] node5754;
	wire [15-1:0] node5755;
	wire [15-1:0] node5756;
	wire [15-1:0] node5757;
	wire [15-1:0] node5761;
	wire [15-1:0] node5764;
	wire [15-1:0] node5766;
	wire [15-1:0] node5769;
	wire [15-1:0] node5770;
	wire [15-1:0] node5772;
	wire [15-1:0] node5774;
	wire [15-1:0] node5778;
	wire [15-1:0] node5779;
	wire [15-1:0] node5780;
	wire [15-1:0] node5781;
	wire [15-1:0] node5784;
	wire [15-1:0] node5786;
	wire [15-1:0] node5789;
	wire [15-1:0] node5790;
	wire [15-1:0] node5792;
	wire [15-1:0] node5795;
	wire [15-1:0] node5796;
	wire [15-1:0] node5798;
	wire [15-1:0] node5802;
	wire [15-1:0] node5803;
	wire [15-1:0] node5804;
	wire [15-1:0] node5806;
	wire [15-1:0] node5809;
	wire [15-1:0] node5810;
	wire [15-1:0] node5814;
	wire [15-1:0] node5815;
	wire [15-1:0] node5816;
	wire [15-1:0] node5820;
	wire [15-1:0] node5822;
	wire [15-1:0] node5823;
	wire [15-1:0] node5825;

	assign outp = (inp[12]) ? node2916 : node1;
		assign node1 = (inp[10]) ? node1473 : node2;
			assign node2 = (inp[5]) ? node780 : node3;
				assign node3 = (inp[2]) ? node385 : node4;
					assign node4 = (inp[6]) ? node206 : node5;
						assign node5 = (inp[1]) ? node111 : node6;
							assign node6 = (inp[0]) ? node66 : node7;
								assign node7 = (inp[14]) ? node47 : node8;
									assign node8 = (inp[8]) ? node26 : node9;
										assign node9 = (inp[9]) ? node17 : node10;
											assign node10 = (inp[11]) ? 15'b001111111111111 : node11;
												assign node11 = (inp[4]) ? 15'b001111111111111 : node12;
													assign node12 = (inp[13]) ? 15'b001111111111111 : 15'b011111111111111;
											assign node17 = (inp[7]) ? node19 : 15'b001111111111111;
												assign node19 = (inp[4]) ? node21 : 15'b000111111111111;
													assign node21 = (inp[13]) ? 15'b000011111111111 : node22;
														assign node22 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node26 = (inp[7]) ? node42 : node27;
											assign node27 = (inp[4]) ? node35 : node28;
												assign node28 = (inp[11]) ? 15'b001111111111111 : node29;
													assign node29 = (inp[9]) ? 15'b000111111111111 : node30;
														assign node30 = (inp[3]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node35 = (inp[9]) ? 15'b000000111111111 : node36;
													assign node36 = (inp[3]) ? 15'b000011111111111 : node37;
														assign node37 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node42 = (inp[3]) ? node44 : 15'b000011111111111;
												assign node44 = (inp[11]) ? 15'b000011111111111 : 15'b000001111111111;
									assign node47 = (inp[11]) ? node57 : node48;
										assign node48 = (inp[7]) ? node50 : 15'b000111111111111;
											assign node50 = (inp[13]) ? node54 : node51;
												assign node51 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node54 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node57 = (inp[8]) ? node59 : 15'b000011111111111;
											assign node59 = (inp[3]) ? node61 : 15'b000001111111111;
												assign node61 = (inp[4]) ? 15'b000000111111111 : node62;
													assign node62 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
								assign node66 = (inp[8]) ? node82 : node67;
									assign node67 = (inp[13]) ? node73 : node68;
										assign node68 = (inp[3]) ? node70 : 15'b000111111111111;
											assign node70 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node73 = (inp[4]) ? node77 : node74;
											assign node74 = (inp[9]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node77 = (inp[14]) ? node79 : 15'b000001111111111;
												assign node79 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node82 = (inp[7]) ? node98 : node83;
										assign node83 = (inp[14]) ? node93 : node84;
											assign node84 = (inp[4]) ? node90 : node85;
												assign node85 = (inp[11]) ? 15'b000011111111111 : node86;
													assign node86 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node90 = (inp[9]) ? 15'b000000111111111 : 15'b000011111111111;
											assign node93 = (inp[4]) ? node95 : 15'b000001111111111;
												assign node95 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node98 = (inp[11]) ? node104 : node99;
											assign node99 = (inp[14]) ? 15'b000000111111111 : node100;
												assign node100 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node104 = (inp[14]) ? 15'b000000011111111 : node105;
												assign node105 = (inp[9]) ? node107 : 15'b000001111111111;
													assign node107 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node111 = (inp[8]) ? node171 : node112;
								assign node112 = (inp[11]) ? node146 : node113;
									assign node113 = (inp[7]) ? node129 : node114;
										assign node114 = (inp[4]) ? node122 : node115;
											assign node115 = (inp[13]) ? 15'b000011111111111 : node116;
												assign node116 = (inp[3]) ? node118 : 15'b000111111111111;
													assign node118 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node122 = (inp[13]) ? node124 : 15'b000011111111111;
												assign node124 = (inp[0]) ? 15'b000001111111111 : node125;
													assign node125 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node129 = (inp[3]) ? node139 : node130;
											assign node130 = (inp[4]) ? node132 : 15'b000011111111111;
												assign node132 = (inp[13]) ? node136 : node133;
													assign node133 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node136 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node139 = (inp[13]) ? node143 : node140;
												assign node140 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node143 = (inp[4]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node146 = (inp[9]) ? node158 : node147;
										assign node147 = (inp[3]) ? node153 : node148;
											assign node148 = (inp[14]) ? node150 : 15'b000011111111111;
												assign node150 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node153 = (inp[7]) ? node155 : 15'b000001111111111;
												assign node155 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node158 = (inp[13]) ? node162 : node159;
											assign node159 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node162 = (inp[3]) ? node168 : node163;
												assign node163 = (inp[4]) ? node165 : 15'b000000111111111;
													assign node165 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node168 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node171 = (inp[0]) ? node191 : node172;
									assign node172 = (inp[9]) ? node184 : node173;
										assign node173 = (inp[4]) ? node179 : node174;
											assign node174 = (inp[7]) ? node176 : 15'b001111111111111;
												assign node176 = (inp[11]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node179 = (inp[14]) ? 15'b000001111111111 : node180;
												assign node180 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node184 = (inp[14]) ? 15'b000000011111111 : node185;
											assign node185 = (inp[13]) ? node187 : 15'b000000111111111;
												assign node187 = (inp[11]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node191 = (inp[4]) ? node197 : node192;
										assign node192 = (inp[13]) ? 15'b000000011111111 : node193;
											assign node193 = (inp[9]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node197 = (inp[11]) ? node201 : node198;
											assign node198 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node201 = (inp[13]) ? 15'b000000000111111 : node202;
												assign node202 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node206 = (inp[0]) ? node296 : node207;
							assign node207 = (inp[4]) ? node253 : node208;
								assign node208 = (inp[7]) ? node228 : node209;
									assign node209 = (inp[9]) ? node217 : node210;
										assign node210 = (inp[14]) ? 15'b000011111111111 : node211;
											assign node211 = (inp[11]) ? 15'b000011111111111 : node212;
												assign node212 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node217 = (inp[14]) ? 15'b000001111111111 : node218;
											assign node218 = (inp[3]) ? node222 : node219;
												assign node219 = (inp[1]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node222 = (inp[13]) ? 15'b000001111111111 : node223;
													assign node223 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node228 = (inp[14]) ? node242 : node229;
										assign node229 = (inp[9]) ? node233 : node230;
											assign node230 = (inp[1]) ? 15'b000001111111111 : 15'b000111111111111;
											assign node233 = (inp[13]) ? node239 : node234;
												assign node234 = (inp[1]) ? 15'b000001111111111 : node235;
													assign node235 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node239 = (inp[11]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node242 = (inp[11]) ? node246 : node243;
											assign node243 = (inp[13]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node246 = (inp[3]) ? node248 : 15'b000000111111111;
												assign node248 = (inp[9]) ? node250 : 15'b000000011111111;
													assign node250 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node253 = (inp[13]) ? node275 : node254;
									assign node254 = (inp[14]) ? node262 : node255;
										assign node255 = (inp[8]) ? 15'b000001111111111 : node256;
											assign node256 = (inp[1]) ? node258 : 15'b001111111111111;
												assign node258 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node262 = (inp[1]) ? node264 : 15'b000001111111111;
											assign node264 = (inp[8]) ? node272 : node265;
												assign node265 = (inp[3]) ? node267 : 15'b000000111111111;
													assign node267 = (inp[9]) ? 15'b000000011111111 : node268;
														assign node268 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node272 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node275 = (inp[1]) ? node283 : node276;
										assign node276 = (inp[11]) ? node280 : node277;
											assign node277 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node280 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node283 = (inp[14]) ? node291 : node284;
											assign node284 = (inp[3]) ? 15'b000000011111111 : node285;
												assign node285 = (inp[8]) ? 15'b000000011111111 : node286;
													assign node286 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node291 = (inp[7]) ? node293 : 15'b000000011111111;
												assign node293 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node296 = (inp[9]) ? node350 : node297;
								assign node297 = (inp[1]) ? node329 : node298;
									assign node298 = (inp[7]) ? node320 : node299;
										assign node299 = (inp[13]) ? node307 : node300;
											assign node300 = (inp[3]) ? node302 : 15'b000000111111111;
												assign node302 = (inp[14]) ? 15'b000001111111111 : node303;
													assign node303 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node307 = (inp[3]) ? node313 : node308;
												assign node308 = (inp[4]) ? node310 : 15'b000001111111111;
													assign node310 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node313 = (inp[8]) ? 15'b000000011111111 : node314;
													assign node314 = (inp[14]) ? 15'b000000111111111 : node315;
														assign node315 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node320 = (inp[3]) ? node326 : node321;
											assign node321 = (inp[14]) ? 15'b000000111111111 : node322;
												assign node322 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node326 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node329 = (inp[3]) ? node337 : node330;
										assign node330 = (inp[14]) ? node334 : node331;
											assign node331 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node334 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node337 = (inp[11]) ? node347 : node338;
											assign node338 = (inp[8]) ? node342 : node339;
												assign node339 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node342 = (inp[4]) ? node344 : 15'b000000111111111;
													assign node344 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node347 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
								assign node350 = (inp[3]) ? node370 : node351;
									assign node351 = (inp[8]) ? node357 : node352;
										assign node352 = (inp[13]) ? node354 : 15'b000001111111111;
											assign node354 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node357 = (inp[4]) ? node363 : node358;
											assign node358 = (inp[11]) ? 15'b000000011111111 : node359;
												assign node359 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node363 = (inp[7]) ? node365 : 15'b000000011111111;
												assign node365 = (inp[11]) ? 15'b000000001111111 : node366;
													assign node366 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node370 = (inp[14]) ? node378 : node371;
										assign node371 = (inp[8]) ? node375 : node372;
											assign node372 = (inp[4]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node375 = (inp[4]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node378 = (inp[7]) ? node382 : node379;
											assign node379 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node382 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node385 = (inp[3]) ? node557 : node386;
						assign node386 = (inp[13]) ? node464 : node387;
							assign node387 = (inp[6]) ? node431 : node388;
								assign node388 = (inp[1]) ? node400 : node389;
									assign node389 = (inp[9]) ? node395 : node390;
										assign node390 = (inp[4]) ? 15'b000011111111111 : node391;
											assign node391 = (inp[14]) ? 15'b000111111111111 : 15'b011111111111111;
										assign node395 = (inp[14]) ? 15'b000001111111111 : node396;
											assign node396 = (inp[11]) ? 15'b000001111111111 : 15'b000111111111111;
									assign node400 = (inp[9]) ? node414 : node401;
										assign node401 = (inp[14]) ? node411 : node402;
											assign node402 = (inp[11]) ? node408 : node403;
												assign node403 = (inp[8]) ? 15'b000011111111111 : node404;
													assign node404 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node408 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node411 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node414 = (inp[0]) ? node428 : node415;
											assign node415 = (inp[8]) ? node423 : node416;
												assign node416 = (inp[11]) ? 15'b000001111111111 : node417;
													assign node417 = (inp[4]) ? node419 : 15'b000011111111111;
														assign node419 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node423 = (inp[7]) ? 15'b000000011111111 : node424;
													assign node424 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node428 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node431 = (inp[8]) ? node455 : node432;
									assign node432 = (inp[14]) ? node442 : node433;
										assign node433 = (inp[1]) ? node437 : node434;
											assign node434 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node437 = (inp[0]) ? node439 : 15'b000001111111111;
												assign node439 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node442 = (inp[0]) ? node450 : node443;
											assign node443 = (inp[4]) ? node445 : 15'b000001111111111;
												assign node445 = (inp[1]) ? 15'b000000011111111 : node446;
													assign node446 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node450 = (inp[7]) ? 15'b000000011111111 : node451;
												assign node451 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node455 = (inp[7]) ? node457 : 15'b000000111111111;
										assign node457 = (inp[9]) ? node459 : 15'b000000011111111;
											assign node459 = (inp[4]) ? 15'b000000000111111 : node460;
												assign node460 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node464 = (inp[0]) ? node514 : node465;
								assign node465 = (inp[9]) ? node487 : node466;
									assign node466 = (inp[11]) ? node480 : node467;
										assign node467 = (inp[14]) ? node473 : node468;
											assign node468 = (inp[4]) ? node470 : 15'b000011111111111;
												assign node470 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node473 = (inp[6]) ? 15'b000000111111111 : node474;
												assign node474 = (inp[1]) ? node476 : 15'b000001111111111;
													assign node476 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node480 = (inp[4]) ? 15'b000000111111111 : node481;
											assign node481 = (inp[1]) ? 15'b000000011111111 : node482;
												assign node482 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node487 = (inp[6]) ? node501 : node488;
										assign node488 = (inp[7]) ? node498 : node489;
											assign node489 = (inp[14]) ? 15'b000000111111111 : node490;
												assign node490 = (inp[8]) ? 15'b000000111111111 : node491;
													assign node491 = (inp[11]) ? node493 : 15'b000001111111111;
														assign node493 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node498 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node501 = (inp[11]) ? node507 : node502;
											assign node502 = (inp[4]) ? 15'b000000011111111 : node503;
												assign node503 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node507 = (inp[1]) ? node509 : 15'b000000011111111;
												assign node509 = (inp[4]) ? node511 : 15'b000000001111111;
													assign node511 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node514 = (inp[4]) ? node544 : node515;
									assign node515 = (inp[6]) ? node527 : node516;
										assign node516 = (inp[11]) ? node524 : node517;
											assign node517 = (inp[14]) ? node521 : node518;
												assign node518 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node521 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node524 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node527 = (inp[9]) ? node537 : node528;
											assign node528 = (inp[11]) ? node530 : 15'b000000111111111;
												assign node530 = (inp[7]) ? 15'b000000011111111 : node531;
													assign node531 = (inp[14]) ? 15'b000000011111111 : node532;
														assign node532 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node537 = (inp[8]) ? node541 : node538;
												assign node538 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node541 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node544 = (inp[11]) ? node550 : node545;
										assign node545 = (inp[8]) ? node547 : 15'b000000011111111;
											assign node547 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node550 = (inp[7]) ? node554 : node551;
											assign node551 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node554 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node557 = (inp[13]) ? node647 : node558;
							assign node558 = (inp[8]) ? node594 : node559;
								assign node559 = (inp[4]) ? node579 : node560;
									assign node560 = (inp[0]) ? node568 : node561;
										assign node561 = (inp[1]) ? 15'b000001111111111 : node562;
											assign node562 = (inp[7]) ? node564 : 15'b000111111111111;
												assign node564 = (inp[11]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node568 = (inp[14]) ? node574 : node569;
											assign node569 = (inp[7]) ? 15'b000000111111111 : node570;
												assign node570 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node574 = (inp[7]) ? node576 : 15'b000000111111111;
												assign node576 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node579 = (inp[0]) ? node585 : node580;
										assign node580 = (inp[14]) ? 15'b000000011111111 : node581;
											assign node581 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node585 = (inp[1]) ? node589 : node586;
											assign node586 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node589 = (inp[9]) ? 15'b000000011111111 : node590;
												assign node590 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node594 = (inp[0]) ? node626 : node595;
									assign node595 = (inp[1]) ? node613 : node596;
										assign node596 = (inp[4]) ? node606 : node597;
											assign node597 = (inp[6]) ? node601 : node598;
												assign node598 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node601 = (inp[14]) ? node603 : 15'b000000111111111;
													assign node603 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node606 = (inp[7]) ? 15'b000000011111111 : node607;
												assign node607 = (inp[14]) ? node609 : 15'b000001111111111;
													assign node609 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node613 = (inp[6]) ? node623 : node614;
											assign node614 = (inp[7]) ? 15'b000000011111111 : node615;
												assign node615 = (inp[11]) ? node617 : 15'b000000111111111;
													assign node617 = (inp[4]) ? 15'b000000011111111 : node618;
														assign node618 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node623 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node626 = (inp[11]) ? node636 : node627;
										assign node627 = (inp[1]) ? node633 : node628;
											assign node628 = (inp[7]) ? 15'b000000011111111 : node629;
												assign node629 = (inp[9]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node633 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node636 = (inp[4]) ? node640 : node637;
											assign node637 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node640 = (inp[9]) ? node644 : node641;
												assign node641 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node644 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node647 = (inp[6]) ? node709 : node648;
								assign node648 = (inp[11]) ? node680 : node649;
									assign node649 = (inp[0]) ? node665 : node650;
										assign node650 = (inp[1]) ? 15'b000000111111111 : node651;
											assign node651 = (inp[9]) ? node657 : node652;
												assign node652 = (inp[8]) ? node654 : 15'b000011111111111;
													assign node654 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node657 = (inp[4]) ? node659 : 15'b000001111111111;
													assign node659 = (inp[14]) ? node661 : 15'b000000111111111;
														assign node661 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node665 = (inp[4]) ? node675 : node666;
											assign node666 = (inp[1]) ? node670 : node667;
												assign node667 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node670 = (inp[8]) ? node672 : 15'b000000011111111;
													assign node672 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node675 = (inp[7]) ? 15'b000000011111111 : node676;
												assign node676 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node680 = (inp[14]) ? node698 : node681;
										assign node681 = (inp[7]) ? node693 : node682;
											assign node682 = (inp[9]) ? node690 : node683;
												assign node683 = (inp[4]) ? 15'b000000111111111 : node684;
													assign node684 = (inp[1]) ? node686 : 15'b000001111111111;
														assign node686 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node690 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node693 = (inp[9]) ? node695 : 15'b000000011111111;
												assign node695 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node698 = (inp[0]) ? node704 : node699;
											assign node699 = (inp[7]) ? node701 : 15'b000000011111111;
												assign node701 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node704 = (inp[4]) ? node706 : 15'b000000000111111;
												assign node706 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node709 = (inp[4]) ? node747 : node710;
									assign node710 = (inp[1]) ? node728 : node711;
										assign node711 = (inp[11]) ? node721 : node712;
											assign node712 = (inp[0]) ? 15'b000000011111111 : node713;
												assign node713 = (inp[14]) ? node717 : node714;
													assign node714 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node717 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node721 = (inp[0]) ? 15'b000000001111111 : node722;
												assign node722 = (inp[7]) ? node724 : 15'b000000011111111;
													assign node724 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node728 = (inp[14]) ? node736 : node729;
											assign node729 = (inp[7]) ? 15'b000000001111111 : node730;
												assign node730 = (inp[11]) ? 15'b000000001111111 : node731;
													assign node731 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node736 = (inp[8]) ? node740 : node737;
												assign node737 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node740 = (inp[0]) ? 15'b000000000111111 : node741;
													assign node741 = (inp[7]) ? node743 : 15'b000000011111111;
														assign node743 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node747 = (inp[11]) ? node767 : node748;
										assign node748 = (inp[8]) ? node760 : node749;
											assign node749 = (inp[9]) ? node755 : node750;
												assign node750 = (inp[14]) ? node752 : 15'b000000011111111;
													assign node752 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node755 = (inp[1]) ? node757 : 15'b000000011111111;
													assign node757 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node760 = (inp[14]) ? node762 : 15'b000000001111111;
												assign node762 = (inp[9]) ? 15'b000000000011111 : node763;
													assign node763 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node767 = (inp[7]) ? node775 : node768;
											assign node768 = (inp[9]) ? 15'b000000000111111 : node769;
												assign node769 = (inp[0]) ? node771 : 15'b000000001111111;
													assign node771 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node775 = (inp[9]) ? 15'b000000000011111 : node776;
												assign node776 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
				assign node780 = (inp[8]) ? node1132 : node781;
					assign node781 = (inp[14]) ? node959 : node782;
						assign node782 = (inp[3]) ? node870 : node783;
							assign node783 = (inp[7]) ? node825 : node784;
								assign node784 = (inp[13]) ? node810 : node785;
									assign node785 = (inp[11]) ? node803 : node786;
										assign node786 = (inp[0]) ? node798 : node787;
											assign node787 = (inp[6]) ? node793 : node788;
												assign node788 = (inp[4]) ? 15'b000111111111111 : node789;
													assign node789 = (inp[9]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node793 = (inp[2]) ? 15'b000001111111111 : node794;
													assign node794 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node798 = (inp[2]) ? node800 : 15'b000011111111111;
												assign node800 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node803 = (inp[2]) ? node805 : 15'b000011111111111;
											assign node805 = (inp[4]) ? node807 : 15'b000001111111111;
												assign node807 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
									assign node810 = (inp[2]) ? node816 : node811;
										assign node811 = (inp[1]) ? node813 : 15'b000001111111111;
											assign node813 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node816 = (inp[4]) ? 15'b000000111111111 : node817;
											assign node817 = (inp[6]) ? 15'b000000011111111 : node818;
												assign node818 = (inp[1]) ? 15'b000001111111111 : node819;
													assign node819 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
								assign node825 = (inp[1]) ? node841 : node826;
									assign node826 = (inp[13]) ? node834 : node827;
										assign node827 = (inp[9]) ? 15'b000001111111111 : node828;
											assign node828 = (inp[11]) ? node830 : 15'b000111111111111;
												assign node830 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node834 = (inp[9]) ? node836 : 15'b000001111111111;
											assign node836 = (inp[4]) ? node838 : 15'b000001111111111;
												assign node838 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node841 = (inp[2]) ? node859 : node842;
										assign node842 = (inp[9]) ? node854 : node843;
											assign node843 = (inp[13]) ? node845 : 15'b000001111111111;
												assign node845 = (inp[0]) ? 15'b000000111111111 : node846;
													assign node846 = (inp[4]) ? node848 : 15'b000001111111111;
														assign node848 = (inp[6]) ? 15'b000000111111111 : node849;
															assign node849 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node854 = (inp[0]) ? node856 : 15'b000000111111111;
												assign node856 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node859 = (inp[4]) ? node863 : node860;
											assign node860 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node863 = (inp[6]) ? node865 : 15'b000000011111111;
												assign node865 = (inp[13]) ? node867 : 15'b000000001111111;
													assign node867 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node870 = (inp[11]) ? node918 : node871;
								assign node871 = (inp[4]) ? node893 : node872;
									assign node872 = (inp[2]) ? node886 : node873;
										assign node873 = (inp[7]) ? node881 : node874;
											assign node874 = (inp[1]) ? 15'b000001111111111 : node875;
												assign node875 = (inp[9]) ? node877 : 15'b000111111111111;
													assign node877 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node881 = (inp[1]) ? node883 : 15'b000001111111111;
												assign node883 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node886 = (inp[7]) ? node890 : node887;
											assign node887 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node890 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node893 = (inp[9]) ? node911 : node894;
										assign node894 = (inp[7]) ? node898 : node895;
											assign node895 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node898 = (inp[2]) ? node904 : node899;
												assign node899 = (inp[6]) ? 15'b000000011111111 : node900;
													assign node900 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node904 = (inp[1]) ? node908 : node905;
													assign node905 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node908 = (inp[6]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node911 = (inp[0]) ? node915 : node912;
											assign node912 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node915 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node918 = (inp[13]) ? node938 : node919;
									assign node919 = (inp[4]) ? node931 : node920;
										assign node920 = (inp[6]) ? node928 : node921;
											assign node921 = (inp[9]) ? 15'b000000111111111 : node922;
												assign node922 = (inp[0]) ? 15'b000001111111111 : node923;
													assign node923 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node928 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node931 = (inp[2]) ? node933 : 15'b000000011111111;
											assign node933 = (inp[7]) ? node935 : 15'b000000011111111;
												assign node935 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node938 = (inp[0]) ? node950 : node939;
										assign node939 = (inp[2]) ? node941 : 15'b000000111111111;
											assign node941 = (inp[9]) ? node943 : 15'b000000011111111;
												assign node943 = (inp[7]) ? node947 : node944;
													assign node944 = (inp[6]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node947 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node950 = (inp[7]) ? node956 : node951;
											assign node951 = (inp[2]) ? 15'b000000001111111 : node952;
												assign node952 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node956 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node959 = (inp[1]) ? node1045 : node960;
							assign node960 = (inp[9]) ? node1006 : node961;
								assign node961 = (inp[3]) ? node985 : node962;
									assign node962 = (inp[4]) ? node970 : node963;
										assign node963 = (inp[2]) ? 15'b000001111111111 : node964;
											assign node964 = (inp[6]) ? 15'b000001111111111 : node965;
												assign node965 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node970 = (inp[7]) ? node976 : node971;
											assign node971 = (inp[11]) ? 15'b000000111111111 : node972;
												assign node972 = (inp[0]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node976 = (inp[2]) ? node982 : node977;
												assign node977 = (inp[13]) ? 15'b000000111111111 : node978;
													assign node978 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node982 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node985 = (inp[13]) ? node999 : node986;
										assign node986 = (inp[7]) ? 15'b000000011111111 : node987;
											assign node987 = (inp[2]) ? node993 : node988;
												assign node988 = (inp[0]) ? 15'b000000111111111 : node989;
													assign node989 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node993 = (inp[11]) ? 15'b000001111111111 : node994;
													assign node994 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node999 = (inp[6]) ? 15'b000000011111111 : node1000;
											assign node1000 = (inp[7]) ? node1002 : 15'b000000111111111;
												assign node1002 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1006 = (inp[6]) ? node1028 : node1007;
									assign node1007 = (inp[4]) ? node1013 : node1008;
										assign node1008 = (inp[0]) ? 15'b000000111111111 : node1009;
											assign node1009 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1013 = (inp[0]) ? node1025 : node1014;
											assign node1014 = (inp[3]) ? node1022 : node1015;
												assign node1015 = (inp[11]) ? node1017 : 15'b000000111111111;
													assign node1017 = (inp[13]) ? 15'b000000011111111 : node1018;
														assign node1018 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1022 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node1025 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node1028 = (inp[7]) ? node1034 : node1029;
										assign node1029 = (inp[13]) ? 15'b000000001111111 : node1030;
											assign node1030 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node1034 = (inp[11]) ? node1042 : node1035;
											assign node1035 = (inp[0]) ? node1037 : 15'b000000011111111;
												assign node1037 = (inp[4]) ? 15'b000000001111111 : node1038;
													assign node1038 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node1042 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
							assign node1045 = (inp[0]) ? node1091 : node1046;
								assign node1046 = (inp[2]) ? node1068 : node1047;
									assign node1047 = (inp[13]) ? node1061 : node1048;
										assign node1048 = (inp[7]) ? node1056 : node1049;
											assign node1049 = (inp[11]) ? node1053 : node1050;
												assign node1050 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node1053 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1056 = (inp[6]) ? node1058 : 15'b000000111111111;
												assign node1058 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node1061 = (inp[3]) ? node1065 : node1062;
											assign node1062 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1065 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1068 = (inp[6]) ? node1076 : node1069;
										assign node1069 = (inp[13]) ? 15'b000000011111111 : node1070;
											assign node1070 = (inp[3]) ? node1072 : 15'b000000111111111;
												assign node1072 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1076 = (inp[4]) ? node1082 : node1077;
											assign node1077 = (inp[9]) ? 15'b000000000111111 : node1078;
												assign node1078 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1082 = (inp[7]) ? node1088 : node1083;
												assign node1083 = (inp[3]) ? 15'b000000001111111 : node1084;
													assign node1084 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1088 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1091 = (inp[7]) ? node1107 : node1092;
									assign node1092 = (inp[11]) ? node1098 : node1093;
										assign node1093 = (inp[13]) ? node1095 : 15'b000000011111111;
											assign node1095 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1098 = (inp[6]) ? node1104 : node1099;
											assign node1099 = (inp[13]) ? node1101 : 15'b000000011111111;
												assign node1101 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node1104 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1107 = (inp[13]) ? node1123 : node1108;
										assign node1108 = (inp[9]) ? node1116 : node1109;
											assign node1109 = (inp[11]) ? node1111 : 15'b000000011111111;
												assign node1111 = (inp[6]) ? 15'b000000001111111 : node1112;
													assign node1112 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1116 = (inp[3]) ? node1120 : node1117;
												assign node1117 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1120 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1123 = (inp[3]) ? node1129 : node1124;
											assign node1124 = (inp[2]) ? node1126 : 15'b000000001111111;
												assign node1126 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1129 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node1132 = (inp[14]) ? node1318 : node1133;
						assign node1133 = (inp[2]) ? node1229 : node1134;
							assign node1134 = (inp[9]) ? node1184 : node1135;
								assign node1135 = (inp[1]) ? node1161 : node1136;
									assign node1136 = (inp[6]) ? node1154 : node1137;
										assign node1137 = (inp[4]) ? node1147 : node1138;
											assign node1138 = (inp[0]) ? node1144 : node1139;
												assign node1139 = (inp[3]) ? node1141 : 15'b000011111111111;
													assign node1141 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1144 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1147 = (inp[3]) ? node1149 : 15'b000001111111111;
												assign node1149 = (inp[0]) ? 15'b000000111111111 : node1150;
													assign node1150 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1154 = (inp[11]) ? 15'b000000011111111 : node1155;
											assign node1155 = (inp[13]) ? node1157 : 15'b000001111111111;
												assign node1157 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node1161 = (inp[13]) ? node1171 : node1162;
										assign node1162 = (inp[6]) ? 15'b000000011111111 : node1163;
											assign node1163 = (inp[3]) ? node1165 : 15'b000001111111111;
												assign node1165 = (inp[7]) ? 15'b000000111111111 : node1166;
													assign node1166 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1171 = (inp[4]) ? node1181 : node1172;
											assign node1172 = (inp[3]) ? node1174 : 15'b000000111111111;
												assign node1174 = (inp[11]) ? node1176 : 15'b000000011111111;
													assign node1176 = (inp[0]) ? 15'b000000011111111 : node1177;
														assign node1177 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1181 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1184 = (inp[11]) ? node1204 : node1185;
									assign node1185 = (inp[13]) ? node1197 : node1186;
										assign node1186 = (inp[0]) ? node1192 : node1187;
											assign node1187 = (inp[7]) ? 15'b000000111111111 : node1188;
												assign node1188 = (inp[6]) ? 15'b000001111111111 : 15'b000111111111111;
											assign node1192 = (inp[6]) ? node1194 : 15'b000000111111111;
												assign node1194 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1197 = (inp[3]) ? node1201 : node1198;
											assign node1198 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1201 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1204 = (inp[1]) ? node1216 : node1205;
										assign node1205 = (inp[13]) ? node1209 : node1206;
											assign node1206 = (inp[0]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node1209 = (inp[0]) ? node1211 : 15'b000000111111111;
												assign node1211 = (inp[4]) ? 15'b000000001111111 : node1212;
													assign node1212 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1216 = (inp[7]) ? 15'b000000000111111 : node1217;
											assign node1217 = (inp[13]) ? node1223 : node1218;
												assign node1218 = (inp[6]) ? 15'b000000011111111 : node1219;
													assign node1219 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1223 = (inp[4]) ? node1225 : 15'b000000001111111;
													assign node1225 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1229 = (inp[9]) ? node1283 : node1230;
								assign node1230 = (inp[13]) ? node1248 : node1231;
									assign node1231 = (inp[11]) ? node1243 : node1232;
										assign node1232 = (inp[3]) ? node1234 : 15'b000000011111111;
											assign node1234 = (inp[1]) ? node1236 : 15'b000000111111111;
												assign node1236 = (inp[0]) ? 15'b000000011111111 : node1237;
													assign node1237 = (inp[7]) ? node1239 : 15'b000000111111111;
														assign node1239 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1243 = (inp[3]) ? 15'b000000011111111 : node1244;
											assign node1244 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node1248 = (inp[1]) ? node1262 : node1249;
										assign node1249 = (inp[0]) ? node1253 : node1250;
											assign node1250 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1253 = (inp[3]) ? node1255 : 15'b000000111111111;
												assign node1255 = (inp[4]) ? 15'b000000001111111 : node1256;
													assign node1256 = (inp[11]) ? node1258 : 15'b000000011111111;
														assign node1258 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1262 = (inp[7]) ? node1272 : node1263;
											assign node1263 = (inp[0]) ? node1267 : node1264;
												assign node1264 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1267 = (inp[4]) ? node1269 : 15'b000000001111111;
													assign node1269 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1272 = (inp[4]) ? node1280 : node1273;
												assign node1273 = (inp[11]) ? node1275 : 15'b000000001111111;
													assign node1275 = (inp[3]) ? 15'b000000000111111 : node1276;
														assign node1276 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1280 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1283 = (inp[4]) ? node1301 : node1284;
									assign node1284 = (inp[0]) ? node1290 : node1285;
										assign node1285 = (inp[3]) ? 15'b000000011111111 : node1286;
											assign node1286 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1290 = (inp[1]) ? node1296 : node1291;
											assign node1291 = (inp[7]) ? 15'b000000011111111 : node1292;
												assign node1292 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1296 = (inp[7]) ? node1298 : 15'b000000001111111;
												assign node1298 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node1301 = (inp[6]) ? node1307 : node1302;
										assign node1302 = (inp[11]) ? node1304 : 15'b000000001111111;
											assign node1304 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node1307 = (inp[11]) ? node1313 : node1308;
											assign node1308 = (inp[7]) ? 15'b000000000111111 : node1309;
												assign node1309 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1313 = (inp[3]) ? 15'b000000000011111 : node1314;
												assign node1314 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node1318 = (inp[4]) ? node1394 : node1319;
							assign node1319 = (inp[1]) ? node1363 : node1320;
								assign node1320 = (inp[6]) ? node1346 : node1321;
									assign node1321 = (inp[2]) ? node1339 : node1322;
										assign node1322 = (inp[9]) ? node1328 : node1323;
											assign node1323 = (inp[11]) ? 15'b000000111111111 : node1324;
												assign node1324 = (inp[0]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node1328 = (inp[11]) ? node1334 : node1329;
												assign node1329 = (inp[13]) ? 15'b000000011111111 : node1330;
													assign node1330 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1334 = (inp[0]) ? 15'b000000011111111 : node1335;
													assign node1335 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1339 = (inp[0]) ? 15'b000000011111111 : node1340;
											assign node1340 = (inp[11]) ? 15'b000000011111111 : node1341;
												assign node1341 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1346 = (inp[7]) ? node1358 : node1347;
										assign node1347 = (inp[2]) ? node1355 : node1348;
											assign node1348 = (inp[3]) ? 15'b000000011111111 : node1349;
												assign node1349 = (inp[11]) ? node1351 : 15'b000000111111111;
													assign node1351 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1355 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1358 = (inp[3]) ? node1360 : 15'b000000001111111;
											assign node1360 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1363 = (inp[9]) ? node1379 : node1364;
									assign node1364 = (inp[7]) ? node1368 : node1365;
										assign node1365 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node1368 = (inp[0]) ? node1374 : node1369;
											assign node1369 = (inp[13]) ? 15'b000000001111111 : node1370;
												assign node1370 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1374 = (inp[6]) ? 15'b000000000011111 : node1375;
												assign node1375 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1379 = (inp[11]) ? node1389 : node1380;
										assign node1380 = (inp[0]) ? node1384 : node1381;
											assign node1381 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node1384 = (inp[2]) ? 15'b000000000111111 : node1385;
												assign node1385 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node1389 = (inp[0]) ? 15'b000000000011111 : node1390;
											assign node1390 = (inp[13]) ? 15'b000000000111111 : 15'b000000000011111;
							assign node1394 = (inp[3]) ? node1440 : node1395;
								assign node1395 = (inp[2]) ? node1419 : node1396;
									assign node1396 = (inp[7]) ? node1402 : node1397;
										assign node1397 = (inp[13]) ? 15'b000000001111111 : node1398;
											assign node1398 = (inp[9]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node1402 = (inp[9]) ? node1414 : node1403;
											assign node1403 = (inp[11]) ? node1409 : node1404;
												assign node1404 = (inp[1]) ? node1406 : 15'b000000011111111;
													assign node1406 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1409 = (inp[1]) ? node1411 : 15'b000000001111111;
													assign node1411 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1414 = (inp[11]) ? node1416 : 15'b000000000111111;
												assign node1416 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1419 = (inp[1]) ? node1431 : node1420;
										assign node1420 = (inp[13]) ? 15'b000000000111111 : node1421;
											assign node1421 = (inp[6]) ? 15'b000000000111111 : node1422;
												assign node1422 = (inp[11]) ? 15'b000000001111111 : node1423;
													assign node1423 = (inp[9]) ? node1425 : 15'b000000011111111;
														assign node1425 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1431 = (inp[11]) ? node1433 : 15'b000000000111111;
											assign node1433 = (inp[6]) ? node1437 : node1434;
												assign node1434 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node1437 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1440 = (inp[7]) ? node1456 : node1441;
									assign node1441 = (inp[13]) ? node1449 : node1442;
										assign node1442 = (inp[11]) ? node1446 : node1443;
											assign node1443 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1446 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1449 = (inp[9]) ? node1451 : 15'b000000000111111;
											assign node1451 = (inp[0]) ? node1453 : 15'b000000000111111;
												assign node1453 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1456 = (inp[2]) ? node1466 : node1457;
										assign node1457 = (inp[0]) ? node1461 : node1458;
											assign node1458 = (inp[13]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node1461 = (inp[1]) ? 15'b000000000011111 : node1462;
												assign node1462 = (inp[11]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node1466 = (inp[6]) ? node1468 : 15'b000000001111111;
											assign node1468 = (inp[13]) ? 15'b000000000001111 : node1469;
												assign node1469 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
			assign node1473 = (inp[1]) ? node2185 : node1474;
				assign node1474 = (inp[7]) ? node1806 : node1475;
					assign node1475 = (inp[4]) ? node1637 : node1476;
						assign node1476 = (inp[13]) ? node1552 : node1477;
							assign node1477 = (inp[9]) ? node1509 : node1478;
								assign node1478 = (inp[2]) ? node1494 : node1479;
									assign node1479 = (inp[14]) ? node1491 : node1480;
										assign node1480 = (inp[11]) ? node1486 : node1481;
											assign node1481 = (inp[8]) ? node1483 : 15'b000111111111111;
												assign node1483 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1486 = (inp[5]) ? 15'b000001111111111 : node1487;
												assign node1487 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node1491 = (inp[6]) ? 15'b000011111111111 : 15'b000001111111111;
									assign node1494 = (inp[8]) ? node1500 : node1495;
										assign node1495 = (inp[0]) ? 15'b000001111111111 : node1496;
											assign node1496 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node1500 = (inp[3]) ? 15'b000000111111111 : node1501;
											assign node1501 = (inp[0]) ? 15'b000000111111111 : node1502;
												assign node1502 = (inp[6]) ? node1504 : 15'b000001111111111;
													assign node1504 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node1509 = (inp[2]) ? node1539 : node1510;
									assign node1510 = (inp[11]) ? node1522 : node1511;
										assign node1511 = (inp[8]) ? 15'b000001111111111 : node1512;
											assign node1512 = (inp[3]) ? node1516 : node1513;
												assign node1513 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1516 = (inp[5]) ? node1518 : 15'b000011111111111;
													assign node1518 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1522 = (inp[14]) ? node1530 : node1523;
											assign node1523 = (inp[6]) ? node1525 : 15'b000001111111111;
												assign node1525 = (inp[3]) ? 15'b000000011111111 : node1526;
													assign node1526 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1530 = (inp[3]) ? node1532 : 15'b000000011111111;
												assign node1532 = (inp[5]) ? 15'b000000111111111 : node1533;
													assign node1533 = (inp[0]) ? 15'b000000111111111 : node1534;
														assign node1534 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1539 = (inp[6]) ? node1545 : node1540;
										assign node1540 = (inp[5]) ? 15'b000000111111111 : node1541;
											assign node1541 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node1545 = (inp[8]) ? 15'b000000001111111 : node1546;
											assign node1546 = (inp[11]) ? 15'b000000011111111 : node1547;
												assign node1547 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node1552 = (inp[14]) ? node1600 : node1553;
								assign node1553 = (inp[3]) ? node1579 : node1554;
									assign node1554 = (inp[0]) ? node1574 : node1555;
										assign node1555 = (inp[5]) ? node1565 : node1556;
											assign node1556 = (inp[2]) ? 15'b000001111111111 : node1557;
												assign node1557 = (inp[8]) ? 15'b000011111111111 : node1558;
													assign node1558 = (inp[11]) ? node1560 : 15'b000111111111111;
														assign node1560 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1565 = (inp[8]) ? 15'b000000111111111 : node1566;
												assign node1566 = (inp[11]) ? node1568 : 15'b000011111111111;
													assign node1568 = (inp[2]) ? node1570 : 15'b000001111111111;
														assign node1570 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1574 = (inp[5]) ? 15'b000000111111111 : node1575;
											assign node1575 = (inp[11]) ? 15'b000000011111111 : 15'b000001111111111;
									assign node1579 = (inp[6]) ? node1589 : node1580;
										assign node1580 = (inp[11]) ? node1586 : node1581;
											assign node1581 = (inp[5]) ? 15'b000000111111111 : node1582;
												assign node1582 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1586 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node1589 = (inp[9]) ? node1595 : node1590;
											assign node1590 = (inp[8]) ? node1592 : 15'b000000111111111;
												assign node1592 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1595 = (inp[2]) ? 15'b000000001111111 : node1596;
												assign node1596 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node1600 = (inp[9]) ? node1616 : node1601;
									assign node1601 = (inp[11]) ? node1607 : node1602;
										assign node1602 = (inp[3]) ? node1604 : 15'b000000111111111;
											assign node1604 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1607 = (inp[0]) ? node1613 : node1608;
											assign node1608 = (inp[3]) ? 15'b000000011111111 : node1609;
												assign node1609 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1613 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node1616 = (inp[8]) ? node1622 : node1617;
										assign node1617 = (inp[0]) ? node1619 : 15'b000000111111111;
											assign node1619 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1622 = (inp[11]) ? node1630 : node1623;
											assign node1623 = (inp[6]) ? node1625 : 15'b000001111111111;
												assign node1625 = (inp[2]) ? 15'b000000001111111 : node1626;
													assign node1626 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1630 = (inp[0]) ? 15'b000000000111111 : node1631;
												assign node1631 = (inp[3]) ? node1633 : 15'b000000001111111;
													assign node1633 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node1637 = (inp[8]) ? node1739 : node1638;
							assign node1638 = (inp[2]) ? node1696 : node1639;
								assign node1639 = (inp[11]) ? node1675 : node1640;
									assign node1640 = (inp[6]) ? node1658 : node1641;
										assign node1641 = (inp[0]) ? node1643 : 15'b000011111111111;
											assign node1643 = (inp[13]) ? node1649 : node1644;
												assign node1644 = (inp[9]) ? node1646 : 15'b000001111111111;
													assign node1646 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1649 = (inp[5]) ? 15'b000000111111111 : node1650;
													assign node1650 = (inp[3]) ? 15'b000000111111111 : node1651;
														assign node1651 = (inp[9]) ? 15'b000001111111111 : node1652;
															assign node1652 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node1658 = (inp[3]) ? node1664 : node1659;
											assign node1659 = (inp[13]) ? 15'b000000011111111 : node1660;
												assign node1660 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1664 = (inp[5]) ? node1670 : node1665;
												assign node1665 = (inp[9]) ? 15'b000000111111111 : node1666;
													assign node1666 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1670 = (inp[14]) ? node1672 : 15'b000000011111111;
													assign node1672 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1675 = (inp[9]) ? node1685 : node1676;
										assign node1676 = (inp[5]) ? node1682 : node1677;
											assign node1677 = (inp[6]) ? node1679 : 15'b000001111111111;
												assign node1679 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1682 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1685 = (inp[0]) ? node1689 : node1686;
											assign node1686 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1689 = (inp[3]) ? 15'b000000000111111 : node1690;
												assign node1690 = (inp[6]) ? node1692 : 15'b000000011111111;
													assign node1692 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1696 = (inp[14]) ? node1716 : node1697;
									assign node1697 = (inp[3]) ? node1703 : node1698;
										assign node1698 = (inp[6]) ? node1700 : 15'b000000111111111;
											assign node1700 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1703 = (inp[13]) ? node1707 : node1704;
											assign node1704 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1707 = (inp[11]) ? node1711 : node1708;
												assign node1708 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1711 = (inp[5]) ? 15'b000000001111111 : node1712;
													assign node1712 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1716 = (inp[9]) ? node1726 : node1717;
										assign node1717 = (inp[5]) ? 15'b000000000111111 : node1718;
											assign node1718 = (inp[3]) ? node1720 : 15'b000000011111111;
												assign node1720 = (inp[13]) ? 15'b000000111111111 : node1721;
													assign node1721 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1726 = (inp[11]) ? node1732 : node1727;
											assign node1727 = (inp[0]) ? 15'b000000001111111 : node1728;
												assign node1728 = (inp[5]) ? 15'b000000000111111 : 15'b000000111111111;
											assign node1732 = (inp[0]) ? node1734 : 15'b000000001111111;
												assign node1734 = (inp[3]) ? 15'b000000000111111 : node1735;
													assign node1735 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1739 = (inp[9]) ? node1767 : node1740;
								assign node1740 = (inp[13]) ? node1752 : node1741;
									assign node1741 = (inp[6]) ? node1747 : node1742;
										assign node1742 = (inp[2]) ? node1744 : 15'b000001111111111;
											assign node1744 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1747 = (inp[0]) ? node1749 : 15'b000000111111111;
											assign node1749 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1752 = (inp[0]) ? node1762 : node1753;
										assign node1753 = (inp[11]) ? node1757 : node1754;
											assign node1754 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1757 = (inp[14]) ? 15'b000000001111111 : node1758;
												assign node1758 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1762 = (inp[14]) ? 15'b000000000111111 : node1763;
											assign node1763 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1767 = (inp[6]) ? node1791 : node1768;
									assign node1768 = (inp[3]) ? node1780 : node1769;
										assign node1769 = (inp[5]) ? node1773 : node1770;
											assign node1770 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1773 = (inp[11]) ? node1775 : 15'b000000001111111;
												assign node1775 = (inp[0]) ? 15'b000000001111111 : node1776;
													assign node1776 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1780 = (inp[2]) ? node1788 : node1781;
											assign node1781 = (inp[11]) ? node1783 : 15'b000000001111111;
												assign node1783 = (inp[0]) ? node1785 : 15'b000000001111111;
													assign node1785 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1788 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1791 = (inp[3]) ? node1801 : node1792;
										assign node1792 = (inp[5]) ? node1796 : node1793;
											assign node1793 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1796 = (inp[14]) ? 15'b000000000111111 : node1797;
												assign node1797 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1801 = (inp[0]) ? node1803 : 15'b000000000111111;
											assign node1803 = (inp[2]) ? 15'b000000000011111 : 15'b000000000001111;
					assign node1806 = (inp[0]) ? node2008 : node1807;
						assign node1807 = (inp[11]) ? node1909 : node1808;
							assign node1808 = (inp[5]) ? node1858 : node1809;
								assign node1809 = (inp[14]) ? node1831 : node1810;
									assign node1810 = (inp[9]) ? node1824 : node1811;
										assign node1811 = (inp[8]) ? node1817 : node1812;
											assign node1812 = (inp[4]) ? 15'b000011111111111 : node1813;
												assign node1813 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1817 = (inp[3]) ? node1821 : node1818;
												assign node1818 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1821 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1824 = (inp[2]) ? 15'b000000001111111 : node1825;
											assign node1825 = (inp[8]) ? 15'b000000111111111 : node1826;
												assign node1826 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1831 = (inp[6]) ? node1847 : node1832;
										assign node1832 = (inp[2]) ? node1836 : node1833;
											assign node1833 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1836 = (inp[13]) ? node1842 : node1837;
												assign node1837 = (inp[8]) ? 15'b000000111111111 : node1838;
													assign node1838 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1842 = (inp[9]) ? 15'b000000011111111 : node1843;
													assign node1843 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1847 = (inp[4]) ? node1853 : node1848;
											assign node1848 = (inp[8]) ? node1850 : 15'b000000111111111;
												assign node1850 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1853 = (inp[2]) ? 15'b000000011111111 : node1854;
												assign node1854 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1858 = (inp[6]) ? node1886 : node1859;
									assign node1859 = (inp[3]) ? node1873 : node1860;
										assign node1860 = (inp[9]) ? node1870 : node1861;
											assign node1861 = (inp[4]) ? node1867 : node1862;
												assign node1862 = (inp[2]) ? 15'b000001111111111 : node1863;
													assign node1863 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1867 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1870 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1873 = (inp[13]) ? node1881 : node1874;
											assign node1874 = (inp[4]) ? 15'b000000011111111 : node1875;
												assign node1875 = (inp[9]) ? node1877 : 15'b000001111111111;
													assign node1877 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1881 = (inp[2]) ? node1883 : 15'b000000011111111;
												assign node1883 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1886 = (inp[13]) ? node1902 : node1887;
										assign node1887 = (inp[8]) ? node1897 : node1888;
											assign node1888 = (inp[14]) ? node1892 : node1889;
												assign node1889 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1892 = (inp[4]) ? 15'b000000011111111 : node1893;
													assign node1893 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1897 = (inp[4]) ? 15'b000000011111111 : node1898;
												assign node1898 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1902 = (inp[4]) ? node1904 : 15'b000000111111111;
											assign node1904 = (inp[3]) ? node1906 : 15'b000000001111111;
												assign node1906 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
							assign node1909 = (inp[9]) ? node1971 : node1910;
								assign node1910 = (inp[3]) ? node1938 : node1911;
									assign node1911 = (inp[4]) ? node1923 : node1912;
										assign node1912 = (inp[13]) ? node1920 : node1913;
											assign node1913 = (inp[14]) ? 15'b000011111111111 : node1914;
												assign node1914 = (inp[8]) ? 15'b000001111111111 : node1915;
													assign node1915 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1920 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1923 = (inp[5]) ? node1931 : node1924;
											assign node1924 = (inp[14]) ? node1926 : 15'b000001111111111;
												assign node1926 = (inp[6]) ? 15'b000000011111111 : node1927;
													assign node1927 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1931 = (inp[14]) ? 15'b000000001111111 : node1932;
												assign node1932 = (inp[6]) ? node1934 : 15'b000000111111111;
													assign node1934 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1938 = (inp[13]) ? node1958 : node1939;
										assign node1939 = (inp[2]) ? node1949 : node1940;
											assign node1940 = (inp[6]) ? node1942 : 15'b000000111111111;
												assign node1942 = (inp[5]) ? node1944 : 15'b000000001111111;
													assign node1944 = (inp[14]) ? 15'b000000011111111 : node1945;
														assign node1945 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1949 = (inp[5]) ? node1953 : node1950;
												assign node1950 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1953 = (inp[14]) ? 15'b000000001111111 : node1954;
													assign node1954 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1958 = (inp[8]) ? node1960 : 15'b000000011111111;
											assign node1960 = (inp[6]) ? node1966 : node1961;
												assign node1961 = (inp[2]) ? 15'b000000000111111 : node1962;
													assign node1962 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1966 = (inp[5]) ? 15'b000000000111111 : node1967;
													assign node1967 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1971 = (inp[14]) ? node1991 : node1972;
									assign node1972 = (inp[4]) ? node1982 : node1973;
										assign node1973 = (inp[2]) ? node1979 : node1974;
											assign node1974 = (inp[13]) ? 15'b000000011111111 : node1975;
												assign node1975 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node1979 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node1982 = (inp[5]) ? node1988 : node1983;
											assign node1983 = (inp[6]) ? 15'b000000001111111 : node1984;
												assign node1984 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1988 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node1991 = (inp[5]) ? node2001 : node1992;
										assign node1992 = (inp[6]) ? 15'b000000000111111 : node1993;
											assign node1993 = (inp[13]) ? node1997 : node1994;
												assign node1994 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1997 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2001 = (inp[3]) ? node2005 : node2002;
											assign node2002 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2005 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node2008 = (inp[14]) ? node2086 : node2009;
							assign node2009 = (inp[6]) ? node2039 : node2010;
								assign node2010 = (inp[8]) ? node2024 : node2011;
									assign node2011 = (inp[3]) ? node2019 : node2012;
										assign node2012 = (inp[13]) ? node2016 : node2013;
											assign node2013 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2016 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node2019 = (inp[13]) ? 15'b000000001111111 : node2020;
											assign node2020 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2024 = (inp[9]) ? 15'b000000001111111 : node2025;
										assign node2025 = (inp[11]) ? node2029 : node2026;
											assign node2026 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2029 = (inp[13]) ? node2033 : node2030;
												assign node2030 = (inp[4]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node2033 = (inp[3]) ? 15'b000000001111111 : node2034;
													assign node2034 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2039 = (inp[5]) ? node2061 : node2040;
									assign node2040 = (inp[9]) ? node2050 : node2041;
										assign node2041 = (inp[11]) ? node2045 : node2042;
											assign node2042 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2045 = (inp[4]) ? 15'b000000001111111 : node2046;
												assign node2046 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2050 = (inp[4]) ? node2058 : node2051;
											assign node2051 = (inp[11]) ? 15'b000000011111111 : node2052;
												assign node2052 = (inp[8]) ? 15'b000000011111111 : node2053;
													assign node2053 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2058 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2061 = (inp[13]) ? node2071 : node2062;
										assign node2062 = (inp[9]) ? 15'b000000000111111 : node2063;
											assign node2063 = (inp[2]) ? node2065 : 15'b000000011111111;
												assign node2065 = (inp[8]) ? 15'b000000001111111 : node2066;
													assign node2066 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2071 = (inp[3]) ? node2077 : node2072;
											assign node2072 = (inp[8]) ? node2074 : 15'b000000001111111;
												assign node2074 = (inp[2]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node2077 = (inp[2]) ? node2079 : 15'b000000001111111;
												assign node2079 = (inp[4]) ? node2081 : 15'b000000000011111;
													assign node2081 = (inp[8]) ? node2083 : 15'b000000000001111;
														assign node2083 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node2086 = (inp[6]) ? node2136 : node2087;
								assign node2087 = (inp[9]) ? node2105 : node2088;
									assign node2088 = (inp[8]) ? node2094 : node2089;
										assign node2089 = (inp[11]) ? node2091 : 15'b000000011111111;
											assign node2091 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2094 = (inp[5]) ? node2098 : node2095;
											assign node2095 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2098 = (inp[2]) ? node2100 : 15'b000000001111111;
												assign node2100 = (inp[3]) ? node2102 : 15'b000000001111111;
													assign node2102 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2105 = (inp[3]) ? node2123 : node2106;
										assign node2106 = (inp[2]) ? node2118 : node2107;
											assign node2107 = (inp[4]) ? node2113 : node2108;
												assign node2108 = (inp[8]) ? 15'b000000011111111 : node2109;
													assign node2109 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2113 = (inp[13]) ? 15'b000000000011111 : node2114;
													assign node2114 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2118 = (inp[13]) ? 15'b000000000111111 : node2119;
												assign node2119 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2123 = (inp[4]) ? node2127 : node2124;
											assign node2124 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2127 = (inp[5]) ? 15'b000000000011111 : node2128;
												assign node2128 = (inp[13]) ? node2130 : 15'b000000000111111;
													assign node2130 = (inp[2]) ? 15'b000000000011111 : node2131;
														assign node2131 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2136 = (inp[13]) ? node2156 : node2137;
									assign node2137 = (inp[11]) ? node2147 : node2138;
										assign node2138 = (inp[5]) ? node2142 : node2139;
											assign node2139 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2142 = (inp[9]) ? node2144 : 15'b000000000111111;
												assign node2144 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2147 = (inp[4]) ? node2153 : node2148;
											assign node2148 = (inp[8]) ? 15'b000000000111111 : node2149;
												assign node2149 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2153 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2156 = (inp[8]) ? node2172 : node2157;
										assign node2157 = (inp[9]) ? 15'b000000000001111 : node2158;
											assign node2158 = (inp[5]) ? node2164 : node2159;
												assign node2159 = (inp[11]) ? 15'b000000001111111 : node2160;
													assign node2160 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2164 = (inp[4]) ? node2168 : node2165;
													assign node2165 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2168 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2172 = (inp[4]) ? node2182 : node2173;
											assign node2173 = (inp[3]) ? node2179 : node2174;
												assign node2174 = (inp[2]) ? node2176 : 15'b000000000111111;
													assign node2176 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node2179 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node2182 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node2185 = (inp[13]) ? node2551 : node2186;
					assign node2186 = (inp[11]) ? node2360 : node2187;
						assign node2187 = (inp[5]) ? node2273 : node2188;
							assign node2188 = (inp[0]) ? node2236 : node2189;
								assign node2189 = (inp[3]) ? node2213 : node2190;
									assign node2190 = (inp[6]) ? node2206 : node2191;
										assign node2191 = (inp[7]) ? node2199 : node2192;
											assign node2192 = (inp[14]) ? node2196 : node2193;
												assign node2193 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2196 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2199 = (inp[8]) ? node2201 : 15'b000001111111111;
												assign node2201 = (inp[14]) ? 15'b000000111111111 : node2202;
													assign node2202 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2206 = (inp[4]) ? node2210 : node2207;
											assign node2207 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2210 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node2213 = (inp[4]) ? node2225 : node2214;
										assign node2214 = (inp[9]) ? node2220 : node2215;
											assign node2215 = (inp[8]) ? node2217 : 15'b000001111111111;
												assign node2217 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2220 = (inp[7]) ? 15'b000000011111111 : node2221;
												assign node2221 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node2225 = (inp[9]) ? node2233 : node2226;
											assign node2226 = (inp[7]) ? node2228 : 15'b000000111111111;
												assign node2228 = (inp[2]) ? 15'b000000011111111 : node2229;
													assign node2229 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2233 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2236 = (inp[7]) ? node2252 : node2237;
									assign node2237 = (inp[14]) ? node2247 : node2238;
										assign node2238 = (inp[6]) ? node2242 : node2239;
											assign node2239 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2242 = (inp[9]) ? 15'b000000011111111 : node2243;
												assign node2243 = (inp[2]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node2247 = (inp[2]) ? node2249 : 15'b000000111111111;
											assign node2249 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2252 = (inp[4]) ? node2258 : node2253;
										assign node2253 = (inp[6]) ? 15'b000000001111111 : node2254;
											assign node2254 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2258 = (inp[2]) ? node2268 : node2259;
											assign node2259 = (inp[14]) ? node2265 : node2260;
												assign node2260 = (inp[8]) ? 15'b000000011111111 : node2261;
													assign node2261 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2265 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2268 = (inp[3]) ? node2270 : 15'b000000000111111;
												assign node2270 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2273 = (inp[14]) ? node2317 : node2274;
								assign node2274 = (inp[6]) ? node2290 : node2275;
									assign node2275 = (inp[7]) ? node2283 : node2276;
										assign node2276 = (inp[2]) ? node2278 : 15'b000000111111111;
											assign node2278 = (inp[4]) ? 15'b000000011111111 : node2279;
												assign node2279 = (inp[0]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node2283 = (inp[0]) ? 15'b000000001111111 : node2284;
											assign node2284 = (inp[4]) ? 15'b000000011111111 : node2285;
												assign node2285 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2290 = (inp[2]) ? node2306 : node2291;
										assign node2291 = (inp[9]) ? node2299 : node2292;
											assign node2292 = (inp[8]) ? node2294 : 15'b000000111111111;
												assign node2294 = (inp[3]) ? 15'b000000011111111 : node2295;
													assign node2295 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2299 = (inp[8]) ? 15'b000000001111111 : node2300;
												assign node2300 = (inp[4]) ? node2302 : 15'b000000111111111;
													assign node2302 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2306 = (inp[4]) ? node2310 : node2307;
											assign node2307 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2310 = (inp[7]) ? node2314 : node2311;
												assign node2311 = (inp[0]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node2314 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2317 = (inp[4]) ? node2341 : node2318;
									assign node2318 = (inp[6]) ? node2330 : node2319;
										assign node2319 = (inp[2]) ? node2325 : node2320;
											assign node2320 = (inp[8]) ? node2322 : 15'b000000011111111;
												assign node2322 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2325 = (inp[7]) ? 15'b000000001111111 : node2326;
												assign node2326 = (inp[8]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node2330 = (inp[9]) ? node2336 : node2331;
											assign node2331 = (inp[7]) ? node2333 : 15'b000000011111111;
												assign node2333 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2336 = (inp[3]) ? 15'b000000000011111 : node2337;
												assign node2337 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2341 = (inp[0]) ? node2347 : node2342;
										assign node2342 = (inp[7]) ? node2344 : 15'b000000111111111;
											assign node2344 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2347 = (inp[2]) ? node2353 : node2348;
											assign node2348 = (inp[3]) ? node2350 : 15'b000000000111111;
												assign node2350 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2353 = (inp[3]) ? node2355 : 15'b000000000111111;
												assign node2355 = (inp[8]) ? 15'b000000000011111 : node2356;
													assign node2356 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node2360 = (inp[8]) ? node2458 : node2361;
							assign node2361 = (inp[3]) ? node2405 : node2362;
								assign node2362 = (inp[6]) ? node2386 : node2363;
									assign node2363 = (inp[4]) ? node2379 : node2364;
										assign node2364 = (inp[9]) ? node2376 : node2365;
											assign node2365 = (inp[5]) ? node2371 : node2366;
												assign node2366 = (inp[0]) ? 15'b000001111111111 : node2367;
													assign node2367 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2371 = (inp[0]) ? 15'b000000111111111 : node2372;
													assign node2372 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2376 = (inp[5]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node2379 = (inp[9]) ? node2383 : node2380;
											assign node2380 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2383 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2386 = (inp[2]) ? node2396 : node2387;
										assign node2387 = (inp[4]) ? node2393 : node2388;
											assign node2388 = (inp[0]) ? node2390 : 15'b000000111111111;
												assign node2390 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2393 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2396 = (inp[4]) ? 15'b000000000111111 : node2397;
											assign node2397 = (inp[0]) ? 15'b000000001111111 : node2398;
												assign node2398 = (inp[5]) ? node2400 : 15'b000000011111111;
													assign node2400 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2405 = (inp[5]) ? node2435 : node2406;
									assign node2406 = (inp[0]) ? node2416 : node2407;
										assign node2407 = (inp[14]) ? node2411 : node2408;
											assign node2408 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2411 = (inp[2]) ? node2413 : 15'b000000011111111;
												assign node2413 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2416 = (inp[6]) ? node2428 : node2417;
											assign node2417 = (inp[9]) ? node2423 : node2418;
												assign node2418 = (inp[4]) ? node2420 : 15'b000000011111111;
													assign node2420 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2423 = (inp[4]) ? node2425 : 15'b000000001111111;
													assign node2425 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2428 = (inp[7]) ? 15'b000000000111111 : node2429;
												assign node2429 = (inp[2]) ? node2431 : 15'b000000001111111;
													assign node2431 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2435 = (inp[6]) ? node2445 : node2436;
										assign node2436 = (inp[9]) ? node2438 : 15'b000000111111111;
											assign node2438 = (inp[4]) ? 15'b000000000111111 : node2439;
												assign node2439 = (inp[0]) ? node2441 : 15'b000000001111111;
													assign node2441 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2445 = (inp[14]) ? node2449 : node2446;
											assign node2446 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2449 = (inp[9]) ? 15'b000000000011111 : node2450;
												assign node2450 = (inp[7]) ? node2452 : 15'b000000000111111;
													assign node2452 = (inp[4]) ? node2454 : 15'b000000000111111;
														assign node2454 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node2458 = (inp[5]) ? node2512 : node2459;
								assign node2459 = (inp[3]) ? node2483 : node2460;
									assign node2460 = (inp[2]) ? node2466 : node2461;
										assign node2461 = (inp[0]) ? 15'b000000001111111 : node2462;
											assign node2462 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2466 = (inp[0]) ? node2474 : node2467;
											assign node2467 = (inp[6]) ? node2471 : node2468;
												assign node2468 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2471 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2474 = (inp[4]) ? node2478 : node2475;
												assign node2475 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2478 = (inp[6]) ? 15'b000000000111111 : node2479;
													assign node2479 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2483 = (inp[4]) ? node2497 : node2484;
										assign node2484 = (inp[0]) ? node2490 : node2485;
											assign node2485 = (inp[7]) ? 15'b000000001111111 : node2486;
												assign node2486 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2490 = (inp[14]) ? node2494 : node2491;
												assign node2491 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2494 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2497 = (inp[9]) ? node2505 : node2498;
											assign node2498 = (inp[7]) ? node2500 : 15'b000000001111111;
												assign node2500 = (inp[6]) ? node2502 : 15'b000000001111111;
													assign node2502 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2505 = (inp[0]) ? 15'b000000000011111 : node2506;
												assign node2506 = (inp[6]) ? node2508 : 15'b000000000111111;
													assign node2508 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2512 = (inp[14]) ? node2534 : node2513;
									assign node2513 = (inp[4]) ? node2521 : node2514;
										assign node2514 = (inp[0]) ? node2516 : 15'b000000111111111;
											assign node2516 = (inp[9]) ? 15'b000000000111111 : node2517;
												assign node2517 = (inp[6]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node2521 = (inp[3]) ? node2529 : node2522;
											assign node2522 = (inp[2]) ? 15'b000000000111111 : node2523;
												assign node2523 = (inp[7]) ? node2525 : 15'b000000001111111;
													assign node2525 = (inp[6]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node2529 = (inp[7]) ? 15'b000000000001111 : node2530;
												assign node2530 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2534 = (inp[6]) ? node2544 : node2535;
										assign node2535 = (inp[4]) ? node2539 : node2536;
											assign node2536 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2539 = (inp[3]) ? node2541 : 15'b000000000111111;
												assign node2541 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node2544 = (inp[4]) ? 15'b000000000001111 : node2545;
											assign node2545 = (inp[3]) ? node2547 : 15'b000000000011111;
												assign node2547 = (inp[7]) ? 15'b000000000000111 : 15'b000000000011111;
					assign node2551 = (inp[2]) ? node2719 : node2552;
						assign node2552 = (inp[14]) ? node2642 : node2553;
							assign node2553 = (inp[7]) ? node2611 : node2554;
								assign node2554 = (inp[3]) ? node2586 : node2555;
									assign node2555 = (inp[0]) ? node2573 : node2556;
										assign node2556 = (inp[8]) ? node2562 : node2557;
											assign node2557 = (inp[9]) ? node2559 : 15'b000001111111111;
												assign node2559 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2562 = (inp[11]) ? node2568 : node2563;
												assign node2563 = (inp[5]) ? 15'b000000111111111 : node2564;
													assign node2564 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2568 = (inp[9]) ? 15'b000000011111111 : node2569;
													assign node2569 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2573 = (inp[11]) ? node2583 : node2574;
											assign node2574 = (inp[6]) ? 15'b000000011111111 : node2575;
												assign node2575 = (inp[8]) ? 15'b000000011111111 : node2576;
													assign node2576 = (inp[4]) ? 15'b000000111111111 : node2577;
														assign node2577 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2583 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2586 = (inp[8]) ? node2598 : node2587;
										assign node2587 = (inp[0]) ? node2591 : node2588;
											assign node2588 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2591 = (inp[6]) ? 15'b000000001111111 : node2592;
												assign node2592 = (inp[9]) ? 15'b000000011111111 : node2593;
													assign node2593 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2598 = (inp[4]) ? node2600 : 15'b000000011111111;
											assign node2600 = (inp[11]) ? node2604 : node2601;
												assign node2601 = (inp[9]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node2604 = (inp[0]) ? 15'b000000000011111 : node2605;
													assign node2605 = (inp[6]) ? node2607 : 15'b000000001111111;
														assign node2607 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2611 = (inp[8]) ? node2625 : node2612;
									assign node2612 = (inp[4]) ? node2618 : node2613;
										assign node2613 = (inp[6]) ? 15'b000001111111111 : node2614;
											assign node2614 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2618 = (inp[0]) ? node2622 : node2619;
											assign node2619 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node2622 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2625 = (inp[6]) ? node2631 : node2626;
										assign node2626 = (inp[9]) ? 15'b000000000111111 : node2627;
											assign node2627 = (inp[5]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node2631 = (inp[0]) ? node2637 : node2632;
											assign node2632 = (inp[4]) ? node2634 : 15'b000000000111111;
												assign node2634 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2637 = (inp[4]) ? 15'b000000000011111 : node2638;
												assign node2638 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node2642 = (inp[5]) ? node2682 : node2643;
								assign node2643 = (inp[11]) ? node2665 : node2644;
									assign node2644 = (inp[6]) ? node2652 : node2645;
										assign node2645 = (inp[0]) ? node2649 : node2646;
											assign node2646 = (inp[8]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node2649 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2652 = (inp[9]) ? node2656 : node2653;
											assign node2653 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2656 = (inp[4]) ? 15'b000000000111111 : node2657;
												assign node2657 = (inp[3]) ? node2659 : 15'b000000011111111;
													assign node2659 = (inp[0]) ? node2661 : 15'b000000001111111;
														assign node2661 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2665 = (inp[8]) ? node2675 : node2666;
										assign node2666 = (inp[3]) ? 15'b000000000111111 : node2667;
											assign node2667 = (inp[6]) ? 15'b000000001111111 : node2668;
												assign node2668 = (inp[0]) ? 15'b000000011111111 : node2669;
													assign node2669 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2675 = (inp[9]) ? node2679 : node2676;
											assign node2676 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node2679 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2682 = (inp[9]) ? node2698 : node2683;
									assign node2683 = (inp[0]) ? node2693 : node2684;
										assign node2684 = (inp[8]) ? node2690 : node2685;
											assign node2685 = (inp[4]) ? node2687 : 15'b000000111111111;
												assign node2687 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node2690 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node2693 = (inp[4]) ? 15'b000000000111111 : node2694;
											assign node2694 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node2698 = (inp[0]) ? node2708 : node2699;
										assign node2699 = (inp[6]) ? node2703 : node2700;
											assign node2700 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node2703 = (inp[4]) ? node2705 : 15'b000000000111111;
												assign node2705 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2708 = (inp[7]) ? node2716 : node2709;
											assign node2709 = (inp[6]) ? 15'b000000000000111 : node2710;
												assign node2710 = (inp[8]) ? 15'b000000000011111 : node2711;
													assign node2711 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2716 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node2719 = (inp[4]) ? node2811 : node2720;
							assign node2720 = (inp[8]) ? node2778 : node2721;
								assign node2721 = (inp[7]) ? node2747 : node2722;
									assign node2722 = (inp[0]) ? node2732 : node2723;
										assign node2723 = (inp[11]) ? node2727 : node2724;
											assign node2724 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2727 = (inp[5]) ? node2729 : 15'b000000011111111;
												assign node2729 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2732 = (inp[11]) ? node2742 : node2733;
											assign node2733 = (inp[6]) ? node2735 : 15'b000000111111111;
												assign node2735 = (inp[3]) ? node2737 : 15'b000000011111111;
													assign node2737 = (inp[14]) ? 15'b000000001111111 : node2738;
														assign node2738 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2742 = (inp[3]) ? node2744 : 15'b000000001111111;
												assign node2744 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2747 = (inp[14]) ? node2761 : node2748;
										assign node2748 = (inp[5]) ? 15'b000000000111111 : node2749;
											assign node2749 = (inp[11]) ? node2753 : node2750;
												assign node2750 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2753 = (inp[0]) ? node2755 : 15'b000000001111111;
													assign node2755 = (inp[6]) ? node2757 : 15'b000000001111111;
														assign node2757 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2761 = (inp[6]) ? node2767 : node2762;
											assign node2762 = (inp[11]) ? 15'b000000000111111 : node2763;
												assign node2763 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2767 = (inp[9]) ? node2769 : 15'b000000000111111;
												assign node2769 = (inp[0]) ? node2775 : node2770;
													assign node2770 = (inp[3]) ? 15'b000000000011111 : node2771;
														assign node2771 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node2775 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node2778 = (inp[11]) ? node2798 : node2779;
									assign node2779 = (inp[14]) ? node2789 : node2780;
										assign node2780 = (inp[6]) ? node2786 : node2781;
											assign node2781 = (inp[7]) ? node2783 : 15'b000000001111111;
												assign node2783 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2786 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2789 = (inp[5]) ? node2791 : 15'b000000000011111;
											assign node2791 = (inp[6]) ? 15'b000000000111111 : node2792;
												assign node2792 = (inp[3]) ? 15'b000000000111111 : node2793;
													assign node2793 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2798 = (inp[9]) ? node2802 : node2799;
										assign node2799 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node2802 = (inp[5]) ? node2806 : node2803;
											assign node2803 = (inp[3]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node2806 = (inp[0]) ? 15'b000000000001111 : node2807;
												assign node2807 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node2811 = (inp[0]) ? node2871 : node2812;
								assign node2812 = (inp[6]) ? node2850 : node2813;
									assign node2813 = (inp[3]) ? node2833 : node2814;
										assign node2814 = (inp[5]) ? node2822 : node2815;
											assign node2815 = (inp[7]) ? 15'b000000001111111 : node2816;
												assign node2816 = (inp[9]) ? node2818 : 15'b000000111111111;
													assign node2818 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2822 = (inp[9]) ? node2828 : node2823;
												assign node2823 = (inp[11]) ? 15'b000000001111111 : node2824;
													assign node2824 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2828 = (inp[7]) ? 15'b000000000111111 : node2829;
													assign node2829 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2833 = (inp[9]) ? node2847 : node2834;
											assign node2834 = (inp[14]) ? node2842 : node2835;
												assign node2835 = (inp[7]) ? node2839 : node2836;
													assign node2836 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2839 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2842 = (inp[11]) ? 15'b000000000011111 : node2843;
													assign node2843 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2847 = (inp[11]) ? 15'b000000000011111 : 15'b000000000001111;
									assign node2850 = (inp[14]) ? node2856 : node2851;
										assign node2851 = (inp[7]) ? 15'b000000000111111 : node2852;
											assign node2852 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node2856 = (inp[9]) ? node2862 : node2857;
											assign node2857 = (inp[11]) ? 15'b000000000011111 : node2858;
												assign node2858 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2862 = (inp[8]) ? 15'b000000000000111 : node2863;
												assign node2863 = (inp[7]) ? node2867 : node2864;
													assign node2864 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node2867 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node2871 = (inp[14]) ? node2889 : node2872;
									assign node2872 = (inp[5]) ? node2882 : node2873;
										assign node2873 = (inp[11]) ? 15'b000000000011111 : node2874;
											assign node2874 = (inp[9]) ? 15'b000000000111111 : node2875;
												assign node2875 = (inp[8]) ? 15'b000000000111111 : node2876;
													assign node2876 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2882 = (inp[7]) ? node2884 : 15'b000000000011111;
											assign node2884 = (inp[11]) ? 15'b000000000001111 : node2885;
												assign node2885 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node2889 = (inp[8]) ? node2903 : node2890;
										assign node2890 = (inp[6]) ? node2896 : node2891;
											assign node2891 = (inp[3]) ? 15'b000000000011111 : node2892;
												assign node2892 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2896 = (inp[9]) ? node2900 : node2897;
												assign node2897 = (inp[5]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node2900 = (inp[3]) ? 15'b000000000001111 : 15'b000000000000111;
										assign node2903 = (inp[9]) ? node2907 : node2904;
											assign node2904 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node2907 = (inp[6]) ? node2911 : node2908;
												assign node2908 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node2911 = (inp[3]) ? 15'b000000000000111 : node2912;
													assign node2912 = (inp[11]) ? 15'b000000000000011 : 15'b000000000000111;
		assign node2916 = (inp[2]) ? node4368 : node2917;
			assign node2917 = (inp[14]) ? node3667 : node2918;
				assign node2918 = (inp[1]) ? node3308 : node2919;
					assign node2919 = (inp[9]) ? node3109 : node2920;
						assign node2920 = (inp[11]) ? node3022 : node2921;
							assign node2921 = (inp[10]) ? node2967 : node2922;
								assign node2922 = (inp[13]) ? node2948 : node2923;
									assign node2923 = (inp[3]) ? node2933 : node2924;
										assign node2924 = (inp[5]) ? 15'b000011111111111 : node2925;
											assign node2925 = (inp[4]) ? node2927 : 15'b001111111111111;
												assign node2927 = (inp[0]) ? 15'b000111111111111 : node2928;
													assign node2928 = (inp[8]) ? 15'b000111111111111 : 15'b001111111111111;
										assign node2933 = (inp[6]) ? node2941 : node2934;
											assign node2934 = (inp[8]) ? node2938 : node2935;
												assign node2935 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2938 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2941 = (inp[7]) ? node2945 : node2942;
												assign node2942 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2945 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node2948 = (inp[0]) ? node2964 : node2949;
										assign node2949 = (inp[4]) ? node2959 : node2950;
											assign node2950 = (inp[7]) ? 15'b000001111111111 : node2951;
												assign node2951 = (inp[3]) ? node2953 : 15'b000111111111111;
													assign node2953 = (inp[6]) ? node2955 : 15'b000011111111111;
														assign node2955 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2959 = (inp[3]) ? node2961 : 15'b000001111111111;
												assign node2961 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2964 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node2967 = (inp[7]) ? node2997 : node2968;
									assign node2968 = (inp[3]) ? node2982 : node2969;
										assign node2969 = (inp[8]) ? node2977 : node2970;
											assign node2970 = (inp[0]) ? node2972 : 15'b000111111111111;
												assign node2972 = (inp[6]) ? 15'b000001111111111 : node2973;
													assign node2973 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2977 = (inp[4]) ? node2979 : 15'b000001111111111;
												assign node2979 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2982 = (inp[0]) ? node2992 : node2983;
											assign node2983 = (inp[6]) ? node2985 : 15'b000001111111111;
												assign node2985 = (inp[8]) ? node2987 : 15'b000001111111111;
													assign node2987 = (inp[5]) ? 15'b000000111111111 : node2988;
														assign node2988 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2992 = (inp[13]) ? 15'b000000111111111 : node2993;
												assign node2993 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2997 = (inp[5]) ? node3011 : node2998;
										assign node2998 = (inp[6]) ? node3004 : node2999;
											assign node2999 = (inp[8]) ? 15'b000000011111111 : node3000;
												assign node3000 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node3004 = (inp[3]) ? node3006 : 15'b000000111111111;
												assign node3006 = (inp[13]) ? 15'b000000011111111 : node3007;
													assign node3007 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3011 = (inp[6]) ? 15'b000000001111111 : node3012;
											assign node3012 = (inp[3]) ? 15'b000000001111111 : node3013;
												assign node3013 = (inp[0]) ? node3015 : 15'b000000111111111;
													assign node3015 = (inp[13]) ? 15'b000000011111111 : node3016;
														assign node3016 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node3022 = (inp[6]) ? node3060 : node3023;
								assign node3023 = (inp[13]) ? node3043 : node3024;
									assign node3024 = (inp[7]) ? node3030 : node3025;
										assign node3025 = (inp[3]) ? node3027 : 15'b000011111111111;
											assign node3027 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3030 = (inp[5]) ? 15'b000000111111111 : node3031;
											assign node3031 = (inp[10]) ? node3033 : 15'b000001111111111;
												assign node3033 = (inp[3]) ? node3035 : 15'b000001111111111;
													assign node3035 = (inp[8]) ? 15'b000000111111111 : node3036;
														assign node3036 = (inp[0]) ? 15'b000000111111111 : node3037;
															assign node3037 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node3043 = (inp[8]) ? node3053 : node3044;
										assign node3044 = (inp[5]) ? node3050 : node3045;
											assign node3045 = (inp[4]) ? node3047 : 15'b000001111111111;
												assign node3047 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3050 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3053 = (inp[7]) ? 15'b000000011111111 : node3054;
											assign node3054 = (inp[4]) ? node3056 : 15'b000000111111111;
												assign node3056 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node3060 = (inp[8]) ? node3090 : node3061;
									assign node3061 = (inp[4]) ? node3081 : node3062;
										assign node3062 = (inp[3]) ? node3070 : node3063;
											assign node3063 = (inp[7]) ? node3065 : 15'b000001111111111;
												assign node3065 = (inp[0]) ? 15'b000000111111111 : node3066;
													assign node3066 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3070 = (inp[5]) ? node3076 : node3071;
												assign node3071 = (inp[13]) ? node3073 : 15'b000000111111111;
													assign node3073 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3076 = (inp[0]) ? node3078 : 15'b000000011111111;
													assign node3078 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3081 = (inp[0]) ? node3085 : node3082;
											assign node3082 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3085 = (inp[3]) ? node3087 : 15'b000000000111111;
												assign node3087 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3090 = (inp[10]) ? node3098 : node3091;
										assign node3091 = (inp[13]) ? 15'b000000001111111 : node3092;
											assign node3092 = (inp[7]) ? node3094 : 15'b000011111111111;
												assign node3094 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3098 = (inp[3]) ? node3102 : node3099;
											assign node3099 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3102 = (inp[5]) ? node3104 : 15'b000000001111111;
												assign node3104 = (inp[13]) ? node3106 : 15'b000000000111111;
													assign node3106 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node3109 = (inp[13]) ? node3199 : node3110;
							assign node3110 = (inp[4]) ? node3162 : node3111;
								assign node3111 = (inp[11]) ? node3139 : node3112;
									assign node3112 = (inp[7]) ? node3128 : node3113;
										assign node3113 = (inp[6]) ? node3121 : node3114;
											assign node3114 = (inp[8]) ? 15'b000011111111111 : node3115;
												assign node3115 = (inp[5]) ? 15'b000011111111111 : node3116;
													assign node3116 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node3121 = (inp[5]) ? 15'b000000011111111 : node3122;
												assign node3122 = (inp[8]) ? node3124 : 15'b000011111111111;
													assign node3124 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3128 = (inp[6]) ? node3136 : node3129;
											assign node3129 = (inp[8]) ? 15'b000000111111111 : node3130;
												assign node3130 = (inp[3]) ? node3132 : 15'b000001111111111;
													assign node3132 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node3136 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3139 = (inp[10]) ? node3147 : node3140;
										assign node3140 = (inp[0]) ? node3144 : node3141;
											assign node3141 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3144 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3147 = (inp[7]) ? node3153 : node3148;
											assign node3148 = (inp[0]) ? node3150 : 15'b000000111111111;
												assign node3150 = (inp[8]) ? 15'b000000000111111 : 15'b000000111111111;
											assign node3153 = (inp[0]) ? node3159 : node3154;
												assign node3154 = (inp[6]) ? 15'b000000001111111 : node3155;
													assign node3155 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3159 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node3162 = (inp[5]) ? node3182 : node3163;
									assign node3163 = (inp[7]) ? node3171 : node3164;
										assign node3164 = (inp[8]) ? node3166 : 15'b000001111111111;
											assign node3166 = (inp[3]) ? node3168 : 15'b000001111111111;
												assign node3168 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3171 = (inp[3]) ? node3177 : node3172;
											assign node3172 = (inp[0]) ? node3174 : 15'b000000111111111;
												assign node3174 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3177 = (inp[11]) ? 15'b000000001111111 : node3178;
												assign node3178 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3182 = (inp[10]) ? node3190 : node3183;
										assign node3183 = (inp[8]) ? node3187 : node3184;
											assign node3184 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3187 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3190 = (inp[0]) ? 15'b000000000011111 : node3191;
											assign node3191 = (inp[7]) ? node3193 : 15'b000000011111111;
												assign node3193 = (inp[11]) ? node3195 : 15'b000000001111111;
													assign node3195 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node3199 = (inp[0]) ? node3257 : node3200;
								assign node3200 = (inp[4]) ? node3228 : node3201;
									assign node3201 = (inp[5]) ? node3217 : node3202;
										assign node3202 = (inp[11]) ? node3208 : node3203;
											assign node3203 = (inp[3]) ? node3205 : 15'b000000111111111;
												assign node3205 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3208 = (inp[3]) ? 15'b000000011111111 : node3209;
												assign node3209 = (inp[7]) ? node3211 : 15'b000000111111111;
													assign node3211 = (inp[10]) ? 15'b000000011111111 : node3212;
														assign node3212 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3217 = (inp[6]) ? node3223 : node3218;
											assign node3218 = (inp[10]) ? 15'b000000011111111 : node3219;
												assign node3219 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3223 = (inp[7]) ? 15'b000000001111111 : node3224;
												assign node3224 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3228 = (inp[10]) ? node3240 : node3229;
										assign node3229 = (inp[5]) ? node3233 : node3230;
											assign node3230 = (inp[11]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node3233 = (inp[11]) ? node3235 : 15'b000000011111111;
												assign node3235 = (inp[8]) ? 15'b000000000111111 : node3236;
													assign node3236 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3240 = (inp[3]) ? node3250 : node3241;
											assign node3241 = (inp[11]) ? node3243 : 15'b000000011111111;
												assign node3243 = (inp[5]) ? node3247 : node3244;
													assign node3244 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3247 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3250 = (inp[8]) ? node3252 : 15'b000000001111111;
												assign node3252 = (inp[11]) ? node3254 : 15'b000000000111111;
													assign node3254 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3257 = (inp[7]) ? node3279 : node3258;
									assign node3258 = (inp[5]) ? node3266 : node3259;
										assign node3259 = (inp[8]) ? node3263 : node3260;
											assign node3260 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node3263 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3266 = (inp[11]) ? node3272 : node3267;
											assign node3267 = (inp[4]) ? 15'b000000001111111 : node3268;
												assign node3268 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3272 = (inp[3]) ? 15'b000000000111111 : node3273;
												assign node3273 = (inp[10]) ? node3275 : 15'b000000001111111;
													assign node3275 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node3279 = (inp[4]) ? node3297 : node3280;
										assign node3280 = (inp[10]) ? node3292 : node3281;
											assign node3281 = (inp[5]) ? node3289 : node3282;
												assign node3282 = (inp[11]) ? 15'b000000001111111 : node3283;
													assign node3283 = (inp[8]) ? node3285 : 15'b000000011111111;
														assign node3285 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3289 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3292 = (inp[6]) ? node3294 : 15'b000000001111111;
												assign node3294 = (inp[5]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node3297 = (inp[6]) ? node3305 : node3298;
											assign node3298 = (inp[11]) ? node3300 : 15'b000000001111111;
												assign node3300 = (inp[3]) ? 15'b000000000111111 : node3301;
													assign node3301 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3305 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node3308 = (inp[7]) ? node3478 : node3309;
						assign node3309 = (inp[6]) ? node3381 : node3310;
							assign node3310 = (inp[11]) ? node3350 : node3311;
								assign node3311 = (inp[0]) ? node3333 : node3312;
									assign node3312 = (inp[4]) ? node3318 : node3313;
										assign node3313 = (inp[13]) ? node3315 : 15'b000001111111111;
											assign node3315 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node3318 = (inp[3]) ? 15'b000000111111111 : node3319;
											assign node3319 = (inp[10]) ? node3325 : node3320;
												assign node3320 = (inp[13]) ? node3322 : 15'b000001111111111;
													assign node3322 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3325 = (inp[13]) ? node3329 : node3326;
													assign node3326 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3329 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3333 = (inp[4]) ? node3341 : node3334;
										assign node3334 = (inp[10]) ? node3338 : node3335;
											assign node3335 = (inp[9]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node3338 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3341 = (inp[9]) ? node3343 : 15'b000000111111111;
											assign node3343 = (inp[13]) ? 15'b000000001111111 : node3344;
												assign node3344 = (inp[3]) ? 15'b000000011111111 : node3345;
													assign node3345 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node3350 = (inp[8]) ? node3364 : node3351;
									assign node3351 = (inp[3]) ? node3357 : node3352;
										assign node3352 = (inp[0]) ? 15'b000000111111111 : node3353;
											assign node3353 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3357 = (inp[9]) ? 15'b000000011111111 : node3358;
											assign node3358 = (inp[4]) ? node3360 : 15'b000000111111111;
												assign node3360 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3364 = (inp[5]) ? node3374 : node3365;
										assign node3365 = (inp[10]) ? node3369 : node3366;
											assign node3366 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3369 = (inp[4]) ? node3371 : 15'b000000011111111;
												assign node3371 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3374 = (inp[9]) ? 15'b000000000011111 : node3375;
											assign node3375 = (inp[10]) ? 15'b000000001111111 : node3376;
												assign node3376 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
							assign node3381 = (inp[13]) ? node3421 : node3382;
								assign node3382 = (inp[0]) ? node3400 : node3383;
									assign node3383 = (inp[8]) ? node3393 : node3384;
										assign node3384 = (inp[5]) ? 15'b000000111111111 : node3385;
											assign node3385 = (inp[11]) ? node3387 : 15'b000001111111111;
												assign node3387 = (inp[10]) ? 15'b000000111111111 : node3388;
													assign node3388 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3393 = (inp[3]) ? 15'b000000001111111 : node3394;
											assign node3394 = (inp[11]) ? 15'b000000011111111 : node3395;
												assign node3395 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3400 = (inp[10]) ? node3410 : node3401;
										assign node3401 = (inp[5]) ? node3403 : 15'b000000111111111;
											assign node3403 = (inp[11]) ? node3405 : 15'b000000011111111;
												assign node3405 = (inp[4]) ? 15'b000000001111111 : node3406;
													assign node3406 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3410 = (inp[4]) ? node3416 : node3411;
											assign node3411 = (inp[5]) ? 15'b000000001111111 : node3412;
												assign node3412 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3416 = (inp[11]) ? node3418 : 15'b000000001111111;
												assign node3418 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3421 = (inp[3]) ? node3445 : node3422;
									assign node3422 = (inp[0]) ? node3436 : node3423;
										assign node3423 = (inp[11]) ? node3431 : node3424;
											assign node3424 = (inp[10]) ? node3426 : 15'b000000111111111;
												assign node3426 = (inp[4]) ? 15'b000000011111111 : node3427;
													assign node3427 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node3431 = (inp[9]) ? node3433 : 15'b000000011111111;
												assign node3433 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node3436 = (inp[9]) ? node3440 : node3437;
											assign node3437 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3440 = (inp[10]) ? node3442 : 15'b000000001111111;
												assign node3442 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3445 = (inp[10]) ? node3463 : node3446;
										assign node3446 = (inp[8]) ? node3450 : node3447;
											assign node3447 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3450 = (inp[9]) ? node3458 : node3451;
												assign node3451 = (inp[0]) ? 15'b000000001111111 : node3452;
													assign node3452 = (inp[11]) ? 15'b000000001111111 : node3453;
														assign node3453 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3458 = (inp[4]) ? 15'b000000000111111 : node3459;
													assign node3459 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3463 = (inp[4]) ? node3469 : node3464;
											assign node3464 = (inp[5]) ? 15'b000000000011111 : node3465;
												assign node3465 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3469 = (inp[9]) ? node3475 : node3470;
												assign node3470 = (inp[11]) ? 15'b000000000111111 : node3471;
													assign node3471 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3475 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node3478 = (inp[3]) ? node3572 : node3479;
							assign node3479 = (inp[6]) ? node3517 : node3480;
								assign node3480 = (inp[4]) ? node3492 : node3481;
									assign node3481 = (inp[5]) ? 15'b000000001111111 : node3482;
										assign node3482 = (inp[0]) ? node3488 : node3483;
											assign node3483 = (inp[11]) ? node3485 : 15'b000001111111111;
												assign node3485 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node3488 = (inp[9]) ? 15'b000000011111111 : 15'b000011111111111;
									assign node3492 = (inp[8]) ? node3508 : node3493;
										assign node3493 = (inp[13]) ? node3505 : node3494;
											assign node3494 = (inp[0]) ? 15'b000000011111111 : node3495;
												assign node3495 = (inp[9]) ? 15'b000000011111111 : node3496;
													assign node3496 = (inp[11]) ? node3498 : 15'b000000111111111;
														assign node3498 = (inp[5]) ? node3500 : 15'b000000111111111;
															assign node3500 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3505 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3508 = (inp[11]) ? node3514 : node3509;
											assign node3509 = (inp[9]) ? node3511 : 15'b000000011111111;
												assign node3511 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3514 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3517 = (inp[10]) ? node3543 : node3518;
									assign node3518 = (inp[0]) ? node3530 : node3519;
										assign node3519 = (inp[5]) ? node3525 : node3520;
											assign node3520 = (inp[4]) ? 15'b000000111111111 : node3521;
												assign node3521 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3525 = (inp[8]) ? node3527 : 15'b000000011111111;
												assign node3527 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3530 = (inp[4]) ? node3534 : node3531;
											assign node3531 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node3534 = (inp[5]) ? node3538 : node3535;
												assign node3535 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3538 = (inp[9]) ? 15'b000000000111111 : node3539;
													assign node3539 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3543 = (inp[5]) ? node3559 : node3544;
										assign node3544 = (inp[4]) ? node3548 : node3545;
											assign node3545 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node3548 = (inp[13]) ? node3550 : 15'b000000001111111;
												assign node3550 = (inp[8]) ? 15'b000000000111111 : node3551;
													assign node3551 = (inp[9]) ? node3553 : 15'b000000001111111;
														assign node3553 = (inp[11]) ? 15'b000000000111111 : node3554;
															assign node3554 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3559 = (inp[0]) ? node3563 : node3560;
											assign node3560 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3563 = (inp[9]) ? node3565 : 15'b000000000111111;
												assign node3565 = (inp[11]) ? node3569 : node3566;
													assign node3566 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3569 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3572 = (inp[4]) ? node3632 : node3573;
								assign node3573 = (inp[11]) ? node3609 : node3574;
									assign node3574 = (inp[13]) ? node3590 : node3575;
										assign node3575 = (inp[10]) ? node3585 : node3576;
											assign node3576 = (inp[0]) ? node3580 : node3577;
												assign node3577 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3580 = (inp[5]) ? node3582 : 15'b000000011111111;
													assign node3582 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3585 = (inp[0]) ? 15'b000000001111111 : node3586;
												assign node3586 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3590 = (inp[8]) ? node3604 : node3591;
											assign node3591 = (inp[6]) ? node3597 : node3592;
												assign node3592 = (inp[10]) ? 15'b000000011111111 : node3593;
													assign node3593 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3597 = (inp[9]) ? node3599 : 15'b000000001111111;
													assign node3599 = (inp[0]) ? 15'b000000000111111 : node3600;
														assign node3600 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3604 = (inp[9]) ? 15'b000000000111111 : node3605;
												assign node3605 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3609 = (inp[10]) ? node3621 : node3610;
										assign node3610 = (inp[0]) ? node3616 : node3611;
											assign node3611 = (inp[8]) ? node3613 : 15'b000000011111111;
												assign node3613 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node3616 = (inp[6]) ? 15'b000000000111111 : node3617;
												assign node3617 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node3621 = (inp[13]) ? node3627 : node3622;
											assign node3622 = (inp[6]) ? 15'b000000000111111 : node3623;
												assign node3623 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3627 = (inp[0]) ? 15'b000000000001111 : node3628;
												assign node3628 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node3632 = (inp[5]) ? node3642 : node3633;
									assign node3633 = (inp[10]) ? node3639 : node3634;
										assign node3634 = (inp[11]) ? node3636 : 15'b000000011111111;
											assign node3636 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3639 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3642 = (inp[13]) ? node3650 : node3643;
										assign node3643 = (inp[6]) ? 15'b000000000011111 : node3644;
											assign node3644 = (inp[11]) ? node3646 : 15'b000000001111111;
												assign node3646 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3650 = (inp[10]) ? node3658 : node3651;
											assign node3651 = (inp[11]) ? 15'b000000000011111 : node3652;
												assign node3652 = (inp[0]) ? node3654 : 15'b000000000111111;
													assign node3654 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node3658 = (inp[11]) ? node3662 : node3659;
												assign node3659 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node3662 = (inp[8]) ? node3664 : 15'b000000000011111;
													assign node3664 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node3667 = (inp[8]) ? node3997 : node3668;
					assign node3668 = (inp[6]) ? node3832 : node3669;
						assign node3669 = (inp[5]) ? node3749 : node3670;
							assign node3670 = (inp[7]) ? node3702 : node3671;
								assign node3671 = (inp[9]) ? node3695 : node3672;
									assign node3672 = (inp[0]) ? node3678 : node3673;
										assign node3673 = (inp[11]) ? 15'b000001111111111 : node3674;
											assign node3674 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node3678 = (inp[1]) ? node3686 : node3679;
											assign node3679 = (inp[10]) ? 15'b000000111111111 : node3680;
												assign node3680 = (inp[11]) ? node3682 : 15'b000001111111111;
													assign node3682 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3686 = (inp[3]) ? node3690 : node3687;
												assign node3687 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3690 = (inp[4]) ? node3692 : 15'b000000111111111;
													assign node3692 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3695 = (inp[11]) ? node3697 : 15'b000000111111111;
										assign node3697 = (inp[3]) ? 15'b000000011111111 : node3698;
											assign node3698 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node3702 = (inp[9]) ? node3724 : node3703;
									assign node3703 = (inp[1]) ? node3709 : node3704;
										assign node3704 = (inp[13]) ? node3706 : 15'b000001111111111;
											assign node3706 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3709 = (inp[0]) ? node3715 : node3710;
											assign node3710 = (inp[13]) ? node3712 : 15'b000000111111111;
												assign node3712 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3715 = (inp[13]) ? 15'b000000001111111 : node3716;
												assign node3716 = (inp[3]) ? node3720 : node3717;
													assign node3717 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3720 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3724 = (inp[0]) ? node3740 : node3725;
										assign node3725 = (inp[10]) ? node3731 : node3726;
											assign node3726 = (inp[3]) ? node3728 : 15'b000000111111111;
												assign node3728 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3731 = (inp[1]) ? node3737 : node3732;
												assign node3732 = (inp[11]) ? node3734 : 15'b000000111111111;
													assign node3734 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3737 = (inp[13]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node3740 = (inp[1]) ? node3744 : node3741;
											assign node3741 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3744 = (inp[11]) ? 15'b000000001111111 : node3745;
												assign node3745 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node3749 = (inp[13]) ? node3793 : node3750;
								assign node3750 = (inp[4]) ? node3774 : node3751;
									assign node3751 = (inp[10]) ? node3761 : node3752;
										assign node3752 = (inp[7]) ? 15'b000000111111111 : node3753;
											assign node3753 = (inp[11]) ? 15'b000000111111111 : node3754;
												assign node3754 = (inp[3]) ? node3756 : 15'b000001111111111;
													assign node3756 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node3761 = (inp[1]) ? node3765 : node3762;
											assign node3762 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3765 = (inp[11]) ? node3771 : node3766;
												assign node3766 = (inp[3]) ? 15'b000000011111111 : node3767;
													assign node3767 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3771 = (inp[3]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node3774 = (inp[11]) ? node3784 : node3775;
										assign node3775 = (inp[10]) ? node3779 : node3776;
											assign node3776 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3779 = (inp[3]) ? node3781 : 15'b000000011111111;
												assign node3781 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node3784 = (inp[1]) ? node3790 : node3785;
											assign node3785 = (inp[10]) ? 15'b000000001111111 : node3786;
												assign node3786 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3790 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3793 = (inp[3]) ? node3807 : node3794;
									assign node3794 = (inp[1]) ? node3802 : node3795;
										assign node3795 = (inp[0]) ? 15'b000000011111111 : node3796;
											assign node3796 = (inp[7]) ? node3798 : 15'b000000111111111;
												assign node3798 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3802 = (inp[4]) ? 15'b000000000111111 : node3803;
											assign node3803 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3807 = (inp[1]) ? node3821 : node3808;
										assign node3808 = (inp[7]) ? node3818 : node3809;
											assign node3809 = (inp[11]) ? node3811 : 15'b000000011111111;
												assign node3811 = (inp[0]) ? node3815 : node3812;
													assign node3812 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3815 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node3818 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3821 = (inp[11]) ? node3825 : node3822;
											assign node3822 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3825 = (inp[0]) ? node3827 : 15'b000000000111111;
												assign node3827 = (inp[9]) ? node3829 : 15'b000000000011111;
													assign node3829 = (inp[10]) ? 15'b000000000011111 : 15'b000000000001111;
						assign node3832 = (inp[0]) ? node3920 : node3833;
							assign node3833 = (inp[7]) ? node3875 : node3834;
								assign node3834 = (inp[9]) ? node3856 : node3835;
									assign node3835 = (inp[1]) ? node3849 : node3836;
										assign node3836 = (inp[3]) ? node3840 : node3837;
											assign node3837 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3840 = (inp[4]) ? node3842 : 15'b000000111111111;
												assign node3842 = (inp[5]) ? 15'b000000001111111 : node3843;
													assign node3843 = (inp[11]) ? 15'b000000011111111 : node3844;
														assign node3844 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3849 = (inp[5]) ? 15'b000000011111111 : node3850;
											assign node3850 = (inp[10]) ? 15'b000000011111111 : node3851;
												assign node3851 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3856 = (inp[4]) ? node3866 : node3857;
										assign node3857 = (inp[5]) ? node3861 : node3858;
											assign node3858 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3861 = (inp[13]) ? node3863 : 15'b000000011111111;
												assign node3863 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3866 = (inp[13]) ? node3872 : node3867;
											assign node3867 = (inp[11]) ? 15'b000000001111111 : node3868;
												assign node3868 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3872 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node3875 = (inp[5]) ? node3893 : node3876;
									assign node3876 = (inp[1]) ? node3886 : node3877;
										assign node3877 = (inp[13]) ? node3883 : node3878;
											assign node3878 = (inp[9]) ? node3880 : 15'b000000111111111;
												assign node3880 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3883 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3886 = (inp[11]) ? node3890 : node3887;
											assign node3887 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3890 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node3893 = (inp[1]) ? node3909 : node3894;
										assign node3894 = (inp[4]) ? node3898 : node3895;
											assign node3895 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3898 = (inp[11]) ? node3902 : node3899;
												assign node3899 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3902 = (inp[9]) ? 15'b000000000111111 : node3903;
													assign node3903 = (inp[13]) ? node3905 : 15'b000000001111111;
														assign node3905 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3909 = (inp[10]) ? node3915 : node3910;
											assign node3910 = (inp[4]) ? node3912 : 15'b000000001111111;
												assign node3912 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3915 = (inp[9]) ? node3917 : 15'b000000000111111;
												assign node3917 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3920 = (inp[10]) ? node3956 : node3921;
								assign node3921 = (inp[9]) ? node3947 : node3922;
									assign node3922 = (inp[13]) ? node3936 : node3923;
										assign node3923 = (inp[3]) ? node3929 : node3924;
											assign node3924 = (inp[11]) ? 15'b000000001111111 : node3925;
												assign node3925 = (inp[5]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node3929 = (inp[7]) ? 15'b000000001111111 : node3930;
												assign node3930 = (inp[5]) ? node3932 : 15'b000000011111111;
													assign node3932 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3936 = (inp[4]) ? node3942 : node3937;
											assign node3937 = (inp[7]) ? 15'b000000000111111 : node3938;
												assign node3938 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3942 = (inp[1]) ? 15'b000000000111111 : node3943;
												assign node3943 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3947 = (inp[1]) ? node3953 : node3948;
										assign node3948 = (inp[13]) ? node3950 : 15'b000000000111111;
											assign node3950 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3953 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3956 = (inp[11]) ? node3980 : node3957;
									assign node3957 = (inp[4]) ? node3969 : node3958;
										assign node3958 = (inp[1]) ? node3962 : node3959;
											assign node3959 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3962 = (inp[7]) ? node3964 : 15'b000000001111111;
												assign node3964 = (inp[13]) ? 15'b000000000111111 : node3965;
													assign node3965 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3969 = (inp[3]) ? node3973 : node3970;
											assign node3970 = (inp[9]) ? 15'b000000000011111 : 15'b000000011111111;
											assign node3973 = (inp[9]) ? node3975 : 15'b000000000111111;
												assign node3975 = (inp[7]) ? node3977 : 15'b000000000111111;
													assign node3977 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3980 = (inp[3]) ? node3990 : node3981;
										assign node3981 = (inp[13]) ? node3987 : node3982;
											assign node3982 = (inp[5]) ? 15'b000000000111111 : node3983;
												assign node3983 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3987 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3990 = (inp[4]) ? node3994 : node3991;
											assign node3991 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3994 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node3997 = (inp[3]) ? node4187 : node3998;
						assign node3998 = (inp[6]) ? node4110 : node3999;
							assign node3999 = (inp[7]) ? node4053 : node4000;
								assign node4000 = (inp[11]) ? node4022 : node4001;
									assign node4001 = (inp[13]) ? node4015 : node4002;
										assign node4002 = (inp[10]) ? node4004 : 15'b000000111111111;
											assign node4004 = (inp[1]) ? node4010 : node4005;
												assign node4005 = (inp[0]) ? 15'b000000011111111 : node4006;
													assign node4006 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4010 = (inp[0]) ? node4012 : 15'b000000011111111;
													assign node4012 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4015 = (inp[0]) ? 15'b000000011111111 : node4016;
											assign node4016 = (inp[9]) ? node4018 : 15'b000000111111111;
												assign node4018 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4022 = (inp[5]) ? node4036 : node4023;
										assign node4023 = (inp[9]) ? node4029 : node4024;
											assign node4024 = (inp[13]) ? 15'b000000111111111 : node4025;
												assign node4025 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4029 = (inp[0]) ? node4031 : 15'b000000111111111;
												assign node4031 = (inp[10]) ? 15'b000000000111111 : node4032;
													assign node4032 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4036 = (inp[1]) ? node4042 : node4037;
											assign node4037 = (inp[10]) ? node4039 : 15'b000000011111111;
												assign node4039 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4042 = (inp[10]) ? node4048 : node4043;
												assign node4043 = (inp[4]) ? 15'b000000001111111 : node4044;
													assign node4044 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4048 = (inp[13]) ? 15'b000000000111111 : node4049;
													assign node4049 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
								assign node4053 = (inp[9]) ? node4079 : node4054;
									assign node4054 = (inp[13]) ? node4068 : node4055;
										assign node4055 = (inp[1]) ? node4061 : node4056;
											assign node4056 = (inp[5]) ? 15'b000000011111111 : node4057;
												assign node4057 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4061 = (inp[11]) ? 15'b000000001111111 : node4062;
												assign node4062 = (inp[0]) ? node4064 : 15'b000000011111111;
													assign node4064 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4068 = (inp[11]) ? node4076 : node4069;
											assign node4069 = (inp[1]) ? node4071 : 15'b000000001111111;
												assign node4071 = (inp[5]) ? node4073 : 15'b000000001111111;
													assign node4073 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4076 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4079 = (inp[1]) ? node4093 : node4080;
										assign node4080 = (inp[4]) ? node4084 : node4081;
											assign node4081 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4084 = (inp[10]) ? 15'b000000000111111 : node4085;
												assign node4085 = (inp[0]) ? node4089 : node4086;
													assign node4086 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4089 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4093 = (inp[0]) ? node4103 : node4094;
											assign node4094 = (inp[11]) ? node4098 : node4095;
												assign node4095 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4098 = (inp[13]) ? 15'b000000000011111 : node4099;
													assign node4099 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4103 = (inp[13]) ? node4105 : 15'b000000000111111;
												assign node4105 = (inp[11]) ? 15'b000000000011111 : node4106;
													assign node4106 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node4110 = (inp[4]) ? node4144 : node4111;
								assign node4111 = (inp[13]) ? node4127 : node4112;
									assign node4112 = (inp[9]) ? node4118 : node4113;
										assign node4113 = (inp[5]) ? node4115 : 15'b000000011111111;
											assign node4115 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node4118 = (inp[1]) ? 15'b000000001111111 : node4119;
											assign node4119 = (inp[0]) ? 15'b000000001111111 : node4120;
												assign node4120 = (inp[5]) ? node4122 : 15'b000000011111111;
													assign node4122 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4127 = (inp[5]) ? node4137 : node4128;
										assign node4128 = (inp[1]) ? node4134 : node4129;
											assign node4129 = (inp[9]) ? node4131 : 15'b000000001111111;
												assign node4131 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4134 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node4137 = (inp[9]) ? node4141 : node4138;
											assign node4138 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4141 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node4144 = (inp[5]) ? node4160 : node4145;
									assign node4145 = (inp[10]) ? node4149 : node4146;
										assign node4146 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4149 = (inp[13]) ? node4157 : node4150;
											assign node4150 = (inp[7]) ? 15'b000000000111111 : node4151;
												assign node4151 = (inp[0]) ? node4153 : 15'b000000001111111;
													assign node4153 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4157 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4160 = (inp[0]) ? node4168 : node4161;
										assign node4161 = (inp[7]) ? node4165 : node4162;
											assign node4162 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4165 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4168 = (inp[1]) ? node4180 : node4169;
											assign node4169 = (inp[7]) ? node4175 : node4170;
												assign node4170 = (inp[13]) ? node4172 : 15'b000000000111111;
													assign node4172 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node4175 = (inp[13]) ? node4177 : 15'b000000000011111;
													assign node4177 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4180 = (inp[9]) ? node4182 : 15'b000000000011111;
												assign node4182 = (inp[7]) ? 15'b000000000000111 : node4183;
													assign node4183 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node4187 = (inp[13]) ? node4277 : node4188;
							assign node4188 = (inp[4]) ? node4234 : node4189;
								assign node4189 = (inp[11]) ? node4209 : node4190;
									assign node4190 = (inp[5]) ? node4198 : node4191;
										assign node4191 = (inp[6]) ? node4193 : 15'b000001111111111;
											assign node4193 = (inp[1]) ? 15'b000000001111111 : node4194;
												assign node4194 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4198 = (inp[6]) ? node4204 : node4199;
											assign node4199 = (inp[10]) ? 15'b000000001111111 : node4200;
												assign node4200 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4204 = (inp[7]) ? node4206 : 15'b000000001111111;
												assign node4206 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4209 = (inp[6]) ? node4225 : node4210;
										assign node4210 = (inp[0]) ? node4222 : node4211;
											assign node4211 = (inp[5]) ? node4215 : node4212;
												assign node4212 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4215 = (inp[10]) ? node4219 : node4216;
													assign node4216 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4219 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4222 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4225 = (inp[1]) ? node4229 : node4226;
											assign node4226 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4229 = (inp[7]) ? node4231 : 15'b000000000111111;
												assign node4231 = (inp[0]) ? 15'b000000000011111 : 15'b000000000001111;
								assign node4234 = (inp[10]) ? node4262 : node4235;
									assign node4235 = (inp[6]) ? node4241 : node4236;
										assign node4236 = (inp[7]) ? node4238 : 15'b000000001111111;
											assign node4238 = (inp[1]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node4241 = (inp[5]) ? node4251 : node4242;
											assign node4242 = (inp[11]) ? 15'b000000000111111 : node4243;
												assign node4243 = (inp[0]) ? node4245 : 15'b000000111111111;
													assign node4245 = (inp[9]) ? 15'b000000000111111 : node4246;
														assign node4246 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4251 = (inp[11]) ? node4259 : node4252;
												assign node4252 = (inp[9]) ? node4256 : node4253;
													assign node4253 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4256 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4259 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node4262 = (inp[6]) ? node4272 : node4263;
										assign node4263 = (inp[7]) ? node4267 : node4264;
											assign node4264 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4267 = (inp[0]) ? 15'b000000000011111 : node4268;
												assign node4268 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4272 = (inp[7]) ? node4274 : 15'b000000000011111;
											assign node4274 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node4277 = (inp[11]) ? node4309 : node4278;
								assign node4278 = (inp[0]) ? node4294 : node4279;
									assign node4279 = (inp[6]) ? node4285 : node4280;
										assign node4280 = (inp[4]) ? 15'b000000001111111 : node4281;
											assign node4281 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4285 = (inp[10]) ? node4291 : node4286;
											assign node4286 = (inp[1]) ? 15'b000000000111111 : node4287;
												assign node4287 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4291 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4294 = (inp[10]) ? node4302 : node4295;
										assign node4295 = (inp[4]) ? 15'b000000000111111 : node4296;
											assign node4296 = (inp[7]) ? node4298 : 15'b000000000111111;
												assign node4298 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4302 = (inp[5]) ? node4306 : node4303;
											assign node4303 = (inp[6]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node4306 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node4309 = (inp[4]) ? node4341 : node4310;
									assign node4310 = (inp[5]) ? node4324 : node4311;
										assign node4311 = (inp[7]) ? node4315 : node4312;
											assign node4312 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4315 = (inp[9]) ? 15'b000000000011111 : node4316;
												assign node4316 = (inp[0]) ? 15'b000000000011111 : node4317;
													assign node4317 = (inp[1]) ? node4319 : 15'b000000001111111;
														assign node4319 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4324 = (inp[7]) ? node4334 : node4325;
											assign node4325 = (inp[6]) ? 15'b000000000011111 : node4326;
												assign node4326 = (inp[1]) ? node4328 : 15'b000000000111111;
													assign node4328 = (inp[10]) ? 15'b000000000001111 : node4329;
														assign node4329 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4334 = (inp[0]) ? node4336 : 15'b000000000011111;
												assign node4336 = (inp[1]) ? 15'b000000000001111 : node4337;
													assign node4337 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node4341 = (inp[9]) ? node4349 : node4342;
										assign node4342 = (inp[5]) ? node4344 : 15'b000000000011111;
											assign node4344 = (inp[7]) ? 15'b000000000001111 : node4345;
												assign node4345 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4349 = (inp[0]) ? node4359 : node4350;
											assign node4350 = (inp[1]) ? node4352 : 15'b000000000011111;
												assign node4352 = (inp[5]) ? 15'b000000000001111 : node4353;
													assign node4353 = (inp[10]) ? 15'b000000000001111 : node4354;
														assign node4354 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4359 = (inp[5]) ? node4365 : node4360;
												assign node4360 = (inp[1]) ? node4362 : 15'b000000000001111;
													assign node4362 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node4365 = (inp[1]) ? 15'b000000000000011 : 15'b000000000000111;
			assign node4368 = (inp[10]) ? node5072 : node4369;
				assign node4369 = (inp[1]) ? node4709 : node4370;
					assign node4370 = (inp[6]) ? node4542 : node4371;
						assign node4371 = (inp[14]) ? node4463 : node4372;
							assign node4372 = (inp[7]) ? node4434 : node4373;
								assign node4373 = (inp[5]) ? node4407 : node4374;
									assign node4374 = (inp[9]) ? node4392 : node4375;
										assign node4375 = (inp[13]) ? node4387 : node4376;
											assign node4376 = (inp[11]) ? 15'b000001111111111 : node4377;
												assign node4377 = (inp[4]) ? 15'b000011111111111 : node4378;
													assign node4378 = (inp[3]) ? node4380 : 15'b000111111111111;
														assign node4380 = (inp[8]) ? 15'b000011111111111 : node4381;
															assign node4381 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node4387 = (inp[0]) ? 15'b000000111111111 : node4388;
												assign node4388 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node4392 = (inp[3]) ? node4404 : node4393;
											assign node4393 = (inp[13]) ? node4399 : node4394;
												assign node4394 = (inp[11]) ? node4396 : 15'b000001111111111;
													assign node4396 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4399 = (inp[4]) ? 15'b000000111111111 : node4400;
													assign node4400 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4404 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
									assign node4407 = (inp[9]) ? node4425 : node4408;
										assign node4408 = (inp[3]) ? node4414 : node4409;
											assign node4409 = (inp[13]) ? node4411 : 15'b000011111111111;
												assign node4411 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node4414 = (inp[13]) ? node4420 : node4415;
												assign node4415 = (inp[4]) ? 15'b000000111111111 : node4416;
													assign node4416 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4420 = (inp[0]) ? node4422 : 15'b000000111111111;
													assign node4422 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4425 = (inp[4]) ? node4431 : node4426;
											assign node4426 = (inp[13]) ? 15'b000000011111111 : node4427;
												assign node4427 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4431 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node4434 = (inp[0]) ? node4448 : node4435;
									assign node4435 = (inp[8]) ? node4445 : node4436;
										assign node4436 = (inp[3]) ? node4442 : node4437;
											assign node4437 = (inp[13]) ? node4439 : 15'b000001111111111;
												assign node4439 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4442 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node4445 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node4448 = (inp[11]) ? node4458 : node4449;
										assign node4449 = (inp[5]) ? node4451 : 15'b000001111111111;
											assign node4451 = (inp[13]) ? 15'b000000000111111 : node4452;
												assign node4452 = (inp[3]) ? 15'b000000011111111 : node4453;
													assign node4453 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node4458 = (inp[13]) ? 15'b000000000111111 : node4459;
											assign node4459 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
							assign node4463 = (inp[13]) ? node4509 : node4464;
								assign node4464 = (inp[11]) ? node4488 : node4465;
									assign node4465 = (inp[5]) ? node4479 : node4466;
										assign node4466 = (inp[3]) ? node4472 : node4467;
											assign node4467 = (inp[0]) ? 15'b000000111111111 : node4468;
												assign node4468 = (inp[8]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node4472 = (inp[4]) ? 15'b000000011111111 : node4473;
												assign node4473 = (inp[9]) ? node4475 : 15'b000000111111111;
													assign node4475 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4479 = (inp[3]) ? 15'b000000011111111 : node4480;
											assign node4480 = (inp[4]) ? node4482 : 15'b000000111111111;
												assign node4482 = (inp[0]) ? 15'b000000001111111 : node4483;
													assign node4483 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node4488 = (inp[7]) ? node4498 : node4489;
										assign node4489 = (inp[5]) ? node4493 : node4490;
											assign node4490 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node4493 = (inp[0]) ? node4495 : 15'b000000011111111;
												assign node4495 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node4498 = (inp[8]) ? 15'b000000000111111 : node4499;
											assign node4499 = (inp[3]) ? node4505 : node4500;
												assign node4500 = (inp[5]) ? node4502 : 15'b000000011111111;
													assign node4502 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4505 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
								assign node4509 = (inp[4]) ? node4527 : node4510;
									assign node4510 = (inp[8]) ? node4518 : node4511;
										assign node4511 = (inp[5]) ? node4515 : node4512;
											assign node4512 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4515 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node4518 = (inp[9]) ? 15'b000000001111111 : node4519;
											assign node4519 = (inp[0]) ? 15'b000000001111111 : node4520;
												assign node4520 = (inp[11]) ? node4522 : 15'b000000011111111;
													assign node4522 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4527 = (inp[7]) ? node4533 : node4528;
										assign node4528 = (inp[11]) ? node4530 : 15'b000000011111111;
											assign node4530 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node4533 = (inp[11]) ? node4537 : node4534;
											assign node4534 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4537 = (inp[8]) ? 15'b000000000001111 : node4538;
												assign node4538 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node4542 = (inp[3]) ? node4632 : node4543;
							assign node4543 = (inp[14]) ? node4591 : node4544;
								assign node4544 = (inp[8]) ? node4572 : node4545;
									assign node4545 = (inp[4]) ? node4563 : node4546;
										assign node4546 = (inp[9]) ? node4556 : node4547;
											assign node4547 = (inp[5]) ? node4553 : node4548;
												assign node4548 = (inp[7]) ? node4550 : 15'b000011111111111;
													assign node4550 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4553 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4556 = (inp[5]) ? 15'b000000000111111 : node4557;
												assign node4557 = (inp[13]) ? node4559 : 15'b000001111111111;
													assign node4559 = (inp[11]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node4563 = (inp[11]) ? 15'b000000011111111 : node4564;
											assign node4564 = (inp[9]) ? 15'b000000011111111 : node4565;
												assign node4565 = (inp[13]) ? node4567 : 15'b000000111111111;
													assign node4567 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node4572 = (inp[5]) ? node4580 : node4573;
										assign node4573 = (inp[11]) ? node4577 : node4574;
											assign node4574 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4577 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4580 = (inp[11]) ? 15'b000000000111111 : node4581;
											assign node4581 = (inp[4]) ? 15'b000000001111111 : node4582;
												assign node4582 = (inp[9]) ? 15'b000000001111111 : node4583;
													assign node4583 = (inp[0]) ? node4585 : 15'b000000011111111;
														assign node4585 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node4591 = (inp[4]) ? node4607 : node4592;
									assign node4592 = (inp[11]) ? node4600 : node4593;
										assign node4593 = (inp[0]) ? node4595 : 15'b000000111111111;
											assign node4595 = (inp[7]) ? node4597 : 15'b000000011111111;
												assign node4597 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node4600 = (inp[5]) ? node4602 : 15'b000000011111111;
											assign node4602 = (inp[0]) ? 15'b000000000011111 : node4603;
												assign node4603 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4607 = (inp[7]) ? node4619 : node4608;
										assign node4608 = (inp[13]) ? node4616 : node4609;
											assign node4609 = (inp[11]) ? 15'b000000001111111 : node4610;
												assign node4610 = (inp[8]) ? node4612 : 15'b000000011111111;
													assign node4612 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4616 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4619 = (inp[5]) ? node4625 : node4620;
											assign node4620 = (inp[13]) ? 15'b000000000111111 : node4621;
												assign node4621 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4625 = (inp[0]) ? node4627 : 15'b000000000111111;
												assign node4627 = (inp[9]) ? node4629 : 15'b000000000011111;
													assign node4629 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node4632 = (inp[7]) ? node4678 : node4633;
								assign node4633 = (inp[9]) ? node4655 : node4634;
									assign node4634 = (inp[13]) ? node4650 : node4635;
										assign node4635 = (inp[5]) ? node4641 : node4636;
											assign node4636 = (inp[14]) ? 15'b000000111111111 : node4637;
												assign node4637 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4641 = (inp[4]) ? node4645 : node4642;
												assign node4642 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4645 = (inp[8]) ? 15'b000000001111111 : node4646;
													assign node4646 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4650 = (inp[5]) ? node4652 : 15'b000000001111111;
											assign node4652 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4655 = (inp[5]) ? node4671 : node4656;
										assign node4656 = (inp[4]) ? node4664 : node4657;
											assign node4657 = (inp[0]) ? node4661 : node4658;
												assign node4658 = (inp[11]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node4661 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4664 = (inp[13]) ? 15'b000000000011111 : node4665;
												assign node4665 = (inp[11]) ? 15'b000000000111111 : node4666;
													assign node4666 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4671 = (inp[0]) ? node4673 : 15'b000000000111111;
											assign node4673 = (inp[8]) ? 15'b000000000011111 : node4674;
												assign node4674 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
								assign node4678 = (inp[5]) ? node4692 : node4679;
									assign node4679 = (inp[4]) ? node4683 : node4680;
										assign node4680 = (inp[11]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node4683 = (inp[13]) ? node4689 : node4684;
											assign node4684 = (inp[8]) ? 15'b000000000111111 : node4685;
												assign node4685 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4689 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4692 = (inp[4]) ? node4698 : node4693;
										assign node4693 = (inp[0]) ? 15'b000000000111111 : node4694;
											assign node4694 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node4698 = (inp[13]) ? node4700 : 15'b000000000011111;
											assign node4700 = (inp[14]) ? node4704 : node4701;
												assign node4701 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node4704 = (inp[9]) ? 15'b000000000001111 : node4705;
													assign node4705 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node4709 = (inp[6]) ? node4891 : node4710;
						assign node4710 = (inp[5]) ? node4794 : node4711;
							assign node4711 = (inp[11]) ? node4753 : node4712;
								assign node4712 = (inp[9]) ? node4736 : node4713;
									assign node4713 = (inp[0]) ? node4721 : node4714;
										assign node4714 = (inp[14]) ? 15'b000000111111111 : node4715;
											assign node4715 = (inp[3]) ? node4717 : 15'b000001111111111;
												assign node4717 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node4721 = (inp[7]) ? node4731 : node4722;
											assign node4722 = (inp[4]) ? node4728 : node4723;
												assign node4723 = (inp[3]) ? 15'b000000111111111 : node4724;
													assign node4724 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4728 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4731 = (inp[13]) ? node4733 : 15'b000000011111111;
												assign node4733 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node4736 = (inp[8]) ? node4746 : node4737;
										assign node4737 = (inp[4]) ? node4743 : node4738;
											assign node4738 = (inp[3]) ? 15'b000000011111111 : node4739;
												assign node4739 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4743 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node4746 = (inp[14]) ? node4750 : node4747;
											assign node4747 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4750 = (inp[0]) ? 15'b000000001111111 : 15'b000000000111111;
								assign node4753 = (inp[3]) ? node4773 : node4754;
									assign node4754 = (inp[14]) ? node4766 : node4755;
										assign node4755 = (inp[13]) ? node4759 : node4756;
											assign node4756 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4759 = (inp[0]) ? node4761 : 15'b000000011111111;
												assign node4761 = (inp[7]) ? 15'b000000001111111 : node4762;
													assign node4762 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4766 = (inp[9]) ? 15'b000000001111111 : node4767;
											assign node4767 = (inp[13]) ? 15'b000000001111111 : node4768;
												assign node4768 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4773 = (inp[0]) ? node4785 : node4774;
										assign node4774 = (inp[7]) ? 15'b000000000111111 : node4775;
											assign node4775 = (inp[13]) ? 15'b000000001111111 : node4776;
												assign node4776 = (inp[8]) ? node4778 : 15'b000000011111111;
													assign node4778 = (inp[14]) ? node4780 : 15'b000000011111111;
														assign node4780 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4785 = (inp[9]) ? node4791 : node4786;
											assign node4786 = (inp[14]) ? 15'b000000000111111 : node4787;
												assign node4787 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4791 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node4794 = (inp[8]) ? node4836 : node4795;
								assign node4795 = (inp[4]) ? node4817 : node4796;
									assign node4796 = (inp[7]) ? node4806 : node4797;
										assign node4797 = (inp[0]) ? node4801 : node4798;
											assign node4798 = (inp[13]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node4801 = (inp[14]) ? node4803 : 15'b000000011111111;
												assign node4803 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4806 = (inp[11]) ? node4812 : node4807;
											assign node4807 = (inp[14]) ? 15'b000000001111111 : node4808;
												assign node4808 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4812 = (inp[13]) ? node4814 : 15'b000000001111111;
												assign node4814 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4817 = (inp[3]) ? node4825 : node4818;
										assign node4818 = (inp[9]) ? 15'b000000000111111 : node4819;
											assign node4819 = (inp[0]) ? node4821 : 15'b000000011111111;
												assign node4821 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4825 = (inp[0]) ? node4827 : 15'b000000001111111;
											assign node4827 = (inp[11]) ? node4831 : node4828;
												assign node4828 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node4831 = (inp[13]) ? node4833 : 15'b000000000011111;
													assign node4833 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node4836 = (inp[11]) ? node4858 : node4837;
									assign node4837 = (inp[0]) ? node4845 : node4838;
										assign node4838 = (inp[4]) ? node4842 : node4839;
											assign node4839 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4842 = (inp[3]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node4845 = (inp[13]) ? node4851 : node4846;
											assign node4846 = (inp[4]) ? node4848 : 15'b000000001111111;
												assign node4848 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4851 = (inp[7]) ? node4853 : 15'b000000000111111;
												assign node4853 = (inp[3]) ? node4855 : 15'b000000000111111;
													assign node4855 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4858 = (inp[14]) ? node4876 : node4859;
										assign node4859 = (inp[0]) ? node4869 : node4860;
											assign node4860 = (inp[3]) ? node4866 : node4861;
												assign node4861 = (inp[13]) ? node4863 : 15'b000000011111111;
													assign node4863 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4866 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node4869 = (inp[13]) ? 15'b000000000001111 : node4870;
												assign node4870 = (inp[3]) ? node4872 : 15'b000000000111111;
													assign node4872 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4876 = (inp[13]) ? node4884 : node4877;
											assign node4877 = (inp[9]) ? node4879 : 15'b000000000111111;
												assign node4879 = (inp[0]) ? 15'b000000000011111 : node4880;
													assign node4880 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4884 = (inp[0]) ? 15'b000000000001111 : node4885;
												assign node4885 = (inp[9]) ? node4887 : 15'b000000000011111;
													assign node4887 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node4891 = (inp[0]) ? node4981 : node4892;
							assign node4892 = (inp[13]) ? node4930 : node4893;
								assign node4893 = (inp[7]) ? node4911 : node4894;
									assign node4894 = (inp[5]) ? node4902 : node4895;
										assign node4895 = (inp[8]) ? node4899 : node4896;
											assign node4896 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4899 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4902 = (inp[3]) ? node4908 : node4903;
											assign node4903 = (inp[11]) ? 15'b000000001111111 : node4904;
												assign node4904 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4908 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4911 = (inp[14]) ? node4923 : node4912;
										assign node4912 = (inp[11]) ? node4918 : node4913;
											assign node4913 = (inp[4]) ? node4915 : 15'b000000111111111;
												assign node4915 = (inp[5]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node4918 = (inp[8]) ? node4920 : 15'b000000001111111;
												assign node4920 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4923 = (inp[3]) ? 15'b000000000111111 : node4924;
											assign node4924 = (inp[8]) ? 15'b000000000111111 : node4925;
												assign node4925 = (inp[4]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node4930 = (inp[9]) ? node4948 : node4931;
									assign node4931 = (inp[5]) ? node4939 : node4932;
										assign node4932 = (inp[8]) ? node4934 : 15'b000000011111111;
											assign node4934 = (inp[14]) ? 15'b000000000111111 : node4935;
												assign node4935 = (inp[11]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node4939 = (inp[4]) ? node4945 : node4940;
											assign node4940 = (inp[7]) ? node4942 : 15'b000000001111111;
												assign node4942 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4945 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4948 = (inp[5]) ? node4968 : node4949;
										assign node4949 = (inp[3]) ? node4957 : node4950;
											assign node4950 = (inp[4]) ? 15'b000000000111111 : node4951;
												assign node4951 = (inp[7]) ? node4953 : 15'b000000001111111;
													assign node4953 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4957 = (inp[7]) ? node4963 : node4958;
												assign node4958 = (inp[4]) ? node4960 : 15'b000000000111111;
													assign node4960 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4963 = (inp[11]) ? 15'b000000000001111 : node4964;
													assign node4964 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4968 = (inp[11]) ? node4974 : node4969;
											assign node4969 = (inp[3]) ? node4971 : 15'b000000011111111;
												assign node4971 = (inp[4]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node4974 = (inp[14]) ? node4976 : 15'b000000000000111;
												assign node4976 = (inp[8]) ? 15'b000000000001111 : node4977;
													assign node4977 = (inp[7]) ? 15'b000000000011111 : 15'b000000000001111;
							assign node4981 = (inp[13]) ? node5023 : node4982;
								assign node4982 = (inp[5]) ? node5006 : node4983;
									assign node4983 = (inp[9]) ? node4999 : node4984;
										assign node4984 = (inp[11]) ? node4990 : node4985;
											assign node4985 = (inp[14]) ? 15'b000000011111111 : node4986;
												assign node4986 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4990 = (inp[3]) ? node4994 : node4991;
												assign node4991 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4994 = (inp[14]) ? node4996 : 15'b000000000111111;
													assign node4996 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4999 = (inp[3]) ? node5003 : node5000;
											assign node5000 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node5003 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5006 = (inp[3]) ? node5014 : node5007;
										assign node5007 = (inp[4]) ? node5011 : node5008;
											assign node5008 = (inp[14]) ? 15'b000000001111111 : 15'b000000000011111;
											assign node5011 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5014 = (inp[9]) ? node5020 : node5015;
											assign node5015 = (inp[8]) ? 15'b000000000011111 : node5016;
												assign node5016 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5020 = (inp[8]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node5023 = (inp[14]) ? node5041 : node5024;
									assign node5024 = (inp[8]) ? node5036 : node5025;
										assign node5025 = (inp[9]) ? node5029 : node5026;
											assign node5026 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5029 = (inp[11]) ? 15'b000000000011111 : node5030;
												assign node5030 = (inp[7]) ? node5032 : 15'b000000001111111;
													assign node5032 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5036 = (inp[11]) ? 15'b000000000011111 : node5037;
											assign node5037 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5041 = (inp[7]) ? node5057 : node5042;
										assign node5042 = (inp[11]) ? node5048 : node5043;
											assign node5043 = (inp[4]) ? node5045 : 15'b000000000111111;
												assign node5045 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node5048 = (inp[9]) ? node5050 : 15'b000000000011111;
												assign node5050 = (inp[5]) ? 15'b000000000001111 : node5051;
													assign node5051 = (inp[8]) ? node5053 : 15'b000000000011111;
														assign node5053 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5057 = (inp[5]) ? node5065 : node5058;
											assign node5058 = (inp[11]) ? node5060 : 15'b000000000011111;
												assign node5060 = (inp[3]) ? 15'b000000000001111 : node5061;
													assign node5061 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5065 = (inp[9]) ? 15'b000000000000111 : node5066;
												assign node5066 = (inp[3]) ? node5068 : 15'b000000000011111;
													assign node5068 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node5072 = (inp[4]) ? node5436 : node5073;
					assign node5073 = (inp[11]) ? node5277 : node5074;
						assign node5074 = (inp[3]) ? node5170 : node5075;
							assign node5075 = (inp[7]) ? node5127 : node5076;
								assign node5076 = (inp[9]) ? node5102 : node5077;
									assign node5077 = (inp[13]) ? node5089 : node5078;
										assign node5078 = (inp[5]) ? 15'b000000111111111 : node5079;
											assign node5079 = (inp[0]) ? node5085 : node5080;
												assign node5080 = (inp[1]) ? 15'b000001111111111 : node5081;
													assign node5081 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5085 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node5089 = (inp[8]) ? node5095 : node5090;
											assign node5090 = (inp[5]) ? 15'b000000011111111 : node5091;
												assign node5091 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5095 = (inp[14]) ? node5097 : 15'b000000011111111;
												assign node5097 = (inp[0]) ? 15'b000000000111111 : node5098;
													assign node5098 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5102 = (inp[13]) ? node5116 : node5103;
										assign node5103 = (inp[14]) ? node5109 : node5104;
											assign node5104 = (inp[1]) ? node5106 : 15'b000001111111111;
												assign node5106 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5109 = (inp[8]) ? 15'b000000001111111 : node5110;
												assign node5110 = (inp[5]) ? 15'b000000011111111 : node5111;
													assign node5111 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5116 = (inp[0]) ? node5120 : node5117;
											assign node5117 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5120 = (inp[6]) ? 15'b000000000111111 : node5121;
												assign node5121 = (inp[5]) ? node5123 : 15'b000000001111111;
													assign node5123 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5127 = (inp[13]) ? node5151 : node5128;
									assign node5128 = (inp[8]) ? node5138 : node5129;
										assign node5129 = (inp[14]) ? node5133 : node5130;
											assign node5130 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node5133 = (inp[5]) ? node5135 : 15'b000000011111111;
												assign node5135 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5138 = (inp[0]) ? node5144 : node5139;
											assign node5139 = (inp[9]) ? 15'b000000001111111 : node5140;
												assign node5140 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node5144 = (inp[9]) ? node5146 : 15'b000000001111111;
												assign node5146 = (inp[6]) ? node5148 : 15'b000000001111111;
													assign node5148 = (inp[14]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node5151 = (inp[0]) ? node5163 : node5152;
										assign node5152 = (inp[1]) ? node5156 : node5153;
											assign node5153 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5156 = (inp[5]) ? 15'b000000000111111 : node5157;
												assign node5157 = (inp[6]) ? node5159 : 15'b000000011111111;
													assign node5159 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5163 = (inp[8]) ? node5167 : node5164;
											assign node5164 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node5167 = (inp[14]) ? 15'b000000000011111 : 15'b000000000001111;
							assign node5170 = (inp[13]) ? node5210 : node5171;
								assign node5171 = (inp[9]) ? node5193 : node5172;
									assign node5172 = (inp[6]) ? node5182 : node5173;
										assign node5173 = (inp[8]) ? node5179 : node5174;
											assign node5174 = (inp[0]) ? 15'b000000111111111 : node5175;
												assign node5175 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5179 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5182 = (inp[7]) ? node5186 : node5183;
											assign node5183 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5186 = (inp[0]) ? 15'b000000000111111 : node5187;
												assign node5187 = (inp[1]) ? node5189 : 15'b000000001111111;
													assign node5189 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5193 = (inp[8]) ? node5195 : 15'b000000001111111;
										assign node5195 = (inp[7]) ? node5205 : node5196;
											assign node5196 = (inp[14]) ? node5202 : node5197;
												assign node5197 = (inp[6]) ? 15'b000000001111111 : node5198;
													assign node5198 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5202 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5205 = (inp[6]) ? 15'b000000000001111 : node5206;
												assign node5206 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5210 = (inp[5]) ? node5244 : node5211;
									assign node5211 = (inp[0]) ? node5227 : node5212;
										assign node5212 = (inp[7]) ? node5220 : node5213;
											assign node5213 = (inp[8]) ? 15'b000000011111111 : node5214;
												assign node5214 = (inp[9]) ? node5216 : 15'b000000111111111;
													assign node5216 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5220 = (inp[8]) ? node5222 : 15'b000000001111111;
												assign node5222 = (inp[14]) ? 15'b000000000111111 : node5223;
													assign node5223 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5227 = (inp[8]) ? node5239 : node5228;
											assign node5228 = (inp[7]) ? node5234 : node5229;
												assign node5229 = (inp[14]) ? 15'b000000001111111 : node5230;
													assign node5230 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5234 = (inp[6]) ? node5236 : 15'b000000001111111;
													assign node5236 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5239 = (inp[6]) ? 15'b000000000011111 : node5240;
												assign node5240 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5244 = (inp[14]) ? node5256 : node5245;
										assign node5245 = (inp[6]) ? node5251 : node5246;
											assign node5246 = (inp[9]) ? node5248 : 15'b000000000011111;
												assign node5248 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5251 = (inp[9]) ? node5253 : 15'b000000000111111;
												assign node5253 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5256 = (inp[6]) ? node5262 : node5257;
											assign node5257 = (inp[1]) ? 15'b000000000001111 : node5258;
												assign node5258 = (inp[0]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node5262 = (inp[0]) ? node5268 : node5263;
												assign node5263 = (inp[1]) ? node5265 : 15'b000000000011111;
													assign node5265 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5268 = (inp[1]) ? 15'b000000000001111 : node5269;
													assign node5269 = (inp[9]) ? 15'b000000000001111 : node5270;
														assign node5270 = (inp[7]) ? node5272 : 15'b000000000011111;
															assign node5272 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node5277 = (inp[5]) ? node5349 : node5278;
							assign node5278 = (inp[1]) ? node5320 : node5279;
								assign node5279 = (inp[0]) ? node5295 : node5280;
									assign node5280 = (inp[8]) ? node5288 : node5281;
										assign node5281 = (inp[3]) ? node5283 : 15'b000001111111111;
											assign node5283 = (inp[6]) ? 15'b000000011111111 : node5284;
												assign node5284 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5288 = (inp[6]) ? node5292 : node5289;
											assign node5289 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node5292 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node5295 = (inp[7]) ? node5307 : node5296;
										assign node5296 = (inp[14]) ? node5304 : node5297;
											assign node5297 = (inp[3]) ? node5301 : node5298;
												assign node5298 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5301 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5304 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5307 = (inp[9]) ? node5311 : node5308;
											assign node5308 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5311 = (inp[3]) ? node5315 : node5312;
												assign node5312 = (inp[14]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node5315 = (inp[6]) ? node5317 : 15'b000000000011111;
													assign node5317 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node5320 = (inp[9]) ? node5338 : node5321;
									assign node5321 = (inp[8]) ? node5323 : 15'b000000111111111;
										assign node5323 = (inp[0]) ? node5335 : node5324;
											assign node5324 = (inp[14]) ? 15'b000000000011111 : node5325;
												assign node5325 = (inp[6]) ? node5329 : node5326;
													assign node5326 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node5329 = (inp[7]) ? node5331 : 15'b000000001111111;
														assign node5331 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5335 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5338 = (inp[13]) ? node5344 : node5339;
										assign node5339 = (inp[3]) ? 15'b000000000011111 : node5340;
											assign node5340 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5344 = (inp[3]) ? node5346 : 15'b000000000001111;
											assign node5346 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
							assign node5349 = (inp[7]) ? node5397 : node5350;
								assign node5350 = (inp[8]) ? node5376 : node5351;
									assign node5351 = (inp[0]) ? node5363 : node5352;
										assign node5352 = (inp[1]) ? node5356 : node5353;
											assign node5353 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5356 = (inp[9]) ? node5358 : 15'b000000001111111;
												assign node5358 = (inp[3]) ? 15'b000000000111111 : node5359;
													assign node5359 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5363 = (inp[6]) ? node5369 : node5364;
											assign node5364 = (inp[14]) ? 15'b000000000111111 : node5365;
												assign node5365 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5369 = (inp[1]) ? node5371 : 15'b000000000111111;
												assign node5371 = (inp[9]) ? node5373 : 15'b000000000111111;
													assign node5373 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5376 = (inp[14]) ? node5392 : node5377;
										assign node5377 = (inp[6]) ? node5381 : node5378;
											assign node5378 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5381 = (inp[3]) ? node5387 : node5382;
												assign node5382 = (inp[13]) ? node5384 : 15'b000000001111111;
													assign node5384 = (inp[0]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node5387 = (inp[13]) ? node5389 : 15'b000000000011111;
													assign node5389 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5392 = (inp[9]) ? node5394 : 15'b000000000011111;
											assign node5394 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node5397 = (inp[3]) ? node5417 : node5398;
									assign node5398 = (inp[14]) ? node5410 : node5399;
										assign node5399 = (inp[9]) ? node5405 : node5400;
											assign node5400 = (inp[0]) ? 15'b000000000111111 : node5401;
												assign node5401 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5405 = (inp[1]) ? node5407 : 15'b000000001111111;
												assign node5407 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5410 = (inp[1]) ? node5414 : node5411;
											assign node5411 = (inp[0]) ? 15'b000000000011111 : 15'b000000011111111;
											assign node5414 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5417 = (inp[0]) ? node5425 : node5418;
										assign node5418 = (inp[9]) ? node5420 : 15'b000000000011111;
											assign node5420 = (inp[8]) ? node5422 : 15'b000000000011111;
												assign node5422 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5425 = (inp[8]) ? node5429 : node5426;
											assign node5426 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5429 = (inp[9]) ? 15'b000000000000111 : node5430;
												assign node5430 = (inp[6]) ? node5432 : 15'b000000000001111;
													assign node5432 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node5436 = (inp[8]) ? node5618 : node5437;
						assign node5437 = (inp[3]) ? node5525 : node5438;
							assign node5438 = (inp[0]) ? node5476 : node5439;
								assign node5439 = (inp[5]) ? node5461 : node5440;
									assign node5440 = (inp[11]) ? node5448 : node5441;
										assign node5441 = (inp[6]) ? 15'b000000011111111 : node5442;
											assign node5442 = (inp[14]) ? node5444 : 15'b000000111111111;
												assign node5444 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5448 = (inp[6]) ? node5456 : node5449;
											assign node5449 = (inp[1]) ? 15'b000000001111111 : node5450;
												assign node5450 = (inp[7]) ? node5452 : 15'b000000111111111;
													assign node5452 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5456 = (inp[14]) ? node5458 : 15'b000000001111111;
												assign node5458 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5461 = (inp[7]) ? node5471 : node5462;
										assign node5462 = (inp[1]) ? node5466 : node5463;
											assign node5463 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5466 = (inp[9]) ? node5468 : 15'b000000001111111;
												assign node5468 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5471 = (inp[11]) ? node5473 : 15'b000000000111111;
											assign node5473 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5476 = (inp[6]) ? node5488 : node5477;
									assign node5477 = (inp[13]) ? node5483 : node5478;
										assign node5478 = (inp[9]) ? node5480 : 15'b000000011111111;
											assign node5480 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5483 = (inp[1]) ? node5485 : 15'b000000000111111;
											assign node5485 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5488 = (inp[14]) ? node5510 : node5489;
										assign node5489 = (inp[7]) ? node5497 : node5490;
											assign node5490 = (inp[9]) ? node5494 : node5491;
												assign node5491 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5494 = (inp[13]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node5497 = (inp[13]) ? node5503 : node5498;
												assign node5498 = (inp[11]) ? node5500 : 15'b000000000111111;
													assign node5500 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5503 = (inp[5]) ? 15'b000000000001111 : node5504;
													assign node5504 = (inp[11]) ? 15'b000000000011111 : node5505;
														assign node5505 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5510 = (inp[11]) ? node5520 : node5511;
											assign node5511 = (inp[13]) ? 15'b000000000001111 : node5512;
												assign node5512 = (inp[1]) ? node5514 : 15'b000000001111111;
													assign node5514 = (inp[9]) ? node5516 : 15'b000000000111111;
														assign node5516 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5520 = (inp[5]) ? 15'b000000000001111 : node5521;
												assign node5521 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node5525 = (inp[1]) ? node5569 : node5526;
								assign node5526 = (inp[9]) ? node5548 : node5527;
									assign node5527 = (inp[0]) ? node5543 : node5528;
										assign node5528 = (inp[11]) ? node5530 : 15'b000000001111111;
											assign node5530 = (inp[6]) ? node5536 : node5531;
												assign node5531 = (inp[13]) ? node5533 : 15'b000000011111111;
													assign node5533 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node5536 = (inp[5]) ? 15'b000000000111111 : node5537;
													assign node5537 = (inp[13]) ? 15'b000000000111111 : node5538;
														assign node5538 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5543 = (inp[7]) ? 15'b000000000011111 : node5544;
											assign node5544 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5548 = (inp[13]) ? node5558 : node5549;
										assign node5549 = (inp[14]) ? node5553 : node5550;
											assign node5550 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5553 = (inp[7]) ? node5555 : 15'b000000000111111;
												assign node5555 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5558 = (inp[0]) ? node5562 : node5559;
											assign node5559 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5562 = (inp[6]) ? 15'b000000000001111 : node5563;
												assign node5563 = (inp[5]) ? 15'b000000000001111 : node5564;
													assign node5564 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5569 = (inp[9]) ? node5593 : node5570;
									assign node5570 = (inp[6]) ? node5582 : node5571;
										assign node5571 = (inp[7]) ? node5575 : node5572;
											assign node5572 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5575 = (inp[14]) ? node5577 : 15'b000000000111111;
												assign node5577 = (inp[13]) ? 15'b000000000011111 : node5578;
													assign node5578 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5582 = (inp[13]) ? node5586 : node5583;
											assign node5583 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node5586 = (inp[5]) ? 15'b000000000001111 : node5587;
												assign node5587 = (inp[11]) ? 15'b000000000001111 : node5588;
													assign node5588 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5593 = (inp[7]) ? node5611 : node5594;
										assign node5594 = (inp[6]) ? node5602 : node5595;
											assign node5595 = (inp[14]) ? node5597 : 15'b000000000011111;
												assign node5597 = (inp[0]) ? node5599 : 15'b000000000011111;
													assign node5599 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5602 = (inp[0]) ? node5608 : node5603;
												assign node5603 = (inp[11]) ? node5605 : 15'b000000000011111;
													assign node5605 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5608 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node5611 = (inp[14]) ? node5613 : 15'b000000000001111;
											assign node5613 = (inp[13]) ? node5615 : 15'b000000000001111;
												assign node5615 = (inp[0]) ? 15'b000000000000011 : 15'b000000000000111;
						assign node5618 = (inp[14]) ? node5728 : node5619;
							assign node5619 = (inp[0]) ? node5665 : node5620;
								assign node5620 = (inp[9]) ? node5646 : node5621;
									assign node5621 = (inp[3]) ? node5635 : node5622;
										assign node5622 = (inp[13]) ? node5632 : node5623;
											assign node5623 = (inp[7]) ? node5625 : 15'b000000011111111;
												assign node5625 = (inp[5]) ? 15'b000000000111111 : node5626;
													assign node5626 = (inp[11]) ? 15'b000000001111111 : node5627;
														assign node5627 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5632 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5635 = (inp[1]) ? node5639 : node5636;
											assign node5636 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5639 = (inp[11]) ? 15'b000000000011111 : node5640;
												assign node5640 = (inp[13]) ? node5642 : 15'b000000001111111;
													assign node5642 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5646 = (inp[7]) ? node5652 : node5647;
										assign node5647 = (inp[13]) ? node5649 : 15'b000000000111111;
											assign node5649 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5652 = (inp[11]) ? node5658 : node5653;
											assign node5653 = (inp[5]) ? node5655 : 15'b000000000111111;
												assign node5655 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5658 = (inp[13]) ? node5662 : node5659;
												assign node5659 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5662 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node5665 = (inp[6]) ? node5703 : node5666;
									assign node5666 = (inp[1]) ? node5684 : node5667;
										assign node5667 = (inp[7]) ? node5677 : node5668;
											assign node5668 = (inp[9]) ? 15'b000000000011111 : node5669;
												assign node5669 = (inp[3]) ? 15'b000000000111111 : node5670;
													assign node5670 = (inp[13]) ? node5672 : 15'b000000001111111;
														assign node5672 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5677 = (inp[5]) ? node5679 : 15'b000000000111111;
												assign node5679 = (inp[3]) ? 15'b000000000011111 : node5680;
													assign node5680 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5684 = (inp[13]) ? node5696 : node5685;
											assign node5685 = (inp[9]) ? node5687 : 15'b000000000001111;
												assign node5687 = (inp[5]) ? node5689 : 15'b000000000111111;
													assign node5689 = (inp[11]) ? 15'b000000000011111 : node5690;
														assign node5690 = (inp[7]) ? 15'b000000000011111 : node5691;
															assign node5691 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5696 = (inp[7]) ? node5698 : 15'b000000000011111;
												assign node5698 = (inp[11]) ? node5700 : 15'b000000000001111;
													assign node5700 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node5703 = (inp[7]) ? node5719 : node5704;
										assign node5704 = (inp[11]) ? node5712 : node5705;
											assign node5705 = (inp[13]) ? 15'b000000000011111 : node5706;
												assign node5706 = (inp[1]) ? node5708 : 15'b000000000111111;
													assign node5708 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5712 = (inp[9]) ? 15'b000000000001111 : node5713;
												assign node5713 = (inp[1]) ? node5715 : 15'b000000000011111;
													assign node5715 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5719 = (inp[11]) ? node5725 : node5720;
											assign node5720 = (inp[3]) ? 15'b000000000001111 : node5721;
												assign node5721 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5725 = (inp[13]) ? 15'b000000000000001 : 15'b000000000001111;
							assign node5728 = (inp[1]) ? node5778 : node5729;
								assign node5729 = (inp[5]) ? node5749 : node5730;
									assign node5730 = (inp[11]) ? node5736 : node5731;
										assign node5731 = (inp[13]) ? node5733 : 15'b000000000111111;
											assign node5733 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node5736 = (inp[7]) ? node5744 : node5737;
											assign node5737 = (inp[6]) ? 15'b000000000011111 : node5738;
												assign node5738 = (inp[0]) ? node5740 : 15'b000000000111111;
													assign node5740 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5744 = (inp[13]) ? node5746 : 15'b000000000011111;
												assign node5746 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5749 = (inp[0]) ? node5769 : node5750;
										assign node5750 = (inp[3]) ? node5754 : node5751;
											assign node5751 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5754 = (inp[11]) ? node5764 : node5755;
												assign node5755 = (inp[9]) ? node5761 : node5756;
													assign node5756 = (inp[7]) ? 15'b000000000011111 : node5757;
														assign node5757 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5761 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5764 = (inp[9]) ? node5766 : 15'b000000000001111;
													assign node5766 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node5769 = (inp[9]) ? 15'b000000000000111 : node5770;
											assign node5770 = (inp[13]) ? node5772 : 15'b000000000011111;
												assign node5772 = (inp[3]) ? node5774 : 15'b000000000001111;
													assign node5774 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node5778 = (inp[7]) ? node5802 : node5779;
									assign node5779 = (inp[11]) ? node5789 : node5780;
										assign node5780 = (inp[5]) ? node5784 : node5781;
											assign node5781 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5784 = (inp[9]) ? node5786 : 15'b000000000011111;
												assign node5786 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5789 = (inp[0]) ? node5795 : node5790;
											assign node5790 = (inp[9]) ? node5792 : 15'b000000000001111;
												assign node5792 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5795 = (inp[5]) ? 15'b000000000000111 : node5796;
												assign node5796 = (inp[6]) ? node5798 : 15'b000000000001111;
													assign node5798 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node5802 = (inp[5]) ? node5814 : node5803;
										assign node5803 = (inp[11]) ? node5809 : node5804;
											assign node5804 = (inp[13]) ? node5806 : 15'b000000000001111;
												assign node5806 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5809 = (inp[6]) ? 15'b000000000000011 : node5810;
												assign node5810 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node5814 = (inp[0]) ? node5820 : node5815;
											assign node5815 = (inp[9]) ? 15'b000000000000111 : node5816;
												assign node5816 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node5820 = (inp[13]) ? node5822 : 15'b000000000000111;
												assign node5822 = (inp[3]) ? 15'b000000000000000 : node5823;
													assign node5823 = (inp[9]) ? node5825 : 15'b000000000000011;
														assign node5825 = (inp[11]) ? 15'b000000000000001 : 15'b000000000000011;

endmodule