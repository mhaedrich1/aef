module dtc_split5_bm12 (
	input  wire [9-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node12;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node17;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node31;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node35;
	wire [1-1:0] node37;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node51;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node67;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node77;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node85;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node92;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node97;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node122;
	wire [1-1:0] node123;
	wire [1-1:0] node124;
	wire [1-1:0] node125;

	assign outp = (inp[1]) ? node60 : node1;
		assign node1 = (inp[4]) ? node31 : node2;
			assign node2 = (inp[3]) ? node12 : node3;
				assign node3 = (inp[7]) ? node5 : 1'b1;
					assign node5 = (inp[5]) ? node7 : 1'b1;
						assign node7 = (inp[8]) ? node9 : 1'b1;
							assign node9 = (inp[6]) ? 1'b0 : 1'b1;
				assign node12 = (inp[7]) ? node20 : node13;
					assign node13 = (inp[6]) ? node15 : 1'b1;
						assign node15 = (inp[5]) ? node17 : 1'b1;
							assign node17 = (inp[0]) ? 1'b0 : 1'b1;
					assign node20 = (inp[6]) ? node26 : node21;
						assign node21 = (inp[0]) ? node23 : 1'b1;
							assign node23 = (inp[8]) ? 1'b0 : 1'b1;
						assign node26 = (inp[5]) ? 1'b0 : node27;
							assign node27 = (inp[8]) ? 1'b0 : 1'b1;
			assign node31 = (inp[0]) ? node51 : node32;
				assign node32 = (inp[3]) ? node40 : node33;
					assign node33 = (inp[7]) ? node35 : 1'b1;
						assign node35 = (inp[6]) ? node37 : 1'b1;
							assign node37 = (inp[2]) ? 1'b0 : 1'b1;
					assign node40 = (inp[6]) ? node46 : node41;
						assign node41 = (inp[5]) ? node43 : 1'b1;
							assign node43 = (inp[8]) ? 1'b0 : 1'b1;
						assign node46 = (inp[7]) ? 1'b0 : node47;
							assign node47 = (inp[5]) ? 1'b0 : 1'b1;
				assign node51 = (inp[3]) ? 1'b0 : node52;
					assign node52 = (inp[2]) ? node54 : 1'b1;
						assign node54 = (inp[6]) ? 1'b0 : node55;
							assign node55 = (inp[7]) ? 1'b0 : 1'b1;
		assign node60 = (inp[8]) ? node102 : node61;
			assign node61 = (inp[0]) ? node81 : node62;
				assign node62 = (inp[6]) ? node70 : node63;
					assign node63 = (inp[4]) ? node65 : 1'b1;
						assign node65 = (inp[7]) ? node67 : 1'b1;
							assign node67 = (inp[3]) ? 1'b0 : 1'b1;
					assign node70 = (inp[3]) ? node76 : node71;
						assign node71 = (inp[2]) ? node73 : 1'b1;
							assign node73 = (inp[5]) ? 1'b0 : 1'b1;
						assign node76 = (inp[7]) ? 1'b0 : node77;
							assign node77 = (inp[5]) ? 1'b0 : 1'b1;
				assign node81 = (inp[7]) ? node95 : node82;
					assign node82 = (inp[2]) ? node88 : node83;
						assign node83 = (inp[5]) ? node85 : 1'b1;
							assign node85 = (inp[6]) ? 1'b0 : 1'b1;
						assign node88 = (inp[4]) ? node92 : node89;
							assign node89 = (inp[5]) ? 1'b0 : 1'b1;
							assign node92 = (inp[3]) ? 1'b0 : 1'b0;
					assign node95 = (inp[3]) ? 1'b0 : node96;
						assign node96 = (inp[5]) ? 1'b0 : node97;
							assign node97 = (inp[2]) ? 1'b0 : 1'b0;
			assign node102 = (inp[5]) ? node122 : node103;
				assign node103 = (inp[2]) ? node115 : node104;
					assign node104 = (inp[7]) ? node110 : node105;
						assign node105 = (inp[4]) ? node107 : 1'b1;
							assign node107 = (inp[6]) ? 1'b0 : 1'b1;
						assign node110 = (inp[0]) ? 1'b0 : node111;
							assign node111 = (inp[6]) ? 1'b0 : 1'b1;
					assign node115 = (inp[0]) ? 1'b0 : node116;
						assign node116 = (inp[4]) ? 1'b0 : node117;
							assign node117 = (inp[6]) ? 1'b0 : 1'b1;
				assign node122 = (inp[0]) ? 1'b0 : node123;
					assign node123 = (inp[3]) ? 1'b0 : node124;
						assign node124 = (inp[6]) ? 1'b0 : node125;
							assign node125 = (inp[2]) ? 1'b0 : 1'b1;

endmodule