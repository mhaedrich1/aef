module dtc_split125_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node28;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node35;
	wire [1-1:0] node38;
	wire [1-1:0] node39;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node77;
	wire [1-1:0] node79;
	wire [1-1:0] node81;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node97;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node107;
	wire [1-1:0] node108;
	wire [1-1:0] node110;
	wire [1-1:0] node112;
	wire [1-1:0] node115;
	wire [1-1:0] node117;
	wire [1-1:0] node120;
	wire [1-1:0] node121;
	wire [1-1:0] node123;
	wire [1-1:0] node124;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node135;
	wire [1-1:0] node137;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node151;
	wire [1-1:0] node154;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node171;
	wire [1-1:0] node173;
	wire [1-1:0] node175;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node181;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node191;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node204;
	wire [1-1:0] node205;
	wire [1-1:0] node209;
	wire [1-1:0] node210;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node215;
	wire [1-1:0] node217;
	wire [1-1:0] node220;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node233;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node237;
	wire [1-1:0] node239;
	wire [1-1:0] node242;
	wire [1-1:0] node243;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node263;
	wire [1-1:0] node265;
	wire [1-1:0] node267;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node273;
	wire [1-1:0] node276;
	wire [1-1:0] node277;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node289;
	wire [1-1:0] node292;
	wire [1-1:0] node293;
	wire [1-1:0] node295;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node311;
	wire [1-1:0] node313;
	wire [1-1:0] node315;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node325;
	wire [1-1:0] node327;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node337;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node347;
	wire [1-1:0] node349;
	wire [1-1:0] node352;
	wire [1-1:0] node353;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node364;
	wire [1-1:0] node365;
	wire [1-1:0] node366;
	wire [1-1:0] node368;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node373;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node385;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node396;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node401;
	wire [1-1:0] node403;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node421;
	wire [1-1:0] node423;
	wire [1-1:0] node425;
	wire [1-1:0] node428;
	wire [1-1:0] node429;
	wire [1-1:0] node431;
	wire [1-1:0] node433;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node442;
	wire [1-1:0] node446;
	wire [1-1:0] node447;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node454;
	wire [1-1:0] node455;
	wire [1-1:0] node457;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node487;
	wire [1-1:0] node488;
	wire [1-1:0] node489;
	wire [1-1:0] node491;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node497;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node504;
	wire [1-1:0] node505;
	wire [1-1:0] node507;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node512;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node525;
	wire [1-1:0] node527;
	wire [1-1:0] node528;
	wire [1-1:0] node530;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node549;
	wire [1-1:0] node551;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node557;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node565;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node569;
	wire [1-1:0] node572;
	wire [1-1:0] node573;
	wire [1-1:0] node578;
	wire [1-1:0] node579;
	wire [1-1:0] node580;
	wire [1-1:0] node581;
	wire [1-1:0] node583;
	wire [1-1:0] node585;
	wire [1-1:0] node588;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node611;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node618;
	wire [1-1:0] node619;
	wire [1-1:0] node620;
	wire [1-1:0] node621;
	wire [1-1:0] node623;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node630;
	wire [1-1:0] node631;
	wire [1-1:0] node632;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node640;
	wire [1-1:0] node642;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node657;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node661;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node667;
	wire [1-1:0] node670;
	wire [1-1:0] node671;
	wire [1-1:0] node673;
	wire [1-1:0] node674;
	wire [1-1:0] node676;
	wire [1-1:0] node680;
	wire [1-1:0] node681;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node693;
	wire [1-1:0] node694;
	wire [1-1:0] node695;
	wire [1-1:0] node697;
	wire [1-1:0] node699;
	wire [1-1:0] node702;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node713;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node718;
	wire [1-1:0] node723;
	wire [1-1:0] node724;
	wire [1-1:0] node728;
	wire [1-1:0] node729;
	wire [1-1:0] node730;
	wire [1-1:0] node731;
	wire [1-1:0] node733;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node743;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node753;
	wire [1-1:0] node754;
	wire [1-1:0] node755;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node763;
	wire [1-1:0] node765;
	wire [1-1:0] node767;
	wire [1-1:0] node769;
	wire [1-1:0] node772;
	wire [1-1:0] node773;
	wire [1-1:0] node774;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node783;
	wire [1-1:0] node784;
	wire [1-1:0] node785;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node792;
	wire [1-1:0] node793;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node807;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node819;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node825;
	wire [1-1:0] node828;
	wire [1-1:0] node829;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node843;
	wire [1-1:0] node844;
	wire [1-1:0] node846;
	wire [1-1:0] node850;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node854;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node864;
	wire [1-1:0] node866;
	wire [1-1:0] node867;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node877;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node898;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node902;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node915;
	wire [1-1:0] node916;
	wire [1-1:0] node924;
	wire [1-1:0] node925;
	wire [1-1:0] node926;
	wire [1-1:0] node927;
	wire [1-1:0] node928;
	wire [1-1:0] node930;
	wire [1-1:0] node932;
	wire [1-1:0] node933;
	wire [1-1:0] node935;
	wire [1-1:0] node938;
	wire [1-1:0] node939;
	wire [1-1:0] node941;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node948;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node952;
	wire [1-1:0] node957;
	wire [1-1:0] node958;
	wire [1-1:0] node959;
	wire [1-1:0] node961;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node966;
	wire [1-1:0] node968;
	wire [1-1:0] node972;
	wire [1-1:0] node973;
	wire [1-1:0] node975;
	wire [1-1:0] node977;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node983;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node993;
	wire [1-1:0] node996;
	wire [1-1:0] node998;
	wire [1-1:0] node999;
	wire [1-1:0] node1001;
	wire [1-1:0] node1002;
	wire [1-1:0] node1007;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1014;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1021;
	wire [1-1:0] node1022;
	wire [1-1:0] node1023;
	wire [1-1:0] node1030;
	wire [1-1:0] node1031;
	wire [1-1:0] node1032;
	wire [1-1:0] node1034;
	wire [1-1:0] node1035;
	wire [1-1:0] node1037;
	wire [1-1:0] node1038;
	wire [1-1:0] node1040;
	wire [1-1:0] node1042;
	wire [1-1:0] node1046;
	wire [1-1:0] node1047;
	wire [1-1:0] node1049;
	wire [1-1:0] node1051;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1059;
	wire [1-1:0] node1060;
	wire [1-1:0] node1061;
	wire [1-1:0] node1063;
	wire [1-1:0] node1065;
	wire [1-1:0] node1066;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1073;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1081;
	wire [1-1:0] node1082;
	wire [1-1:0] node1083;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1092;
	wire [1-1:0] node1093;
	wire [1-1:0] node1094;
	wire [1-1:0] node1095;
	wire [1-1:0] node1097;
	wire [1-1:0] node1099;
	wire [1-1:0] node1102;
	wire [1-1:0] node1104;
	wire [1-1:0] node1105;
	wire [1-1:0] node1107;
	wire [1-1:0] node1111;
	wire [1-1:0] node1112;
	wire [1-1:0] node1113;
	wire [1-1:0] node1115;
	wire [1-1:0] node1119;
	wire [1-1:0] node1120;
	wire [1-1:0] node1121;
	wire [1-1:0] node1123;
	wire [1-1:0] node1128;
	wire [1-1:0] node1129;
	wire [1-1:0] node1130;
	wire [1-1:0] node1131;
	wire [1-1:0] node1133;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1139;
	wire [1-1:0] node1143;
	wire [1-1:0] node1144;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1150;
	wire [1-1:0] node1151;
	wire [1-1:0] node1157;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1160;
	wire [1-1:0] node1161;
	wire [1-1:0] node1163;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1168;
	wire [1-1:0] node1172;
	wire [1-1:0] node1173;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1177;
	wire [1-1:0] node1179;
	wire [1-1:0] node1183;
	wire [1-1:0] node1186;
	wire [1-1:0] node1189;
	wire [1-1:0] node1190;
	wire [1-1:0] node1191;
	wire [1-1:0] node1193;
	wire [1-1:0] node1195;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1201;
	wire [1-1:0] node1204;
	wire [1-1:0] node1206;
	wire [1-1:0] node1209;
	wire [1-1:0] node1210;
	wire [1-1:0] node1211;
	wire [1-1:0] node1213;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1222;
	wire [1-1:0] node1223;
	wire [1-1:0] node1224;
	wire [1-1:0] node1225;
	wire [1-1:0] node1227;
	wire [1-1:0] node1229;
	wire [1-1:0] node1232;
	wire [1-1:0] node1233;
	wire [1-1:0] node1235;
	wire [1-1:0] node1239;
	wire [1-1:0] node1240;
	wire [1-1:0] node1241;
	wire [1-1:0] node1243;
	wire [1-1:0] node1246;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1265;
	wire [1-1:0] node1266;
	wire [1-1:0] node1268;
	wire [1-1:0] node1272;
	wire [1-1:0] node1273;
	wire [1-1:0] node1274;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1281;
	wire [1-1:0] node1282;
	wire [1-1:0] node1283;
	wire [1-1:0] node1285;
	wire [1-1:0] node1287;
	wire [1-1:0] node1290;
	wire [1-1:0] node1291;
	wire [1-1:0] node1293;
	wire [1-1:0] node1294;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1303;
	wire [1-1:0] node1304;
	wire [1-1:0] node1305;
	wire [1-1:0] node1307;
	wire [1-1:0] node1310;
	wire [1-1:0] node1314;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1319;
	wire [1-1:0] node1320;
	wire [1-1:0] node1324;
	wire [1-1:0] node1325;
	wire [1-1:0] node1329;
	wire [1-1:0] node1330;
	wire [1-1:0] node1331;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1347;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1351;
	wire [1-1:0] node1354;
	wire [1-1:0] node1355;
	wire [1-1:0] node1359;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1370;
	wire [1-1:0] node1372;
	wire [1-1:0] node1376;
	wire [1-1:0] node1377;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1385;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1396;
	wire [1-1:0] node1397;
	wire [1-1:0] node1398;
	wire [1-1:0] node1399;
	wire [1-1:0] node1401;
	wire [1-1:0] node1403;
	wire [1-1:0] node1406;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1411;
	wire [1-1:0] node1412;
	wire [1-1:0] node1414;
	wire [1-1:0] node1417;
	wire [1-1:0] node1418;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1431;
	wire [1-1:0] node1434;
	wire [1-1:0] node1435;
	wire [1-1:0] node1437;
	wire [1-1:0] node1440;
	wire [1-1:0] node1441;
	wire [1-1:0] node1445;
	wire [1-1:0] node1446;
	wire [1-1:0] node1447;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1456;
	wire [1-1:0] node1457;
	wire [1-1:0] node1458;
	wire [1-1:0] node1460;
	wire [1-1:0] node1461;
	wire [1-1:0] node1463;
	wire [1-1:0] node1466;
	wire [1-1:0] node1469;
	wire [1-1:0] node1470;
	wire [1-1:0] node1471;
	wire [1-1:0] node1473;
	wire [1-1:0] node1476;
	wire [1-1:0] node1477;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1487;
	wire [1-1:0] node1489;
	wire [1-1:0] node1492;
	wire [1-1:0] node1493;
	wire [1-1:0] node1495;
	wire [1-1:0] node1496;
	wire [1-1:0] node1501;
	wire [1-1:0] node1502;
	wire [1-1:0] node1504;
	wire [1-1:0] node1505;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1512;
	wire [1-1:0] node1514;
	wire [1-1:0] node1515;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1526;
	wire [1-1:0] node1528;
	wire [1-1:0] node1529;
	wire [1-1:0] node1531;
	wire [1-1:0] node1532;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1541;
	wire [1-1:0] node1544;
	wire [1-1:0] node1545;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1555;
	wire [1-1:0] node1558;
	wire [1-1:0] node1560;
	wire [1-1:0] node1561;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1572;
	wire [1-1:0] node1573;
	wire [1-1:0] node1574;
	wire [1-1:0] node1579;
	wire [1-1:0] node1580;
	wire [1-1:0] node1581;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1585;
	wire [1-1:0] node1588;
	wire [1-1:0] node1589;
	wire [1-1:0] node1593;
	wire [1-1:0] node1594;
	wire [1-1:0] node1595;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1603;
	wire [1-1:0] node1610;
	wire [1-1:0] node1611;
	wire [1-1:0] node1612;
	wire [1-1:0] node1613;
	wire [1-1:0] node1614;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1619;
	wire [1-1:0] node1620;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1627;
	wire [1-1:0] node1629;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1635;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1641;
	wire [1-1:0] node1643;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1650;
	wire [1-1:0] node1652;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1660;
	wire [1-1:0] node1661;
	wire [1-1:0] node1662;
	wire [1-1:0] node1663;
	wire [1-1:0] node1665;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1673;
	wire [1-1:0] node1674;
	wire [1-1:0] node1675;
	wire [1-1:0] node1677;
	wire [1-1:0] node1680;
	wire [1-1:0] node1681;
	wire [1-1:0] node1683;
	wire [1-1:0] node1688;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1693;
	wire [1-1:0] node1699;
	wire [1-1:0] node1700;
	wire [1-1:0] node1701;
	wire [1-1:0] node1702;
	wire [1-1:0] node1708;
	wire [1-1:0] node1709;
	wire [1-1:0] node1710;
	wire [1-1:0] node1711;
	wire [1-1:0] node1712;
	wire [1-1:0] node1713;
	wire [1-1:0] node1715;
	wire [1-1:0] node1716;
	wire [1-1:0] node1720;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1725;
	wire [1-1:0] node1728;
	wire [1-1:0] node1730;
	wire [1-1:0] node1734;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1737;
	wire [1-1:0] node1739;
	wire [1-1:0] node1742;
	wire [1-1:0] node1743;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1753;
	wire [1-1:0] node1760;
	wire [1-1:0] node1761;
	wire [1-1:0] node1762;
	wire [1-1:0] node1763;
	wire [1-1:0] node1764;

	assign outp = (inp[4]) ? node924 : node1;
		assign node1 = (inp[2]) ? node391 : node2;
			assign node2 = (inp[10]) ? node166 : node3;
				assign node3 = (inp[1]) ? node47 : node4;
					assign node4 = (inp[8]) ? node6 : 1'b1;
						assign node6 = (inp[12]) ? node18 : node7;
							assign node7 = (inp[13]) ? node9 : 1'b1;
								assign node9 = (inp[3]) ? node11 : 1'b1;
									assign node11 = (inp[6]) ? node13 : 1'b1;
										assign node13 = (inp[9]) ? node15 : 1'b1;
											assign node15 = (inp[7]) ? 1'b1 : 1'b0;
							assign node18 = (inp[9]) ? node32 : node19;
								assign node19 = (inp[5]) ? node21 : 1'b1;
									assign node21 = (inp[14]) ? node23 : 1'b1;
										assign node23 = (inp[3]) ? node25 : 1'b1;
											assign node25 = (inp[11]) ? 1'b0 : node26;
												assign node26 = (inp[13]) ? node28 : 1'b1;
													assign node28 = (inp[7]) ? 1'b0 : 1'b1;
								assign node32 = (inp[5]) ? node38 : node33;
									assign node33 = (inp[13]) ? node35 : 1'b1;
										assign node35 = (inp[6]) ? 1'b0 : 1'b1;
									assign node38 = (inp[0]) ? 1'b0 : node39;
										assign node39 = (inp[3]) ? node41 : 1'b1;
											assign node41 = (inp[11]) ? 1'b0 : node42;
												assign node42 = (inp[14]) ? 1'b0 : 1'b1;
					assign node47 = (inp[9]) ? node93 : node48;
						assign node48 = (inp[3]) ? node68 : node49;
							assign node49 = (inp[14]) ? node51 : 1'b1;
								assign node51 = (inp[11]) ? node53 : 1'b1;
									assign node53 = (inp[12]) ? node55 : 1'b1;
										assign node55 = (inp[0]) ? node63 : node56;
											assign node56 = (inp[8]) ? node58 : 1'b1;
												assign node58 = (inp[5]) ? node60 : 1'b1;
													assign node60 = (inp[13]) ? 1'b0 : 1'b1;
											assign node63 = (inp[5]) ? 1'b0 : node64;
												assign node64 = (inp[7]) ? 1'b0 : 1'b1;
							assign node68 = (inp[13]) ? node76 : node69;
								assign node69 = (inp[0]) ? node71 : 1'b1;
									assign node71 = (inp[6]) ? node73 : 1'b1;
										assign node73 = (inp[11]) ? 1'b0 : 1'b1;
								assign node76 = (inp[7]) ? node84 : node77;
									assign node77 = (inp[5]) ? node79 : 1'b1;
										assign node79 = (inp[8]) ? node81 : 1'b1;
											assign node81 = (inp[6]) ? 1'b1 : 1'b0;
									assign node84 = (inp[6]) ? node88 : node85;
										assign node85 = (inp[14]) ? 1'b0 : 1'b1;
										assign node88 = (inp[8]) ? 1'b0 : node89;
											assign node89 = (inp[0]) ? 1'b0 : 1'b1;
						assign node93 = (inp[14]) ? node133 : node94;
							assign node94 = (inp[13]) ? node104 : node95;
								assign node95 = (inp[3]) ? node97 : 1'b1;
									assign node97 = (inp[0]) ? node99 : 1'b1;
										assign node99 = (inp[11]) ? node101 : 1'b1;
											assign node101 = (inp[7]) ? 1'b0 : 1'b1;
								assign node104 = (inp[0]) ? node120 : node105;
									assign node105 = (inp[6]) ? node107 : 1'b1;
										assign node107 = (inp[3]) ? node115 : node108;
											assign node108 = (inp[8]) ? node110 : 1'b1;
												assign node110 = (inp[11]) ? node112 : 1'b1;
													assign node112 = (inp[5]) ? 1'b0 : 1'b1;
											assign node115 = (inp[5]) ? node117 : 1'b0;
												assign node117 = (inp[8]) ? 1'b0 : 1'b1;
									assign node120 = (inp[5]) ? node128 : node121;
										assign node121 = (inp[3]) ? node123 : 1'b1;
											assign node123 = (inp[11]) ? 1'b0 : node124;
												assign node124 = (inp[6]) ? 1'b0 : 1'b1;
										assign node128 = (inp[6]) ? 1'b0 : node129;
											assign node129 = (inp[3]) ? 1'b0 : 1'b1;
							assign node133 = (inp[5]) ? node149 : node134;
								assign node134 = (inp[0]) ? node144 : node135;
									assign node135 = (inp[3]) ? node137 : 1'b1;
										assign node137 = (inp[13]) ? node139 : 1'b1;
											assign node139 = (inp[6]) ? 1'b0 : node140;
												assign node140 = (inp[7]) ? 1'b1 : 1'b0;
									assign node144 = (inp[11]) ? 1'b0 : node145;
										assign node145 = (inp[6]) ? 1'b0 : 1'b1;
								assign node149 = (inp[12]) ? node161 : node150;
									assign node150 = (inp[0]) ? node154 : node151;
										assign node151 = (inp[6]) ? 1'b0 : 1'b1;
										assign node154 = (inp[8]) ? 1'b0 : node155;
											assign node155 = (inp[6]) ? 1'b0 : node156;
												assign node156 = (inp[3]) ? 1'b0 : 1'b1;
									assign node161 = (inp[7]) ? 1'b0 : node162;
										assign node162 = (inp[13]) ? 1'b0 : 1'b1;
				assign node166 = (inp[11]) ? node258 : node167;
					assign node167 = (inp[9]) ? node209 : node168;
						assign node168 = (inp[1]) ? node178 : node169;
							assign node169 = (inp[12]) ? node171 : 1'b1;
								assign node171 = (inp[14]) ? node173 : 1'b1;
									assign node173 = (inp[6]) ? node175 : 1'b1;
										assign node175 = (inp[0]) ? 1'b0 : 1'b1;
							assign node178 = (inp[6]) ? node188 : node179;
								assign node179 = (inp[5]) ? node181 : 1'b1;
									assign node181 = (inp[13]) ? node183 : 1'b1;
										assign node183 = (inp[3]) ? 1'b1 : node184;
											assign node184 = (inp[0]) ? 1'b0 : 1'b1;
								assign node188 = (inp[14]) ? node198 : node189;
									assign node189 = (inp[3]) ? node191 : 1'b1;
										assign node191 = (inp[7]) ? node193 : 1'b1;
											assign node193 = (inp[0]) ? 1'b0 : node194;
												assign node194 = (inp[13]) ? 1'b0 : 1'b1;
									assign node198 = (inp[8]) ? node204 : node199;
										assign node199 = (inp[3]) ? node201 : 1'b1;
											assign node201 = (inp[12]) ? 1'b0 : 1'b1;
										assign node204 = (inp[13]) ? 1'b0 : node205;
											assign node205 = (inp[5]) ? 1'b1 : 1'b0;
						assign node209 = (inp[3]) ? node233 : node210;
							assign node210 = (inp[6]) ? node212 : 1'b1;
								assign node212 = (inp[5]) ? node220 : node213;
									assign node213 = (inp[7]) ? node215 : 1'b1;
										assign node215 = (inp[14]) ? node217 : 1'b1;
											assign node217 = (inp[13]) ? 1'b0 : 1'b1;
									assign node220 = (inp[14]) ? node228 : node221;
										assign node221 = (inp[1]) ? node223 : 1'b1;
											assign node223 = (inp[7]) ? 1'b0 : node224;
												assign node224 = (inp[12]) ? 1'b0 : 1'b1;
										assign node228 = (inp[12]) ? 1'b0 : node229;
											assign node229 = (inp[8]) ? 1'b0 : 1'b1;
							assign node233 = (inp[13]) ? node253 : node234;
								assign node234 = (inp[7]) ? node242 : node235;
									assign node235 = (inp[1]) ? node237 : 1'b1;
										assign node237 = (inp[5]) ? node239 : 1'b1;
											assign node239 = (inp[12]) ? 1'b0 : 1'b1;
									assign node242 = (inp[14]) ? 1'b0 : node243;
										assign node243 = (inp[12]) ? node245 : 1'b1;
											assign node245 = (inp[8]) ? 1'b0 : node246;
												assign node246 = (inp[0]) ? node248 : 1'b1;
													assign node248 = (inp[5]) ? 1'b0 : 1'b1;
								assign node253 = (inp[5]) ? 1'b0 : node254;
									assign node254 = (inp[12]) ? 1'b0 : 1'b1;
					assign node258 = (inp[5]) ? node320 : node259;
						assign node259 = (inp[8]) ? node285 : node260;
							assign node260 = (inp[1]) ? node270 : node261;
								assign node261 = (inp[14]) ? node263 : 1'b1;
									assign node263 = (inp[12]) ? node265 : 1'b1;
										assign node265 = (inp[9]) ? node267 : 1'b1;
											assign node267 = (inp[3]) ? 1'b0 : 1'b1;
								assign node270 = (inp[7]) ? node276 : node271;
									assign node271 = (inp[13]) ? node273 : 1'b1;
										assign node273 = (inp[6]) ? 1'b0 : 1'b1;
									assign node276 = (inp[12]) ? node280 : node277;
										assign node277 = (inp[9]) ? 1'b0 : 1'b1;
										assign node280 = (inp[6]) ? 1'b0 : node281;
											assign node281 = (inp[14]) ? 1'b0 : 1'b1;
							assign node285 = (inp[0]) ? node309 : node286;
								assign node286 = (inp[7]) ? node292 : node287;
									assign node287 = (inp[1]) ? node289 : 1'b1;
										assign node289 = (inp[6]) ? 1'b0 : 1'b1;
									assign node292 = (inp[12]) ? node298 : node293;
										assign node293 = (inp[13]) ? node295 : 1'b1;
											assign node295 = (inp[6]) ? 1'b0 : 1'b1;
										assign node298 = (inp[3]) ? 1'b0 : node299;
											assign node299 = (inp[6]) ? node303 : node300;
												assign node300 = (inp[9]) ? 1'b0 : 1'b1;
												assign node303 = (inp[13]) ? 1'b0 : node304;
													assign node304 = (inp[1]) ? 1'b0 : 1'b1;
								assign node309 = (inp[13]) ? 1'b0 : node310;
									assign node310 = (inp[14]) ? 1'b0 : node311;
										assign node311 = (inp[9]) ? node313 : 1'b1;
											assign node313 = (inp[7]) ? node315 : 1'b1;
												assign node315 = (inp[6]) ? 1'b0 : 1'b1;
						assign node320 = (inp[1]) ? node364 : node321;
							assign node321 = (inp[8]) ? node345 : node322;
								assign node322 = (inp[3]) ? node334 : node323;
									assign node323 = (inp[9]) ? node325 : 1'b1;
										assign node325 = (inp[14]) ? node327 : 1'b1;
											assign node327 = (inp[0]) ? node329 : 1'b1;
												assign node329 = (inp[12]) ? 1'b0 : node330;
													assign node330 = (inp[6]) ? 1'b0 : 1'b1;
									assign node334 = (inp[9]) ? node340 : node335;
										assign node335 = (inp[12]) ? node337 : 1'b1;
											assign node337 = (inp[7]) ? 1'b0 : 1'b1;
										assign node340 = (inp[12]) ? 1'b0 : node341;
											assign node341 = (inp[14]) ? 1'b0 : 1'b1;
								assign node345 = (inp[0]) ? node357 : node346;
									assign node346 = (inp[6]) ? node352 : node347;
										assign node347 = (inp[14]) ? node349 : 1'b1;
											assign node349 = (inp[12]) ? 1'b0 : 1'b1;
										assign node352 = (inp[3]) ? 1'b0 : node353;
											assign node353 = (inp[13]) ? 1'b0 : 1'b1;
									assign node357 = (inp[12]) ? 1'b0 : node358;
										assign node358 = (inp[7]) ? 1'b0 : node359;
											assign node359 = (inp[14]) ? 1'b0 : 1'b1;
							assign node364 = (inp[6]) ? node382 : node365;
								assign node365 = (inp[12]) ? node371 : node366;
									assign node366 = (inp[13]) ? node368 : 1'b1;
										assign node368 = (inp[14]) ? 1'b0 : 1'b1;
									assign node371 = (inp[0]) ? 1'b0 : node372;
										assign node372 = (inp[9]) ? node376 : node373;
											assign node373 = (inp[3]) ? 1'b0 : 1'b1;
											assign node376 = (inp[14]) ? 1'b0 : node377;
												assign node377 = (inp[7]) ? 1'b0 : 1'b1;
								assign node382 = (inp[9]) ? 1'b0 : node383;
									assign node383 = (inp[13]) ? 1'b0 : node384;
										assign node384 = (inp[3]) ? 1'b0 : node385;
											assign node385 = (inp[12]) ? 1'b0 : 1'b1;
			assign node391 = (inp[13]) ? node657 : node392;
				assign node392 = (inp[11]) ? node502 : node393;
					assign node393 = (inp[12]) ? node417 : node394;
						assign node394 = (inp[10]) ? node396 : 1'b1;
							assign node396 = (inp[9]) ? node398 : 1'b1;
								assign node398 = (inp[5]) ? node406 : node399;
									assign node399 = (inp[1]) ? node401 : 1'b1;
										assign node401 = (inp[6]) ? node403 : 1'b1;
											assign node403 = (inp[0]) ? 1'b0 : 1'b1;
									assign node406 = (inp[0]) ? node412 : node407;
										assign node407 = (inp[8]) ? 1'b1 : node408;
											assign node408 = (inp[7]) ? 1'b0 : 1'b1;
										assign node412 = (inp[3]) ? 1'b0 : node413;
											assign node413 = (inp[6]) ? 1'b1 : 1'b0;
						assign node417 = (inp[8]) ? node451 : node418;
							assign node418 = (inp[0]) ? node428 : node419;
								assign node419 = (inp[6]) ? node421 : 1'b1;
									assign node421 = (inp[14]) ? node423 : 1'b1;
										assign node423 = (inp[5]) ? node425 : 1'b1;
											assign node425 = (inp[7]) ? 1'b0 : 1'b1;
								assign node428 = (inp[9]) ? node436 : node429;
									assign node429 = (inp[6]) ? node431 : 1'b1;
										assign node431 = (inp[3]) ? node433 : 1'b1;
											assign node433 = (inp[5]) ? 1'b0 : 1'b1;
									assign node436 = (inp[14]) ? node446 : node437;
										assign node437 = (inp[5]) ? node439 : 1'b1;
											assign node439 = (inp[6]) ? 1'b0 : node440;
												assign node440 = (inp[10]) ? node442 : 1'b1;
													assign node442 = (inp[1]) ? 1'b0 : 1'b1;
										assign node446 = (inp[10]) ? 1'b0 : node447;
											assign node447 = (inp[3]) ? 1'b0 : 1'b1;
							assign node451 = (inp[14]) ? node469 : node452;
								assign node452 = (inp[5]) ? node454 : 1'b1;
									assign node454 = (inp[1]) ? node464 : node455;
										assign node455 = (inp[6]) ? node457 : 1'b1;
											assign node457 = (inp[7]) ? node459 : 1'b1;
												assign node459 = (inp[9]) ? 1'b0 : node460;
													assign node460 = (inp[3]) ? 1'b0 : 1'b1;
										assign node464 = (inp[3]) ? 1'b0 : node465;
											assign node465 = (inp[6]) ? 1'b0 : 1'b1;
								assign node469 = (inp[7]) ? node487 : node470;
									assign node470 = (inp[5]) ? node482 : node471;
										assign node471 = (inp[10]) ? node477 : node472;
											assign node472 = (inp[3]) ? 1'b1 : node473;
												assign node473 = (inp[6]) ? 1'b0 : 1'b1;
											assign node477 = (inp[1]) ? 1'b0 : node478;
												assign node478 = (inp[9]) ? 1'b0 : 1'b1;
										assign node482 = (inp[9]) ? 1'b0 : node483;
											assign node483 = (inp[1]) ? 1'b0 : 1'b1;
									assign node487 = (inp[6]) ? 1'b0 : node488;
										assign node488 = (inp[1]) ? node494 : node489;
											assign node489 = (inp[3]) ? node491 : 1'b1;
												assign node491 = (inp[9]) ? 1'b0 : 1'b1;
											assign node494 = (inp[10]) ? 1'b0 : node495;
												assign node495 = (inp[5]) ? node497 : 1'b0;
													assign node497 = (inp[9]) ? 1'b0 : 1'b1;
					assign node502 = (inp[6]) ? node578 : node503;
						assign node503 = (inp[0]) ? node545 : node504;
							assign node504 = (inp[14]) ? node522 : node505;
								assign node505 = (inp[10]) ? node507 : 1'b1;
									assign node507 = (inp[3]) ? node509 : 1'b1;
										assign node509 = (inp[9]) ? node517 : node510;
											assign node510 = (inp[1]) ? node512 : 1'b1;
												assign node512 = (inp[8]) ? node514 : 1'b1;
													assign node514 = (inp[12]) ? 1'b0 : 1'b1;
											assign node517 = (inp[5]) ? 1'b0 : node518;
												assign node518 = (inp[12]) ? 1'b0 : 1'b1;
								assign node522 = (inp[12]) ? node534 : node523;
									assign node523 = (inp[10]) ? node525 : 1'b1;
										assign node525 = (inp[5]) ? node527 : 1'b1;
											assign node527 = (inp[9]) ? 1'b0 : node528;
												assign node528 = (inp[7]) ? node530 : 1'b1;
													assign node530 = (inp[3]) ? 1'b0 : 1'b1;
									assign node534 = (inp[7]) ? node540 : node535;
										assign node535 = (inp[8]) ? node537 : 1'b1;
											assign node537 = (inp[5]) ? 1'b0 : 1'b1;
										assign node540 = (inp[1]) ? 1'b0 : node541;
											assign node541 = (inp[5]) ? 1'b0 : 1'b1;
							assign node545 = (inp[7]) ? node565 : node546;
								assign node546 = (inp[8]) ? node554 : node547;
									assign node547 = (inp[3]) ? node549 : 1'b1;
										assign node549 = (inp[9]) ? node551 : 1'b1;
											assign node551 = (inp[5]) ? 1'b0 : 1'b1;
									assign node554 = (inp[14]) ? node560 : node555;
										assign node555 = (inp[5]) ? node557 : 1'b1;
											assign node557 = (inp[10]) ? 1'b0 : 1'b1;
										assign node560 = (inp[12]) ? 1'b0 : node561;
											assign node561 = (inp[5]) ? 1'b0 : 1'b1;
								assign node565 = (inp[14]) ? 1'b0 : node566;
									assign node566 = (inp[12]) ? node572 : node567;
										assign node567 = (inp[10]) ? node569 : 1'b1;
											assign node569 = (inp[3]) ? 1'b0 : 1'b1;
										assign node572 = (inp[8]) ? 1'b0 : node573;
											assign node573 = (inp[1]) ? 1'b1 : 1'b0;
						assign node578 = (inp[0]) ? node618 : node579;
							assign node579 = (inp[10]) ? node595 : node580;
								assign node580 = (inp[8]) ? node588 : node581;
									assign node581 = (inp[7]) ? node583 : 1'b1;
										assign node583 = (inp[1]) ? node585 : 1'b1;
											assign node585 = (inp[5]) ? 1'b0 : 1'b1;
									assign node588 = (inp[1]) ? 1'b0 : node589;
										assign node589 = (inp[5]) ? 1'b1 : node590;
											assign node590 = (inp[3]) ? 1'b0 : 1'b1;
								assign node595 = (inp[9]) ? node611 : node596;
									assign node596 = (inp[12]) ? node602 : node597;
										assign node597 = (inp[8]) ? node599 : 1'b1;
											assign node599 = (inp[1]) ? 1'b0 : 1'b1;
										assign node602 = (inp[7]) ? 1'b0 : node603;
											assign node603 = (inp[1]) ? node605 : 1'b1;
												assign node605 = (inp[3]) ? 1'b0 : node606;
													assign node606 = (inp[5]) ? 1'b0 : 1'b1;
									assign node611 = (inp[1]) ? 1'b0 : node612;
										assign node612 = (inp[8]) ? 1'b0 : node613;
											assign node613 = (inp[7]) ? 1'b0 : 1'b1;
							assign node618 = (inp[12]) ? node648 : node619;
								assign node619 = (inp[9]) ? node637 : node620;
									assign node620 = (inp[3]) ? node630 : node621;
										assign node621 = (inp[8]) ? node623 : 1'b1;
											assign node623 = (inp[7]) ? node625 : 1'b1;
												assign node625 = (inp[14]) ? 1'b0 : node626;
													assign node626 = (inp[10]) ? 1'b0 : 1'b1;
										assign node630 = (inp[5]) ? 1'b0 : node631;
											assign node631 = (inp[10]) ? 1'b0 : node632;
												assign node632 = (inp[1]) ? 1'b0 : 1'b1;
									assign node637 = (inp[7]) ? 1'b0 : node638;
										assign node638 = (inp[5]) ? 1'b0 : node639;
											assign node639 = (inp[14]) ? 1'b0 : node640;
												assign node640 = (inp[1]) ? node642 : 1'b1;
													assign node642 = (inp[10]) ? 1'b0 : 1'b1;
								assign node648 = (inp[14]) ? 1'b0 : node649;
									assign node649 = (inp[9]) ? 1'b0 : node650;
										assign node650 = (inp[3]) ? 1'b0 : node651;
											assign node651 = (inp[7]) ? 1'b0 : 1'b1;
				assign node657 = (inp[3]) ? node799 : node658;
					assign node658 = (inp[12]) ? node728 : node659;
						assign node659 = (inp[14]) ? node693 : node660;
							assign node660 = (inp[9]) ? node670 : node661;
								assign node661 = (inp[10]) ? node663 : 1'b1;
									assign node663 = (inp[1]) ? node665 : 1'b1;
										assign node665 = (inp[7]) ? node667 : 1'b1;
											assign node667 = (inp[5]) ? 1'b0 : 1'b1;
								assign node670 = (inp[0]) ? node680 : node671;
									assign node671 = (inp[8]) ? node673 : 1'b1;
										assign node673 = (inp[1]) ? 1'b0 : node674;
											assign node674 = (inp[5]) ? node676 : 1'b1;
												assign node676 = (inp[6]) ? 1'b1 : 1'b0;
									assign node680 = (inp[5]) ? node688 : node681;
										assign node681 = (inp[6]) ? node683 : 1'b1;
											assign node683 = (inp[11]) ? 1'b0 : node684;
												assign node684 = (inp[1]) ? 1'b0 : 1'b1;
										assign node688 = (inp[1]) ? 1'b0 : node689;
											assign node689 = (inp[10]) ? 1'b0 : 1'b1;
							assign node693 = (inp[0]) ? node709 : node694;
								assign node694 = (inp[6]) ? node702 : node695;
									assign node695 = (inp[10]) ? node697 : 1'b1;
										assign node697 = (inp[8]) ? node699 : 1'b1;
											assign node699 = (inp[7]) ? 1'b0 : 1'b1;
									assign node702 = (inp[7]) ? node704 : 1'b1;
										assign node704 = (inp[8]) ? 1'b0 : node705;
											assign node705 = (inp[9]) ? 1'b0 : 1'b1;
								assign node709 = (inp[1]) ? node723 : node710;
									assign node710 = (inp[9]) ? node716 : node711;
										assign node711 = (inp[8]) ? node713 : 1'b1;
											assign node713 = (inp[11]) ? 1'b0 : 1'b1;
										assign node716 = (inp[10]) ? 1'b0 : node717;
											assign node717 = (inp[7]) ? 1'b0 : node718;
												assign node718 = (inp[8]) ? 1'b0 : 1'b1;
									assign node723 = (inp[10]) ? 1'b0 : node724;
										assign node724 = (inp[5]) ? 1'b0 : 1'b1;
						assign node728 = (inp[9]) ? node760 : node729;
							assign node729 = (inp[1]) ? node743 : node730;
								assign node730 = (inp[10]) ? node736 : node731;
									assign node731 = (inp[5]) ? node733 : 1'b1;
										assign node733 = (inp[0]) ? 1'b0 : 1'b1;
									assign node736 = (inp[6]) ? 1'b0 : node737;
										assign node737 = (inp[8]) ? node739 : 1'b1;
											assign node739 = (inp[11]) ? 1'b0 : 1'b1;
								assign node743 = (inp[7]) ? node753 : node744;
									assign node744 = (inp[11]) ? node748 : node745;
										assign node745 = (inp[6]) ? 1'b0 : 1'b1;
										assign node748 = (inp[8]) ? 1'b0 : node749;
											assign node749 = (inp[10]) ? 1'b0 : 1'b1;
									assign node753 = (inp[14]) ? 1'b0 : node754;
										assign node754 = (inp[11]) ? 1'b0 : node755;
											assign node755 = (inp[0]) ? 1'b0 : 1'b1;
							assign node760 = (inp[7]) ? node790 : node761;
								assign node761 = (inp[10]) ? node783 : node762;
									assign node762 = (inp[11]) ? node772 : node763;
										assign node763 = (inp[1]) ? node765 : 1'b1;
											assign node765 = (inp[14]) ? node767 : 1'b1;
												assign node767 = (inp[6]) ? node769 : 1'b0;
													assign node769 = (inp[8]) ? 1'b0 : 1'b1;
										assign node772 = (inp[0]) ? 1'b0 : node773;
											assign node773 = (inp[1]) ? 1'b0 : node774;
												assign node774 = (inp[8]) ? node776 : 1'b1;
													assign node776 = (inp[14]) ? 1'b0 : node777;
														assign node777 = (inp[6]) ? 1'b0 : 1'b1;
									assign node783 = (inp[6]) ? 1'b0 : node784;
										assign node784 = (inp[8]) ? 1'b0 : node785;
											assign node785 = (inp[14]) ? 1'b0 : 1'b1;
								assign node790 = (inp[5]) ? 1'b0 : node791;
									assign node791 = (inp[14]) ? 1'b0 : node792;
										assign node792 = (inp[6]) ? 1'b0 : node793;
											assign node793 = (inp[0]) ? 1'b0 : 1'b1;
					assign node799 = (inp[7]) ? node871 : node800;
						assign node800 = (inp[11]) ? node838 : node801;
							assign node801 = (inp[5]) ? node815 : node802;
								assign node802 = (inp[10]) ? node804 : 1'b1;
									assign node804 = (inp[6]) ? node810 : node805;
										assign node805 = (inp[12]) ? node807 : 1'b1;
											assign node807 = (inp[8]) ? 1'b0 : 1'b1;
										assign node810 = (inp[1]) ? 1'b0 : node811;
											assign node811 = (inp[0]) ? 1'b0 : 1'b1;
								assign node815 = (inp[14]) ? node833 : node816;
									assign node816 = (inp[8]) ? node822 : node817;
										assign node817 = (inp[0]) ? node819 : 1'b1;
											assign node819 = (inp[9]) ? 1'b0 : 1'b1;
										assign node822 = (inp[6]) ? node828 : node823;
											assign node823 = (inp[1]) ? node825 : 1'b1;
												assign node825 = (inp[10]) ? 1'b0 : 1'b1;
											assign node828 = (inp[12]) ? 1'b0 : node829;
												assign node829 = (inp[10]) ? 1'b0 : 1'b1;
									assign node833 = (inp[1]) ? 1'b0 : node834;
										assign node834 = (inp[6]) ? 1'b0 : 1'b1;
							assign node838 = (inp[8]) ? node864 : node839;
								assign node839 = (inp[6]) ? node859 : node840;
									assign node840 = (inp[9]) ? node850 : node841;
										assign node841 = (inp[10]) ? node843 : 1'b1;
											assign node843 = (inp[12]) ? 1'b0 : node844;
												assign node844 = (inp[14]) ? node846 : 1'b1;
													assign node846 = (inp[5]) ? 1'b0 : 1'b1;
										assign node850 = (inp[1]) ? 1'b0 : node851;
											assign node851 = (inp[5]) ? node853 : 1'b1;
												assign node853 = (inp[14]) ? 1'b0 : node854;
													assign node854 = (inp[10]) ? 1'b0 : 1'b1;
									assign node859 = (inp[1]) ? 1'b0 : node860;
										assign node860 = (inp[10]) ? 1'b0 : 1'b1;
								assign node864 = (inp[6]) ? node866 : 1'b0;
									assign node866 = (inp[9]) ? 1'b0 : node867;
										assign node867 = (inp[0]) ? 1'b0 : 1'b1;
						assign node871 = (inp[8]) ? node909 : node872;
							assign node872 = (inp[9]) ? node896 : node873;
								assign node873 = (inp[14]) ? node889 : node874;
									assign node874 = (inp[6]) ? node880 : node875;
										assign node875 = (inp[12]) ? node877 : 1'b1;
											assign node877 = (inp[5]) ? 1'b0 : 1'b1;
										assign node880 = (inp[10]) ? node884 : node881;
											assign node881 = (inp[11]) ? 1'b0 : 1'b1;
											assign node884 = (inp[5]) ? 1'b0 : node885;
												assign node885 = (inp[11]) ? 1'b0 : 1'b1;
									assign node889 = (inp[11]) ? 1'b0 : node890;
										assign node890 = (inp[6]) ? 1'b0 : node891;
											assign node891 = (inp[10]) ? 1'b0 : 1'b1;
								assign node896 = (inp[5]) ? 1'b0 : node897;
									assign node897 = (inp[10]) ? 1'b0 : node898;
										assign node898 = (inp[1]) ? 1'b0 : node899;
											assign node899 = (inp[11]) ? 1'b0 : node900;
												assign node900 = (inp[12]) ? node902 : 1'b1;
													assign node902 = (inp[6]) ? 1'b0 : 1'b1;
							assign node909 = (inp[14]) ? 1'b0 : node910;
								assign node910 = (inp[12]) ? 1'b0 : node911;
									assign node911 = (inp[10]) ? 1'b0 : node912;
										assign node912 = (inp[9]) ? 1'b0 : node913;
											assign node913 = (inp[5]) ? node915 : 1'b1;
												assign node915 = (inp[6]) ? 1'b0 : node916;
													assign node916 = (inp[0]) ? 1'b0 : 1'b1;
		assign node924 = (inp[5]) ? node1394 : node925;
			assign node925 = (inp[13]) ? node1157 : node926;
				assign node926 = (inp[6]) ? node1030 : node927;
					assign node927 = (inp[12]) ? node957 : node928;
						assign node928 = (inp[11]) ? node930 : 1'b1;
							assign node930 = (inp[14]) ? node932 : 1'b1;
								assign node932 = (inp[9]) ? node938 : node933;
									assign node933 = (inp[3]) ? node935 : 1'b1;
										assign node935 = (inp[2]) ? 1'b0 : 1'b1;
									assign node938 = (inp[2]) ? node948 : node939;
										assign node939 = (inp[8]) ? node941 : 1'b1;
											assign node941 = (inp[3]) ? node943 : 1'b1;
												assign node943 = (inp[7]) ? 1'b0 : node944;
													assign node944 = (inp[1]) ? 1'b0 : 1'b1;
										assign node948 = (inp[10]) ? 1'b0 : node949;
											assign node949 = (inp[8]) ? 1'b0 : node950;
												assign node950 = (inp[7]) ? node952 : 1'b1;
													assign node952 = (inp[3]) ? 1'b0 : 1'b1;
						assign node957 = (inp[0]) ? node987 : node958;
							assign node958 = (inp[8]) ? node972 : node959;
								assign node959 = (inp[10]) ? node961 : 1'b1;
									assign node961 = (inp[3]) ? node963 : 1'b1;
										assign node963 = (inp[14]) ? 1'b0 : node964;
											assign node964 = (inp[7]) ? node966 : 1'b1;
												assign node966 = (inp[11]) ? node968 : 1'b1;
													assign node968 = (inp[2]) ? 1'b0 : 1'b1;
								assign node972 = (inp[9]) ? node980 : node973;
									assign node973 = (inp[7]) ? node975 : 1'b1;
										assign node975 = (inp[3]) ? node977 : 1'b1;
											assign node977 = (inp[1]) ? 1'b0 : 1'b1;
									assign node980 = (inp[14]) ? 1'b0 : node981;
										assign node981 = (inp[7]) ? node983 : 1'b1;
											assign node983 = (inp[11]) ? 1'b0 : 1'b1;
							assign node987 = (inp[1]) ? node1007 : node988;
								assign node988 = (inp[7]) ? node996 : node989;
									assign node989 = (inp[11]) ? node991 : 1'b1;
										assign node991 = (inp[2]) ? node993 : 1'b1;
											assign node993 = (inp[14]) ? 1'b0 : 1'b1;
									assign node996 = (inp[8]) ? node998 : 1'b1;
										assign node998 = (inp[11]) ? 1'b0 : node999;
											assign node999 = (inp[2]) ? node1001 : 1'b1;
												assign node1001 = (inp[14]) ? 1'b0 : node1002;
													assign node1002 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1007 = (inp[2]) ? node1017 : node1008;
									assign node1008 = (inp[9]) ? node1014 : node1009;
										assign node1009 = (inp[10]) ? node1011 : 1'b1;
											assign node1011 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1014 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1017 = (inp[3]) ? 1'b0 : node1018;
										assign node1018 = (inp[9]) ? 1'b0 : node1019;
											assign node1019 = (inp[7]) ? node1021 : 1'b1;
												assign node1021 = (inp[14]) ? 1'b0 : node1022;
													assign node1022 = (inp[10]) ? 1'b0 : node1023;
														assign node1023 = (inp[8]) ? 1'b0 : 1'b1;
					assign node1030 = (inp[2]) ? node1092 : node1031;
						assign node1031 = (inp[9]) ? node1059 : node1032;
							assign node1032 = (inp[0]) ? node1034 : 1'b1;
								assign node1034 = (inp[1]) ? node1046 : node1035;
									assign node1035 = (inp[11]) ? node1037 : 1'b1;
										assign node1037 = (inp[10]) ? 1'b0 : node1038;
											assign node1038 = (inp[12]) ? node1040 : 1'b1;
												assign node1040 = (inp[3]) ? node1042 : 1'b1;
													assign node1042 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1046 = (inp[10]) ? node1054 : node1047;
										assign node1047 = (inp[11]) ? node1049 : 1'b1;
											assign node1049 = (inp[8]) ? node1051 : 1'b1;
												assign node1051 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1054 = (inp[8]) ? 1'b0 : node1055;
											assign node1055 = (inp[14]) ? 1'b0 : 1'b1;
							assign node1059 = (inp[1]) ? node1081 : node1060;
								assign node1060 = (inp[8]) ? node1070 : node1061;
									assign node1061 = (inp[3]) ? node1063 : 1'b1;
										assign node1063 = (inp[7]) ? node1065 : 1'b1;
											assign node1065 = (inp[12]) ? 1'b0 : node1066;
												assign node1066 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1070 = (inp[7]) ? node1076 : node1071;
										assign node1071 = (inp[12]) ? node1073 : 1'b1;
											assign node1073 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1076 = (inp[12]) ? 1'b0 : node1077;
											assign node1077 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1081 = (inp[14]) ? 1'b0 : node1082;
									assign node1082 = (inp[0]) ? node1086 : node1083;
										assign node1083 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1086 = (inp[8]) ? 1'b0 : node1087;
											assign node1087 = (inp[7]) ? 1'b1 : 1'b0;
						assign node1092 = (inp[11]) ? node1128 : node1093;
							assign node1093 = (inp[12]) ? node1111 : node1094;
								assign node1094 = (inp[9]) ? node1102 : node1095;
									assign node1095 = (inp[7]) ? node1097 : 1'b1;
										assign node1097 = (inp[10]) ? node1099 : 1'b1;
											assign node1099 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1102 = (inp[1]) ? node1104 : 1'b1;
										assign node1104 = (inp[3]) ? 1'b0 : node1105;
											assign node1105 = (inp[14]) ? node1107 : 1'b1;
												assign node1107 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1111 = (inp[7]) ? node1119 : node1112;
									assign node1112 = (inp[0]) ? 1'b0 : node1113;
										assign node1113 = (inp[3]) ? node1115 : 1'b1;
											assign node1115 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1119 = (inp[1]) ? 1'b0 : node1120;
										assign node1120 = (inp[8]) ? 1'b0 : node1121;
											assign node1121 = (inp[14]) ? node1123 : 1'b0;
												assign node1123 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1128 = (inp[1]) ? node1148 : node1129;
								assign node1129 = (inp[0]) ? node1143 : node1130;
									assign node1130 = (inp[7]) ? node1136 : node1131;
										assign node1131 = (inp[9]) ? node1133 : 1'b1;
											assign node1133 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1136 = (inp[10]) ? 1'b0 : node1137;
											assign node1137 = (inp[8]) ? node1139 : 1'b1;
												assign node1139 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1143 = (inp[9]) ? 1'b0 : node1144;
										assign node1144 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1148 = (inp[8]) ? 1'b0 : node1149;
									assign node1149 = (inp[3]) ? 1'b0 : node1150;
										assign node1150 = (inp[10]) ? 1'b0 : node1151;
											assign node1151 = (inp[9]) ? 1'b0 : 1'b1;
				assign node1157 = (inp[2]) ? node1279 : node1158;
					assign node1158 = (inp[12]) ? node1222 : node1159;
						assign node1159 = (inp[10]) ? node1189 : node1160;
							assign node1160 = (inp[7]) ? node1172 : node1161;
								assign node1161 = (inp[6]) ? node1163 : 1'b1;
									assign node1163 = (inp[8]) ? node1165 : 1'b1;
										assign node1165 = (inp[11]) ? 1'b0 : node1166;
											assign node1166 = (inp[14]) ? node1168 : 1'b1;
												assign node1168 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1172 = (inp[0]) ? node1186 : node1173;
									assign node1173 = (inp[9]) ? node1183 : node1174;
										assign node1174 = (inp[6]) ? 1'b1 : node1175;
											assign node1175 = (inp[1]) ? node1177 : 1'b1;
												assign node1177 = (inp[11]) ? node1179 : 1'b1;
													assign node1179 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1183 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1186 = (inp[1]) ? 1'b0 : 1'b1;
							assign node1189 = (inp[1]) ? node1209 : node1190;
								assign node1190 = (inp[14]) ? node1198 : node1191;
									assign node1191 = (inp[7]) ? node1193 : 1'b1;
										assign node1193 = (inp[8]) ? node1195 : 1'b1;
											assign node1195 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1198 = (inp[0]) ? node1204 : node1199;
										assign node1199 = (inp[6]) ? node1201 : 1'b1;
											assign node1201 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1204 = (inp[9]) ? node1206 : 1'b0;
											assign node1206 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1209 = (inp[6]) ? 1'b0 : node1210;
									assign node1210 = (inp[11]) ? node1216 : node1211;
										assign node1211 = (inp[8]) ? node1213 : 1'b1;
											assign node1213 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1216 = (inp[9]) ? 1'b0 : node1217;
											assign node1217 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1222 = (inp[9]) ? node1256 : node1223;
							assign node1223 = (inp[10]) ? node1239 : node1224;
								assign node1224 = (inp[1]) ? node1232 : node1225;
									assign node1225 = (inp[3]) ? node1227 : 1'b1;
										assign node1227 = (inp[0]) ? node1229 : 1'b1;
											assign node1229 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1232 = (inp[6]) ? 1'b0 : node1233;
										assign node1233 = (inp[7]) ? node1235 : 1'b1;
											assign node1235 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1239 = (inp[11]) ? node1249 : node1240;
									assign node1240 = (inp[8]) ? node1246 : node1241;
										assign node1241 = (inp[14]) ? node1243 : 1'b1;
											assign node1243 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1246 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1249 = (inp[14]) ? 1'b0 : node1250;
										assign node1250 = (inp[3]) ? 1'b0 : node1251;
											assign node1251 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1256 = (inp[1]) ? node1272 : node1257;
								assign node1257 = (inp[8]) ? node1265 : node1258;
									assign node1258 = (inp[11]) ? node1260 : 1'b1;
										assign node1260 = (inp[0]) ? 1'b0 : node1261;
											assign node1261 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1265 = (inp[7]) ? 1'b0 : node1266;
										assign node1266 = (inp[11]) ? node1268 : 1'b0;
											assign node1268 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1272 = (inp[10]) ? 1'b0 : node1273;
									assign node1273 = (inp[0]) ? 1'b0 : node1274;
										assign node1274 = (inp[6]) ? 1'b0 : 1'b1;
					assign node1279 = (inp[6]) ? node1345 : node1280;
						assign node1280 = (inp[14]) ? node1314 : node1281;
							assign node1281 = (inp[12]) ? node1303 : node1282;
								assign node1282 = (inp[3]) ? node1290 : node1283;
									assign node1283 = (inp[7]) ? node1285 : 1'b1;
										assign node1285 = (inp[0]) ? node1287 : 1'b1;
											assign node1287 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1290 = (inp[10]) ? node1298 : node1291;
										assign node1291 = (inp[0]) ? node1293 : 1'b1;
											assign node1293 = (inp[1]) ? 1'b0 : node1294;
												assign node1294 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1298 = (inp[9]) ? 1'b0 : node1299;
											assign node1299 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1303 = (inp[8]) ? 1'b0 : node1304;
									assign node1304 = (inp[11]) ? node1310 : node1305;
										assign node1305 = (inp[7]) ? node1307 : 1'b1;
											assign node1307 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1310 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1314 = (inp[8]) ? node1336 : node1315;
								assign node1315 = (inp[11]) ? node1329 : node1316;
									assign node1316 = (inp[12]) ? node1324 : node1317;
										assign node1317 = (inp[0]) ? node1319 : 1'b1;
											assign node1319 = (inp[9]) ? 1'b0 : node1320;
												assign node1320 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1324 = (inp[7]) ? 1'b0 : node1325;
											assign node1325 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1329 = (inp[3]) ? 1'b0 : node1330;
										assign node1330 = (inp[10]) ? 1'b0 : node1331;
											assign node1331 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1336 = (inp[7]) ? 1'b0 : node1337;
									assign node1337 = (inp[3]) ? 1'b0 : node1338;
										assign node1338 = (inp[10]) ? 1'b0 : node1339;
											assign node1339 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1345 = (inp[0]) ? node1383 : node1346;
							assign node1346 = (inp[7]) ? node1366 : node1347;
								assign node1347 = (inp[9]) ? node1359 : node1348;
									assign node1348 = (inp[8]) ? node1354 : node1349;
										assign node1349 = (inp[12]) ? node1351 : 1'b1;
											assign node1351 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1354 = (inp[11]) ? 1'b0 : node1355;
											assign node1355 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1359 = (inp[14]) ? 1'b0 : node1360;
										assign node1360 = (inp[1]) ? 1'b0 : node1361;
											assign node1361 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1366 = (inp[8]) ? 1'b0 : node1367;
									assign node1367 = (inp[11]) ? 1'b0 : node1368;
										assign node1368 = (inp[12]) ? node1376 : node1369;
											assign node1369 = (inp[3]) ? 1'b0 : node1370;
												assign node1370 = (inp[9]) ? node1372 : 1'b1;
													assign node1372 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1376 = (inp[1]) ? 1'b0 : node1377;
												assign node1377 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1383 = (inp[8]) ? 1'b0 : node1384;
								assign node1384 = (inp[10]) ? 1'b0 : node1385;
									assign node1385 = (inp[3]) ? 1'b0 : node1386;
										assign node1386 = (inp[9]) ? 1'b0 : node1387;
											assign node1387 = (inp[7]) ? 1'b0 : 1'b1;
			assign node1394 = (inp[9]) ? node1610 : node1395;
				assign node1395 = (inp[1]) ? node1521 : node1396;
					assign node1396 = (inp[3]) ? node1456 : node1397;
						assign node1397 = (inp[6]) ? node1427 : node1398;
							assign node1398 = (inp[11]) ? node1406 : node1399;
								assign node1399 = (inp[10]) ? node1401 : 1'b1;
									assign node1401 = (inp[0]) ? node1403 : 1'b1;
										assign node1403 = (inp[14]) ? 1'b0 : 1'b1;
								assign node1406 = (inp[8]) ? node1408 : 1'b1;
									assign node1408 = (inp[10]) ? node1422 : node1409;
										assign node1409 = (inp[2]) ? node1411 : 1'b1;
											assign node1411 = (inp[14]) ? node1417 : node1412;
												assign node1412 = (inp[7]) ? node1414 : 1'b1;
													assign node1414 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1417 = (inp[7]) ? 1'b0 : node1418;
													assign node1418 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1422 = (inp[13]) ? 1'b0 : node1423;
											assign node1423 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1427 = (inp[2]) ? node1445 : node1428;
								assign node1428 = (inp[7]) ? node1434 : node1429;
									assign node1429 = (inp[13]) ? node1431 : 1'b1;
										assign node1431 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1434 = (inp[14]) ? node1440 : node1435;
										assign node1435 = (inp[8]) ? node1437 : 1'b1;
											assign node1437 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1440 = (inp[10]) ? 1'b0 : node1441;
											assign node1441 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1445 = (inp[13]) ? 1'b0 : node1446;
									assign node1446 = (inp[0]) ? node1450 : node1447;
										assign node1447 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1450 = (inp[14]) ? 1'b0 : node1451;
											assign node1451 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1456 = (inp[12]) ? node1482 : node1457;
							assign node1457 = (inp[0]) ? node1469 : node1458;
								assign node1458 = (inp[6]) ? node1460 : 1'b1;
									assign node1460 = (inp[8]) ? node1466 : node1461;
										assign node1461 = (inp[14]) ? node1463 : 1'b1;
											assign node1463 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1466 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1469 = (inp[13]) ? 1'b0 : node1470;
									assign node1470 = (inp[2]) ? node1476 : node1471;
										assign node1471 = (inp[7]) ? node1473 : 1'b1;
											assign node1473 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1476 = (inp[10]) ? 1'b0 : node1477;
											assign node1477 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1482 = (inp[14]) ? node1510 : node1483;
								assign node1483 = (inp[6]) ? node1501 : node1484;
									assign node1484 = (inp[8]) ? node1492 : node1485;
										assign node1485 = (inp[2]) ? node1487 : 1'b1;
											assign node1487 = (inp[11]) ? node1489 : 1'b1;
												assign node1489 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1492 = (inp[11]) ? 1'b0 : node1493;
											assign node1493 = (inp[13]) ? node1495 : 1'b1;
												assign node1495 = (inp[7]) ? 1'b0 : node1496;
													assign node1496 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1501 = (inp[10]) ? 1'b0 : node1502;
										assign node1502 = (inp[8]) ? node1504 : 1'b1;
											assign node1504 = (inp[0]) ? 1'b0 : node1505;
												assign node1505 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1510 = (inp[8]) ? 1'b0 : node1511;
									assign node1511 = (inp[7]) ? 1'b0 : node1512;
										assign node1512 = (inp[10]) ? node1514 : 1'b1;
											assign node1514 = (inp[2]) ? 1'b0 : node1515;
												assign node1515 = (inp[11]) ? 1'b0 : 1'b1;
					assign node1521 = (inp[12]) ? node1579 : node1522;
						assign node1522 = (inp[11]) ? node1550 : node1523;
							assign node1523 = (inp[13]) ? node1537 : node1524;
								assign node1524 = (inp[6]) ? node1526 : 1'b1;
									assign node1526 = (inp[14]) ? node1528 : 1'b1;
										assign node1528 = (inp[0]) ? 1'b0 : node1529;
											assign node1529 = (inp[10]) ? node1531 : 1'b1;
												assign node1531 = (inp[3]) ? 1'b0 : node1532;
													assign node1532 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1537 = (inp[2]) ? 1'b0 : node1538;
									assign node1538 = (inp[10]) ? node1544 : node1539;
										assign node1539 = (inp[3]) ? node1541 : 1'b1;
											assign node1541 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1544 = (inp[6]) ? 1'b0 : node1545;
											assign node1545 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1550 = (inp[6]) ? node1572 : node1551;
								assign node1551 = (inp[3]) ? node1565 : node1552;
									assign node1552 = (inp[7]) ? node1558 : node1553;
										assign node1553 = (inp[10]) ? node1555 : 1'b1;
											assign node1555 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1558 = (inp[0]) ? node1560 : 1'b1;
											assign node1560 = (inp[13]) ? 1'b0 : node1561;
												assign node1561 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1565 = (inp[7]) ? 1'b0 : node1566;
										assign node1566 = (inp[14]) ? 1'b0 : node1567;
											assign node1567 = (inp[8]) ? 1'b1 : 1'b0;
								assign node1572 = (inp[14]) ? 1'b0 : node1573;
									assign node1573 = (inp[8]) ? 1'b0 : node1574;
										assign node1574 = (inp[0]) ? 1'b0 : 1'b1;
						assign node1579 = (inp[10]) ? 1'b0 : node1580;
							assign node1580 = (inp[14]) ? node1600 : node1581;
								assign node1581 = (inp[7]) ? node1593 : node1582;
									assign node1582 = (inp[8]) ? node1588 : node1583;
										assign node1583 = (inp[2]) ? node1585 : 1'b1;
											assign node1585 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1588 = (inp[6]) ? 1'b0 : node1589;
											assign node1589 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1593 = (inp[2]) ? 1'b0 : node1594;
										assign node1594 = (inp[13]) ? 1'b0 : node1595;
											assign node1595 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1600 = (inp[11]) ? 1'b0 : node1601;
									assign node1601 = (inp[7]) ? 1'b0 : node1602;
										assign node1602 = (inp[3]) ? 1'b0 : node1603;
											assign node1603 = (inp[2]) ? 1'b0 : 1'b1;
				assign node1610 = (inp[8]) ? node1708 : node1611;
					assign node1611 = (inp[10]) ? node1671 : node1612;
						assign node1612 = (inp[3]) ? node1648 : node1613;
							assign node1613 = (inp[6]) ? node1625 : node1614;
								assign node1614 = (inp[1]) ? node1616 : 1'b1;
									assign node1616 = (inp[2]) ? 1'b0 : node1617;
										assign node1617 = (inp[11]) ? node1619 : 1'b1;
											assign node1619 = (inp[7]) ? 1'b0 : node1620;
												assign node1620 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1625 = (inp[12]) ? node1639 : node1626;
									assign node1626 = (inp[13]) ? node1632 : node1627;
										assign node1627 = (inp[2]) ? node1629 : 1'b1;
											assign node1629 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1632 = (inp[11]) ? 1'b0 : node1633;
											assign node1633 = (inp[14]) ? node1635 : 1'b1;
												assign node1635 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1639 = (inp[14]) ? 1'b0 : node1640;
										assign node1640 = (inp[2]) ? 1'b0 : node1641;
											assign node1641 = (inp[7]) ? node1643 : 1'b1;
												assign node1643 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1648 = (inp[7]) ? node1660 : node1649;
								assign node1649 = (inp[14]) ? node1655 : node1650;
									assign node1650 = (inp[6]) ? node1652 : 1'b1;
										assign node1652 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1655 = (inp[11]) ? 1'b0 : node1656;
										assign node1656 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1660 = (inp[0]) ? 1'b0 : node1661;
									assign node1661 = (inp[14]) ? 1'b0 : node1662;
										assign node1662 = (inp[12]) ? 1'b0 : node1663;
											assign node1663 = (inp[13]) ? node1665 : 1'b1;
												assign node1665 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1671 = (inp[1]) ? node1699 : node1672;
							assign node1672 = (inp[3]) ? node1688 : node1673;
								assign node1673 = (inp[11]) ? 1'b0 : node1674;
									assign node1674 = (inp[0]) ? node1680 : node1675;
										assign node1675 = (inp[13]) ? node1677 : 1'b1;
											assign node1677 = (inp[12]) ? 1'b1 : 1'b0;
										assign node1680 = (inp[14]) ? 1'b0 : node1681;
											assign node1681 = (inp[13]) ? node1683 : 1'b1;
												assign node1683 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1688 = (inp[7]) ? 1'b0 : node1689;
									assign node1689 = (inp[13]) ? 1'b0 : node1690;
										assign node1690 = (inp[12]) ? 1'b0 : node1691;
											assign node1691 = (inp[2]) ? node1693 : 1'b1;
												assign node1693 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1699 = (inp[14]) ? 1'b0 : node1700;
								assign node1700 = (inp[6]) ? 1'b0 : node1701;
									assign node1701 = (inp[7]) ? 1'b0 : node1702;
										assign node1702 = (inp[11]) ? 1'b0 : 1'b1;
					assign node1708 = (inp[0]) ? node1760 : node1709;
						assign node1709 = (inp[1]) ? node1749 : node1710;
							assign node1710 = (inp[7]) ? node1734 : node1711;
								assign node1711 = (inp[14]) ? node1723 : node1712;
									assign node1712 = (inp[3]) ? node1720 : node1713;
										assign node1713 = (inp[11]) ? node1715 : 1'b1;
											assign node1715 = (inp[2]) ? 1'b0 : node1716;
												assign node1716 = (inp[12]) ? 1'b1 : 1'b0;
										assign node1720 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1723 = (inp[13]) ? 1'b0 : node1724;
										assign node1724 = (inp[6]) ? node1728 : node1725;
											assign node1725 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1728 = (inp[10]) ? node1730 : 1'b0;
												assign node1730 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1734 = (inp[10]) ? 1'b0 : node1735;
									assign node1735 = (inp[11]) ? 1'b0 : node1736;
										assign node1736 = (inp[2]) ? node1742 : node1737;
											assign node1737 = (inp[3]) ? node1739 : 1'b1;
												assign node1739 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1742 = (inp[3]) ? 1'b0 : node1743;
												assign node1743 = (inp[14]) ? 1'b0 : 1'b1;
							assign node1749 = (inp[13]) ? 1'b0 : node1750;
								assign node1750 = (inp[10]) ? 1'b0 : node1751;
									assign node1751 = (inp[11]) ? 1'b0 : node1752;
										assign node1752 = (inp[3]) ? 1'b0 : node1753;
											assign node1753 = (inp[12]) ? 1'b0 : 1'b1;
						assign node1760 = (inp[3]) ? 1'b0 : node1761;
							assign node1761 = (inp[14]) ? 1'b0 : node1762;
								assign node1762 = (inp[2]) ? 1'b0 : node1763;
									assign node1763 = (inp[11]) ? 1'b0 : node1764;
										assign node1764 = (inp[13]) ? 1'b0 : 1'b1;

endmodule