module dtc_split125_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;

	assign outp = (inp[3]) ? node100 : node1;
		assign node1 = (inp[9]) ? node35 : node2;
			assign node2 = (inp[4]) ? node22 : node3;
				assign node3 = (inp[1]) ? node17 : node4;
					assign node4 = (inp[0]) ? node10 : node5;
						assign node5 = (inp[5]) ? 3'b000 : node6;
							assign node6 = (inp[6]) ? 3'b000 : 3'b001;
						assign node10 = (inp[6]) ? 3'b001 : node11;
							assign node11 = (inp[11]) ? node13 : 3'b000;
								assign node13 = (inp[2]) ? 3'b000 : 3'b001;
					assign node17 = (inp[6]) ? node19 : 3'b001;
						assign node19 = (inp[0]) ? 3'b001 : 3'b000;
				assign node22 = (inp[0]) ? node24 : 3'b000;
					assign node24 = (inp[5]) ? node30 : node25;
						assign node25 = (inp[1]) ? node27 : 3'b000;
							assign node27 = (inp[6]) ? 3'b000 : 3'b001;
						assign node30 = (inp[1]) ? 3'b000 : node31;
							assign node31 = (inp[6]) ? 3'b001 : 3'b000;
			assign node35 = (inp[6]) ? node75 : node36;
				assign node36 = (inp[4]) ? node58 : node37;
					assign node37 = (inp[7]) ? node49 : node38;
						assign node38 = (inp[0]) ? node44 : node39;
							assign node39 = (inp[5]) ? 3'b010 : node40;
								assign node40 = (inp[1]) ? 3'b110 : 3'b010;
							assign node44 = (inp[5]) ? node46 : 3'b001;
								assign node46 = (inp[1]) ? 3'b110 : 3'b001;
						assign node49 = (inp[5]) ? node51 : 3'b110;
							assign node51 = (inp[1]) ? node55 : node52;
								assign node52 = (inp[0]) ? 3'b001 : 3'b100;
								assign node55 = (inp[0]) ? 3'b110 : 3'b010;
					assign node58 = (inp[0]) ? node66 : node59;
						assign node59 = (inp[8]) ? 3'b000 : node60;
							assign node60 = (inp[11]) ? 3'b000 : node61;
								assign node61 = (inp[10]) ? 3'b100 : 3'b000;
						assign node66 = (inp[8]) ? node68 : 3'b100;
							assign node68 = (inp[11]) ? node70 : 3'b100;
								assign node70 = (inp[10]) ? node72 : 3'b100;
									assign node72 = (inp[7]) ? 3'b010 : 3'b100;
				assign node75 = (inp[0]) ? node77 : 3'b001;
					assign node77 = (inp[4]) ? node89 : node78;
						assign node78 = (inp[5]) ? node82 : node79;
							assign node79 = (inp[1]) ? 3'b111 : 3'b011;
							assign node82 = (inp[7]) ? node84 : 3'b011;
								assign node84 = (inp[1]) ? 3'b011 : node85;
									assign node85 = (inp[10]) ? 3'b111 : 3'b011;
						assign node89 = (inp[5]) ? node97 : node90;
							assign node90 = (inp[1]) ? 3'b101 : node91;
								assign node91 = (inp[2]) ? node93 : 3'b001;
									assign node93 = (inp[11]) ? 3'b101 : 3'b001;
							assign node97 = (inp[1]) ? 3'b001 : 3'b010;
		assign node100 = (inp[6]) ? node102 : 3'b000;
			assign node102 = (inp[0]) ? node114 : node103;
				assign node103 = (inp[9]) ? node111 : node104;
					assign node104 = (inp[4]) ? node106 : 3'b000;
						assign node106 = (inp[1]) ? node108 : 3'b010;
							assign node108 = (inp[10]) ? 3'b100 : 3'b010;
					assign node111 = (inp[4]) ? 3'b000 : 3'b100;
				assign node114 = (inp[4]) ? node118 : node115;
					assign node115 = (inp[9]) ? 3'b010 : 3'b001;
					assign node118 = (inp[9]) ? node128 : node119;
						assign node119 = (inp[10]) ? node125 : node120;
							assign node120 = (inp[8]) ? 3'b110 : node121;
								assign node121 = (inp[5]) ? 3'b110 : 3'b010;
							assign node125 = (inp[1]) ? 3'b110 : 3'b010;
						assign node128 = (inp[7]) ? node130 : 3'b000;
							assign node130 = (inp[10]) ? 3'b000 : node131;
								assign node131 = (inp[5]) ? node133 : 3'b100;
									assign node133 = (inp[8]) ? 3'b100 : 3'b000;

endmodule