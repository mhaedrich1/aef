module dtc_split66_bm72 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node952;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1077;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1143;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1176;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1243;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;
	wire [3-1:0] node1261;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1283;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1290;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1297;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1302;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1340;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1356;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1388;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1393;
	wire [3-1:0] node1396;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1442;
	wire [3-1:0] node1445;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1453;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1473;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1482;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1498;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1505;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1513;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;
	wire [3-1:0] node1521;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1546;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1553;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1562;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1574;
	wire [3-1:0] node1577;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;

	assign outp = (inp[3]) ? node874 : node1;
		assign node1 = (inp[6]) ? node459 : node2;
			assign node2 = (inp[9]) ? node246 : node3;
				assign node3 = (inp[0]) ? node125 : node4;
					assign node4 = (inp[4]) ? node66 : node5;
						assign node5 = (inp[8]) ? node37 : node6;
							assign node6 = (inp[5]) ? node22 : node7;
								assign node7 = (inp[7]) ? node15 : node8;
									assign node8 = (inp[11]) ? node12 : node9;
										assign node9 = (inp[1]) ? 3'b001 : 3'b001;
										assign node12 = (inp[1]) ? 3'b001 : 3'b001;
									assign node15 = (inp[11]) ? node19 : node16;
										assign node16 = (inp[1]) ? 3'b011 : 3'b011;
										assign node19 = (inp[2]) ? 3'b101 : 3'b011;
								assign node22 = (inp[7]) ? node30 : node23;
									assign node23 = (inp[1]) ? node27 : node24;
										assign node24 = (inp[10]) ? 3'b001 : 3'b101;
										assign node27 = (inp[10]) ? 3'b110 : 3'b001;
									assign node30 = (inp[11]) ? node34 : node31;
										assign node31 = (inp[2]) ? 3'b101 : 3'b101;
										assign node34 = (inp[1]) ? 3'b001 : 3'b001;
							assign node37 = (inp[7]) ? node51 : node38;
								assign node38 = (inp[5]) ? node46 : node39;
									assign node39 = (inp[1]) ? node43 : node40;
										assign node40 = (inp[2]) ? 3'b001 : 3'b011;
										assign node43 = (inp[10]) ? 3'b001 : 3'b101;
									assign node46 = (inp[10]) ? node48 : 3'b101;
										assign node48 = (inp[2]) ? 3'b110 : 3'b001;
								assign node51 = (inp[10]) ? node59 : node52;
									assign node52 = (inp[5]) ? node56 : node53;
										assign node53 = (inp[11]) ? 3'b111 : 3'b111;
										assign node56 = (inp[1]) ? 3'b011 : 3'b111;
									assign node59 = (inp[1]) ? node63 : node60;
										assign node60 = (inp[5]) ? 3'b011 : 3'b011;
										assign node63 = (inp[5]) ? 3'b101 : 3'b011;
						assign node66 = (inp[7]) ? node98 : node67;
							assign node67 = (inp[8]) ? node83 : node68;
								assign node68 = (inp[11]) ? node76 : node69;
									assign node69 = (inp[10]) ? node73 : node70;
										assign node70 = (inp[1]) ? 3'b010 : 3'b001;
										assign node73 = (inp[1]) ? 3'b010 : 3'b110;
									assign node76 = (inp[10]) ? node80 : node77;
										assign node77 = (inp[5]) ? 3'b010 : 3'b110;
										assign node80 = (inp[2]) ? 3'b010 : 3'b110;
								assign node83 = (inp[1]) ? node91 : node84;
									assign node84 = (inp[10]) ? node88 : node85;
										assign node85 = (inp[5]) ? 3'b001 : 3'b101;
										assign node88 = (inp[5]) ? 3'b110 : 3'b001;
									assign node91 = (inp[5]) ? node95 : node92;
										assign node92 = (inp[10]) ? 3'b110 : 3'b001;
										assign node95 = (inp[10]) ? 3'b010 : 3'b110;
							assign node98 = (inp[1]) ? node112 : node99;
								assign node99 = (inp[10]) ? node105 : node100;
									assign node100 = (inp[5]) ? 3'b101 : node101;
										assign node101 = (inp[8]) ? 3'b011 : 3'b101;
									assign node105 = (inp[8]) ? node109 : node106;
										assign node106 = (inp[5]) ? 3'b110 : 3'b001;
										assign node109 = (inp[5]) ? 3'b001 : 3'b101;
								assign node112 = (inp[10]) ? node120 : node113;
									assign node113 = (inp[2]) ? node117 : node114;
										assign node114 = (inp[8]) ? 3'b001 : 3'b001;
										assign node117 = (inp[5]) ? 3'b000 : 3'b001;
									assign node120 = (inp[2]) ? node122 : 3'b110;
										assign node122 = (inp[8]) ? 3'b110 : 3'b110;
					assign node125 = (inp[7]) ? node185 : node126;
						assign node126 = (inp[4]) ? node156 : node127;
							assign node127 = (inp[10]) ? node143 : node128;
								assign node128 = (inp[1]) ? node136 : node129;
									assign node129 = (inp[8]) ? node133 : node130;
										assign node130 = (inp[5]) ? 3'b010 : 3'b001;
										assign node133 = (inp[11]) ? 3'b001 : 3'b001;
									assign node136 = (inp[5]) ? node140 : node137;
										assign node137 = (inp[2]) ? 3'b110 : 3'b110;
										assign node140 = (inp[8]) ? 3'b110 : 3'b010;
								assign node143 = (inp[8]) ? node149 : node144;
									assign node144 = (inp[1]) ? 3'b100 : node145;
										assign node145 = (inp[5]) ? 3'b010 : 3'b110;
									assign node149 = (inp[1]) ? node153 : node150;
										assign node150 = (inp[2]) ? 3'b110 : 3'b000;
										assign node153 = (inp[11]) ? 3'b010 : 3'b010;
							assign node156 = (inp[10]) ? node170 : node157;
								assign node157 = (inp[1]) ? node165 : node158;
									assign node158 = (inp[11]) ? node162 : node159;
										assign node159 = (inp[2]) ? 3'b010 : 3'b110;
										assign node162 = (inp[5]) ? 3'b000 : 3'b010;
									assign node165 = (inp[5]) ? 3'b100 : node166;
										assign node166 = (inp[2]) ? 3'b100 : 3'b010;
								assign node170 = (inp[8]) ? node178 : node171;
									assign node171 = (inp[1]) ? node175 : node172;
										assign node172 = (inp[5]) ? 3'b000 : 3'b100;
										assign node175 = (inp[2]) ? 3'b000 : 3'b000;
									assign node178 = (inp[5]) ? node182 : node179;
										assign node179 = (inp[1]) ? 3'b100 : 3'b010;
										assign node182 = (inp[1]) ? 3'b000 : 3'b100;
						assign node185 = (inp[4]) ? node217 : node186;
							assign node186 = (inp[5]) ? node202 : node187;
								assign node187 = (inp[10]) ? node195 : node188;
									assign node188 = (inp[1]) ? node192 : node189;
										assign node189 = (inp[11]) ? 3'b101 : 3'b001;
										assign node192 = (inp[8]) ? 3'b101 : 3'b001;
									assign node195 = (inp[8]) ? node199 : node196;
										assign node196 = (inp[1]) ? 3'b110 : 3'b001;
										assign node199 = (inp[1]) ? 3'b001 : 3'b101;
								assign node202 = (inp[1]) ? node210 : node203;
									assign node203 = (inp[8]) ? node207 : node204;
										assign node204 = (inp[10]) ? 3'b110 : 3'b001;
										assign node207 = (inp[10]) ? 3'b001 : 3'b101;
									assign node210 = (inp[8]) ? node214 : node211;
										assign node211 = (inp[10]) ? 3'b010 : 3'b110;
										assign node214 = (inp[11]) ? 3'b110 : 3'b001;
							assign node217 = (inp[1]) ? node233 : node218;
								assign node218 = (inp[10]) ? node226 : node219;
									assign node219 = (inp[11]) ? node223 : node220;
										assign node220 = (inp[2]) ? 3'b001 : 3'b001;
										assign node223 = (inp[8]) ? 3'b000 : 3'b110;
									assign node226 = (inp[5]) ? node230 : node227;
										assign node227 = (inp[8]) ? 3'b000 : 3'b110;
										assign node230 = (inp[8]) ? 3'b110 : 3'b010;
								assign node233 = (inp[10]) ? node239 : node234;
									assign node234 = (inp[8]) ? node236 : 3'b010;
										assign node236 = (inp[5]) ? 3'b010 : 3'b110;
									assign node239 = (inp[11]) ? node243 : node240;
										assign node240 = (inp[2]) ? 3'b010 : 3'b110;
										assign node243 = (inp[2]) ? 3'b100 : 3'b010;
				assign node246 = (inp[0]) ? node368 : node247;
					assign node247 = (inp[7]) ? node307 : node248;
						assign node248 = (inp[4]) ? node280 : node249;
							assign node249 = (inp[8]) ? node265 : node250;
								assign node250 = (inp[11]) ? node258 : node251;
									assign node251 = (inp[1]) ? node255 : node252;
										assign node252 = (inp[10]) ? 3'b010 : 3'b110;
										assign node255 = (inp[10]) ? 3'b010 : 3'b010;
									assign node258 = (inp[1]) ? node262 : node259;
										assign node259 = (inp[5]) ? 3'b010 : 3'b010;
										assign node262 = (inp[10]) ? 3'b100 : 3'b010;
								assign node265 = (inp[5]) ? node273 : node266;
									assign node266 = (inp[10]) ? node270 : node267;
										assign node267 = (inp[11]) ? 3'b001 : 3'b001;
										assign node270 = (inp[1]) ? 3'b010 : 3'b110;
									assign node273 = (inp[1]) ? node277 : node274;
										assign node274 = (inp[10]) ? 3'b010 : 3'b110;
										assign node277 = (inp[10]) ? 3'b100 : 3'b010;
							assign node280 = (inp[1]) ? node294 : node281;
								assign node281 = (inp[8]) ? node289 : node282;
									assign node282 = (inp[11]) ? node286 : node283;
										assign node283 = (inp[10]) ? 3'b100 : 3'b010;
										assign node286 = (inp[10]) ? 3'b000 : 3'b100;
									assign node289 = (inp[11]) ? node291 : 3'b010;
										assign node291 = (inp[5]) ? 3'b100 : 3'b010;
								assign node294 = (inp[10]) ? node302 : node295;
									assign node295 = (inp[8]) ? node299 : node296;
										assign node296 = (inp[5]) ? 3'b000 : 3'b100;
										assign node299 = (inp[5]) ? 3'b100 : 3'b000;
									assign node302 = (inp[5]) ? 3'b000 : node303;
										assign node303 = (inp[2]) ? 3'b000 : 3'b100;
						assign node307 = (inp[4]) ? node339 : node308;
							assign node308 = (inp[10]) ? node324 : node309;
								assign node309 = (inp[1]) ? node317 : node310;
									assign node310 = (inp[2]) ? node314 : node311;
										assign node311 = (inp[5]) ? 3'b101 : 3'b101;
										assign node314 = (inp[5]) ? 3'b101 : 3'b001;
									assign node317 = (inp[11]) ? node321 : node318;
										assign node318 = (inp[2]) ? 3'b001 : 3'b001;
										assign node321 = (inp[5]) ? 3'b110 : 3'b001;
								assign node324 = (inp[5]) ? node332 : node325;
									assign node325 = (inp[2]) ? node329 : node326;
										assign node326 = (inp[8]) ? 3'b001 : 3'b000;
										assign node329 = (inp[11]) ? 3'b110 : 3'b101;
									assign node332 = (inp[8]) ? node336 : node333;
										assign node333 = (inp[1]) ? 3'b010 : 3'b110;
										assign node336 = (inp[11]) ? 3'b110 : 3'b001;
							assign node339 = (inp[2]) ? node353 : node340;
								assign node340 = (inp[1]) ? node348 : node341;
									assign node341 = (inp[8]) ? node345 : node342;
										assign node342 = (inp[11]) ? 3'b110 : 3'b010;
										assign node345 = (inp[10]) ? 3'b000 : 3'b001;
									assign node348 = (inp[10]) ? 3'b100 : node349;
										assign node349 = (inp[8]) ? 3'b110 : 3'b010;
								assign node353 = (inp[1]) ? node361 : node354;
									assign node354 = (inp[10]) ? node358 : node355;
										assign node355 = (inp[8]) ? 3'b000 : 3'b110;
										assign node358 = (inp[5]) ? 3'b010 : 3'b010;
									assign node361 = (inp[5]) ? node365 : node362;
										assign node362 = (inp[8]) ? 3'b010 : 3'b010;
										assign node365 = (inp[10]) ? 3'b000 : 3'b000;
					assign node368 = (inp[7]) ? node404 : node369;
						assign node369 = (inp[4]) ? node395 : node370;
							assign node370 = (inp[1]) ? node386 : node371;
								assign node371 = (inp[10]) ? node379 : node372;
									assign node372 = (inp[5]) ? node376 : node373;
										assign node373 = (inp[11]) ? 3'b010 : 3'b010;
										assign node376 = (inp[8]) ? 3'b010 : 3'b100;
									assign node379 = (inp[5]) ? node383 : node380;
										assign node380 = (inp[2]) ? 3'b100 : 3'b100;
										assign node383 = (inp[8]) ? 3'b100 : 3'b000;
								assign node386 = (inp[10]) ? 3'b000 : node387;
									assign node387 = (inp[5]) ? node391 : node388;
										assign node388 = (inp[11]) ? 3'b100 : 3'b100;
										assign node391 = (inp[8]) ? 3'b100 : 3'b000;
							assign node395 = (inp[10]) ? 3'b000 : node396;
								assign node396 = (inp[1]) ? 3'b000 : node397;
									assign node397 = (inp[5]) ? 3'b000 : node398;
										assign node398 = (inp[8]) ? 3'b100 : 3'b000;
						assign node404 = (inp[4]) ? node430 : node405;
							assign node405 = (inp[10]) ? node419 : node406;
								assign node406 = (inp[5]) ? node412 : node407;
									assign node407 = (inp[8]) ? node409 : 3'b110;
										assign node409 = (inp[1]) ? 3'b110 : 3'b001;
									assign node412 = (inp[8]) ? node416 : node413;
										assign node413 = (inp[1]) ? 3'b100 : 3'b010;
										assign node416 = (inp[1]) ? 3'b010 : 3'b110;
								assign node419 = (inp[5]) ? node425 : node420;
									assign node420 = (inp[2]) ? node422 : 3'b010;
										assign node422 = (inp[1]) ? 3'b100 : 3'b010;
									assign node425 = (inp[8]) ? node427 : 3'b100;
										assign node427 = (inp[1]) ? 3'b100 : 3'b010;
							assign node430 = (inp[10]) ? node446 : node431;
								assign node431 = (inp[1]) ? node439 : node432;
									assign node432 = (inp[8]) ? node436 : node433;
										assign node433 = (inp[11]) ? 3'b100 : 3'b010;
										assign node436 = (inp[11]) ? 3'b010 : 3'b010;
									assign node439 = (inp[5]) ? node443 : node440;
										assign node440 = (inp[11]) ? 3'b100 : 3'b100;
										assign node443 = (inp[8]) ? 3'b100 : 3'b000;
								assign node446 = (inp[1]) ? node454 : node447;
									assign node447 = (inp[5]) ? node451 : node448;
										assign node448 = (inp[11]) ? 3'b100 : 3'b100;
										assign node451 = (inp[8]) ? 3'b100 : 3'b000;
									assign node454 = (inp[5]) ? 3'b000 : node455;
										assign node455 = (inp[8]) ? 3'b000 : 3'b000;
			assign node459 = (inp[9]) ? node635 : node460;
				assign node460 = (inp[0]) ? node524 : node461;
					assign node461 = (inp[4]) ? node477 : node462;
						assign node462 = (inp[5]) ? node464 : 3'b111;
							assign node464 = (inp[7]) ? 3'b111 : node465;
								assign node465 = (inp[10]) ? node471 : node466;
									assign node466 = (inp[2]) ? node468 : 3'b111;
										assign node468 = (inp[1]) ? 3'b011 : 3'b111;
									assign node471 = (inp[1]) ? 3'b011 : node472;
										assign node472 = (inp[8]) ? 3'b111 : 3'b011;
						assign node477 = (inp[7]) ? node509 : node478;
							assign node478 = (inp[10]) ? node494 : node479;
								assign node479 = (inp[1]) ? node487 : node480;
									assign node480 = (inp[8]) ? node484 : node481;
										assign node481 = (inp[2]) ? 3'b011 : 3'b111;
										assign node484 = (inp[5]) ? 3'b111 : 3'b111;
									assign node487 = (inp[5]) ? node491 : node488;
										assign node488 = (inp[8]) ? 3'b111 : 3'b011;
										assign node491 = (inp[11]) ? 3'b101 : 3'b011;
								assign node494 = (inp[5]) ? node502 : node495;
									assign node495 = (inp[8]) ? node499 : node496;
										assign node496 = (inp[1]) ? 3'b101 : 3'b001;
										assign node499 = (inp[1]) ? 3'b011 : 3'b011;
									assign node502 = (inp[1]) ? node506 : node503;
										assign node503 = (inp[8]) ? 3'b001 : 3'b101;
										assign node506 = (inp[8]) ? 3'b101 : 3'b001;
							assign node509 = (inp[10]) ? node511 : 3'b111;
								assign node511 = (inp[8]) ? node519 : node512;
									assign node512 = (inp[11]) ? node516 : node513;
										assign node513 = (inp[5]) ? 3'b011 : 3'b111;
										assign node516 = (inp[2]) ? 3'b011 : 3'b011;
									assign node519 = (inp[1]) ? node521 : 3'b111;
										assign node521 = (inp[2]) ? 3'b011 : 3'b111;
					assign node524 = (inp[4]) ? node574 : node525;
						assign node525 = (inp[7]) ? node555 : node526;
							assign node526 = (inp[10]) ? node542 : node527;
								assign node527 = (inp[1]) ? node535 : node528;
									assign node528 = (inp[5]) ? node532 : node529;
										assign node529 = (inp[8]) ? 3'b111 : 3'b011;
										assign node532 = (inp[11]) ? 3'b011 : 3'b011;
									assign node535 = (inp[11]) ? node539 : node536;
										assign node536 = (inp[8]) ? 3'b011 : 3'b001;
										assign node539 = (inp[8]) ? 3'b001 : 3'b101;
								assign node542 = (inp[11]) ? node550 : node543;
									assign node543 = (inp[2]) ? node547 : node544;
										assign node544 = (inp[5]) ? 3'b001 : 3'b011;
										assign node547 = (inp[8]) ? 3'b101 : 3'b101;
									assign node550 = (inp[1]) ? node552 : 3'b101;
										assign node552 = (inp[5]) ? 3'b001 : 3'b101;
							assign node555 = (inp[10]) ? node563 : node556;
								assign node556 = (inp[2]) ? node558 : 3'b111;
									assign node558 = (inp[1]) ? node560 : 3'b111;
										assign node560 = (inp[11]) ? 3'b011 : 3'b111;
								assign node563 = (inp[1]) ? node569 : node564;
									assign node564 = (inp[11]) ? node566 : 3'b111;
										assign node566 = (inp[8]) ? 3'b111 : 3'b011;
									assign node569 = (inp[5]) ? 3'b011 : node570;
										assign node570 = (inp[8]) ? 3'b111 : 3'b011;
						assign node574 = (inp[7]) ? node606 : node575;
							assign node575 = (inp[1]) ? node591 : node576;
								assign node576 = (inp[11]) ? node584 : node577;
									assign node577 = (inp[10]) ? node581 : node578;
										assign node578 = (inp[5]) ? 3'b101 : 3'b001;
										assign node581 = (inp[5]) ? 3'b001 : 3'b101;
									assign node584 = (inp[10]) ? node588 : node585;
										assign node585 = (inp[5]) ? 3'b001 : 3'b101;
										assign node588 = (inp[5]) ? 3'b110 : 3'b001;
								assign node591 = (inp[5]) ? node599 : node592;
									assign node592 = (inp[10]) ? node596 : node593;
										assign node593 = (inp[11]) ? 3'b001 : 3'b101;
										assign node596 = (inp[11]) ? 3'b110 : 3'b001;
									assign node599 = (inp[2]) ? node603 : node600;
										assign node600 = (inp[11]) ? 3'b010 : 3'b001;
										assign node603 = (inp[10]) ? 3'b110 : 3'b110;
							assign node606 = (inp[10]) ? node622 : node607;
								assign node607 = (inp[1]) ? node615 : node608;
									assign node608 = (inp[5]) ? node612 : node609;
										assign node609 = (inp[8]) ? 3'b111 : 3'b011;
										assign node612 = (inp[2]) ? 3'b011 : 3'b011;
									assign node615 = (inp[5]) ? node619 : node616;
										assign node616 = (inp[8]) ? 3'b011 : 3'b101;
										assign node619 = (inp[11]) ? 3'b001 : 3'b101;
								assign node622 = (inp[1]) ? node628 : node623;
									assign node623 = (inp[5]) ? 3'b101 : node624;
										assign node624 = (inp[2]) ? 3'b101 : 3'b011;
									assign node628 = (inp[8]) ? node632 : node629;
										assign node629 = (inp[2]) ? 3'b000 : 3'b001;
										assign node632 = (inp[5]) ? 3'b001 : 3'b101;
				assign node635 = (inp[0]) ? node751 : node636;
					assign node636 = (inp[4]) ? node690 : node637;
						assign node637 = (inp[7]) ? node667 : node638;
							assign node638 = (inp[10]) ? node652 : node639;
								assign node639 = (inp[5]) ? node647 : node640;
									assign node640 = (inp[1]) ? node644 : node641;
										assign node641 = (inp[11]) ? 3'b011 : 3'b111;
										assign node644 = (inp[2]) ? 3'b001 : 3'b011;
									assign node647 = (inp[1]) ? 3'b101 : node648;
										assign node648 = (inp[8]) ? 3'b011 : 3'b101;
								assign node652 = (inp[5]) ? node660 : node653;
									assign node653 = (inp[1]) ? node657 : node654;
										assign node654 = (inp[2]) ? 3'b101 : 3'b001;
										assign node657 = (inp[8]) ? 3'b101 : 3'b001;
									assign node660 = (inp[8]) ? node664 : node661;
										assign node661 = (inp[2]) ? 3'b001 : 3'b001;
										assign node664 = (inp[1]) ? 3'b001 : 3'b001;
							assign node667 = (inp[10]) ? node677 : node668;
								assign node668 = (inp[5]) ? node670 : 3'b111;
									assign node670 = (inp[11]) ? node674 : node671;
										assign node671 = (inp[8]) ? 3'b111 : 3'b011;
										assign node674 = (inp[1]) ? 3'b011 : 3'b111;
								assign node677 = (inp[5]) ? node683 : node678;
									assign node678 = (inp[1]) ? 3'b011 : node679;
										assign node679 = (inp[11]) ? 3'b111 : 3'b111;
									assign node683 = (inp[8]) ? node687 : node684;
										assign node684 = (inp[1]) ? 3'b101 : 3'b001;
										assign node687 = (inp[1]) ? 3'b011 : 3'b111;
						assign node690 = (inp[7]) ? node722 : node691;
							assign node691 = (inp[10]) ? node707 : node692;
								assign node692 = (inp[1]) ? node700 : node693;
									assign node693 = (inp[11]) ? node697 : node694;
										assign node694 = (inp[5]) ? 3'b101 : 3'b101;
										assign node697 = (inp[2]) ? 3'b001 : 3'b101;
									assign node700 = (inp[5]) ? node704 : node701;
										assign node701 = (inp[8]) ? 3'b101 : 3'b001;
										assign node704 = (inp[11]) ? 3'b110 : 3'b001;
								assign node707 = (inp[8]) ? node715 : node708;
									assign node708 = (inp[1]) ? node712 : node709;
										assign node709 = (inp[5]) ? 3'b110 : 3'b001;
										assign node712 = (inp[5]) ? 3'b010 : 3'b110;
									assign node715 = (inp[5]) ? node719 : node716;
										assign node716 = (inp[1]) ? 3'b001 : 3'b001;
										assign node719 = (inp[2]) ? 3'b010 : 3'b001;
							assign node722 = (inp[10]) ? node738 : node723;
								assign node723 = (inp[1]) ? node731 : node724;
									assign node724 = (inp[2]) ? node728 : node725;
										assign node725 = (inp[5]) ? 3'b011 : 3'b111;
										assign node728 = (inp[11]) ? 3'b011 : 3'b011;
									assign node731 = (inp[8]) ? node735 : node732;
										assign node732 = (inp[2]) ? 3'b101 : 3'b101;
										assign node735 = (inp[5]) ? 3'b101 : 3'b011;
								assign node738 = (inp[5]) ? node746 : node739;
									assign node739 = (inp[1]) ? node743 : node740;
										assign node740 = (inp[11]) ? 3'b101 : 3'b011;
										assign node743 = (inp[8]) ? 3'b101 : 3'b001;
									assign node746 = (inp[2]) ? 3'b001 : node747;
										assign node747 = (inp[11]) ? 3'b001 : 3'b101;
					assign node751 = (inp[4]) ? node811 : node752;
						assign node752 = (inp[7]) ? node782 : node753;
							assign node753 = (inp[10]) ? node769 : node754;
								assign node754 = (inp[5]) ? node762 : node755;
									assign node755 = (inp[1]) ? node759 : node756;
										assign node756 = (inp[8]) ? 3'b101 : 3'b001;
										assign node759 = (inp[11]) ? 3'b001 : 3'b001;
									assign node762 = (inp[1]) ? node766 : node763;
										assign node763 = (inp[8]) ? 3'b001 : 3'b000;
										assign node766 = (inp[2]) ? 3'b010 : 3'b110;
								assign node769 = (inp[8]) ? node775 : node770;
									assign node770 = (inp[1]) ? node772 : 3'b110;
										assign node772 = (inp[5]) ? 3'b010 : 3'b110;
									assign node775 = (inp[1]) ? node779 : node776;
										assign node776 = (inp[2]) ? 3'b001 : 3'b001;
										assign node779 = (inp[5]) ? 3'b110 : 3'b110;
							assign node782 = (inp[10]) ? node798 : node783;
								assign node783 = (inp[8]) ? node791 : node784;
									assign node784 = (inp[11]) ? node788 : node785;
										assign node785 = (inp[1]) ? 3'b101 : 3'b011;
										assign node788 = (inp[1]) ? 3'b001 : 3'b101;
									assign node791 = (inp[1]) ? node795 : node792;
										assign node792 = (inp[2]) ? 3'b011 : 3'b111;
										assign node795 = (inp[5]) ? 3'b101 : 3'b011;
								assign node798 = (inp[1]) ? node804 : node799;
									assign node799 = (inp[2]) ? node801 : 3'b101;
										assign node801 = (inp[11]) ? 3'b001 : 3'b101;
									assign node804 = (inp[5]) ? node808 : node805;
										assign node805 = (inp[8]) ? 3'b101 : 3'b001;
										assign node808 = (inp[2]) ? 3'b110 : 3'b000;
						assign node811 = (inp[7]) ? node843 : node812;
							assign node812 = (inp[10]) ? node828 : node813;
								assign node813 = (inp[5]) ? node821 : node814;
									assign node814 = (inp[1]) ? node818 : node815;
										assign node815 = (inp[8]) ? 3'b000 : 3'b110;
										assign node818 = (inp[2]) ? 3'b010 : 3'b110;
									assign node821 = (inp[2]) ? node825 : node822;
										assign node822 = (inp[8]) ? 3'b110 : 3'b010;
										assign node825 = (inp[8]) ? 3'b110 : 3'b100;
								assign node828 = (inp[11]) ? node836 : node829;
									assign node829 = (inp[8]) ? node833 : node830;
										assign node830 = (inp[1]) ? 3'b000 : 3'b010;
										assign node833 = (inp[1]) ? 3'b010 : 3'b110;
									assign node836 = (inp[1]) ? node840 : node837;
										assign node837 = (inp[5]) ? 3'b100 : 3'b010;
										assign node840 = (inp[2]) ? 3'b100 : 3'b000;
							assign node843 = (inp[10]) ? node859 : node844;
								assign node844 = (inp[11]) ? node852 : node845;
									assign node845 = (inp[1]) ? node849 : node846;
										assign node846 = (inp[8]) ? 3'b001 : 3'b001;
										assign node849 = (inp[8]) ? 3'b001 : 3'b000;
									assign node852 = (inp[1]) ? node856 : node853;
										assign node853 = (inp[5]) ? 3'b110 : 3'b001;
										assign node856 = (inp[8]) ? 3'b110 : 3'b010;
								assign node859 = (inp[1]) ? node867 : node860;
									assign node860 = (inp[5]) ? node864 : node861;
										assign node861 = (inp[8]) ? 3'b001 : 3'b110;
										assign node864 = (inp[2]) ? 3'b010 : 3'b110;
									assign node867 = (inp[5]) ? node871 : node868;
										assign node868 = (inp[11]) ? 3'b110 : 3'b110;
										assign node871 = (inp[2]) ? 3'b010 : 3'b010;
		assign node874 = (inp[6]) ? node1130 : node875;
			assign node875 = (inp[9]) ? node1047 : node876;
				assign node876 = (inp[0]) ? node986 : node877;
					assign node877 = (inp[4]) ? node937 : node878;
						assign node878 = (inp[7]) ? node908 : node879;
							assign node879 = (inp[10]) ? node893 : node880;
								assign node880 = (inp[5]) ? node888 : node881;
									assign node881 = (inp[1]) ? node885 : node882;
										assign node882 = (inp[2]) ? 3'b010 : 3'b110;
										assign node885 = (inp[8]) ? 3'b010 : 3'b010;
									assign node888 = (inp[8]) ? 3'b010 : node889;
										assign node889 = (inp[1]) ? 3'b100 : 3'b010;
								assign node893 = (inp[8]) ? node901 : node894;
									assign node894 = (inp[5]) ? node898 : node895;
										assign node895 = (inp[11]) ? 3'b100 : 3'b100;
										assign node898 = (inp[11]) ? 3'b000 : 3'b000;
									assign node901 = (inp[5]) ? node905 : node902;
										assign node902 = (inp[1]) ? 3'b000 : 3'b010;
										assign node905 = (inp[2]) ? 3'b000 : 3'b100;
							assign node908 = (inp[1]) ? node922 : node909;
								assign node909 = (inp[5]) ? node917 : node910;
									assign node910 = (inp[2]) ? node914 : node911;
										assign node911 = (inp[8]) ? 3'b001 : 3'b001;
										assign node914 = (inp[8]) ? 3'b001 : 3'b010;
									assign node917 = (inp[8]) ? node919 : 3'b110;
										assign node919 = (inp[10]) ? 3'b110 : 3'b001;
								assign node922 = (inp[5]) ? node930 : node923;
									assign node923 = (inp[10]) ? node927 : node924;
										assign node924 = (inp[2]) ? 3'b010 : 3'b001;
										assign node927 = (inp[8]) ? 3'b110 : 3'b010;
									assign node930 = (inp[10]) ? node934 : node931;
										assign node931 = (inp[2]) ? 3'b010 : 3'b110;
										assign node934 = (inp[11]) ? 3'b100 : 3'b010;
						assign node937 = (inp[7]) ? node959 : node938;
							assign node938 = (inp[2]) ? node952 : node939;
								assign node939 = (inp[5]) ? node947 : node940;
									assign node940 = (inp[8]) ? node944 : node941;
										assign node941 = (inp[11]) ? 3'b000 : 3'b100;
										assign node944 = (inp[1]) ? 3'b100 : 3'b000;
									assign node947 = (inp[10]) ? 3'b000 : node948;
										assign node948 = (inp[11]) ? 3'b000 : 3'b100;
								assign node952 = (inp[8]) ? node954 : 3'b000;
									assign node954 = (inp[5]) ? 3'b000 : node955;
										assign node955 = (inp[1]) ? 3'b000 : 3'b010;
							assign node959 = (inp[10]) ? node971 : node960;
								assign node960 = (inp[8]) ? node966 : node961;
									assign node961 = (inp[1]) ? node963 : 3'b010;
										assign node963 = (inp[5]) ? 3'b100 : 3'b000;
									assign node966 = (inp[5]) ? 3'b010 : node967;
										assign node967 = (inp[1]) ? 3'b010 : 3'b110;
								assign node971 = (inp[5]) ? node979 : node972;
									assign node972 = (inp[1]) ? node976 : node973;
										assign node973 = (inp[8]) ? 3'b010 : 3'b000;
										assign node976 = (inp[2]) ? 3'b100 : 3'b000;
									assign node979 = (inp[1]) ? node983 : node980;
										assign node980 = (inp[2]) ? 3'b100 : 3'b100;
										assign node983 = (inp[8]) ? 3'b100 : 3'b000;
					assign node986 = (inp[4]) ? node1034 : node987;
						assign node987 = (inp[7]) ? node1003 : node988;
							assign node988 = (inp[10]) ? 3'b000 : node989;
								assign node989 = (inp[1]) ? node997 : node990;
									assign node990 = (inp[5]) ? node994 : node991;
										assign node991 = (inp[2]) ? 3'b100 : 3'b100;
										assign node994 = (inp[11]) ? 3'b000 : 3'b000;
									assign node997 = (inp[11]) ? 3'b000 : node998;
										assign node998 = (inp[5]) ? 3'b000 : 3'b100;
							assign node1003 = (inp[1]) ? node1019 : node1004;
								assign node1004 = (inp[8]) ? node1012 : node1005;
									assign node1005 = (inp[11]) ? node1009 : node1006;
										assign node1006 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1009 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1012 = (inp[11]) ? node1016 : node1013;
										assign node1013 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1016 = (inp[5]) ? 3'b100 : 3'b010;
								assign node1019 = (inp[5]) ? node1027 : node1020;
									assign node1020 = (inp[10]) ? node1024 : node1021;
										assign node1021 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1024 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1027 = (inp[8]) ? node1031 : node1028;
										assign node1028 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1031 = (inp[10]) ? 3'b000 : 3'b100;
						assign node1034 = (inp[10]) ? 3'b000 : node1035;
							assign node1035 = (inp[1]) ? 3'b000 : node1036;
								assign node1036 = (inp[7]) ? node1038 : 3'b000;
									assign node1038 = (inp[5]) ? node1042 : node1039;
										assign node1039 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1042 = (inp[2]) ? 3'b000 : 3'b000;
				assign node1047 = (inp[0]) ? node1115 : node1048;
					assign node1048 = (inp[4]) ? node1098 : node1049;
						assign node1049 = (inp[7]) ? node1071 : node1050;
							assign node1050 = (inp[10]) ? node1064 : node1051;
								assign node1051 = (inp[5]) ? node1059 : node1052;
									assign node1052 = (inp[2]) ? node1056 : node1053;
										assign node1053 = (inp[1]) ? 3'b100 : 3'b100;
										assign node1056 = (inp[1]) ? 3'b000 : 3'b000;
									assign node1059 = (inp[11]) ? 3'b000 : node1060;
										assign node1060 = (inp[2]) ? 3'b000 : 3'b000;
								assign node1064 = (inp[8]) ? node1066 : 3'b000;
									assign node1066 = (inp[1]) ? 3'b000 : node1067;
										assign node1067 = (inp[11]) ? 3'b000 : 3'b000;
							assign node1071 = (inp[10]) ? node1085 : node1072;
								assign node1072 = (inp[1]) ? node1080 : node1073;
									assign node1073 = (inp[2]) ? node1077 : node1074;
										assign node1074 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1077 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1080 = (inp[2]) ? node1082 : 3'b100;
										assign node1082 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1085 = (inp[8]) ? node1091 : node1086;
									assign node1086 = (inp[1]) ? 3'b000 : node1087;
										assign node1087 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1091 = (inp[11]) ? node1095 : node1092;
										assign node1092 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1095 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1098 = (inp[7]) ? node1100 : 3'b000;
							assign node1100 = (inp[8]) ? node1102 : 3'b000;
								assign node1102 = (inp[1]) ? node1110 : node1103;
									assign node1103 = (inp[10]) ? node1107 : node1104;
										assign node1104 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1107 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1110 = (inp[11]) ? 3'b000 : node1111;
										assign node1111 = (inp[10]) ? 3'b000 : 3'b000;
					assign node1115 = (inp[4]) ? 3'b000 : node1116;
						assign node1116 = (inp[7]) ? node1118 : 3'b000;
							assign node1118 = (inp[10]) ? 3'b000 : node1119;
								assign node1119 = (inp[1]) ? 3'b000 : node1120;
									assign node1120 = (inp[11]) ? node1124 : node1121;
										assign node1121 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1124 = (inp[8]) ? 3'b000 : 3'b000;
			assign node1130 = (inp[9]) ? node1374 : node1131;
				assign node1131 = (inp[0]) ? node1253 : node1132;
					assign node1132 = (inp[7]) ? node1194 : node1133;
						assign node1133 = (inp[4]) ? node1163 : node1134;
							assign node1134 = (inp[1]) ? node1148 : node1135;
								assign node1135 = (inp[2]) ? node1143 : node1136;
									assign node1136 = (inp[8]) ? node1140 : node1137;
										assign node1137 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1140 = (inp[11]) ? 3'b101 : 3'b011;
									assign node1143 = (inp[5]) ? node1145 : 3'b101;
										assign node1145 = (inp[10]) ? 3'b000 : 3'b101;
								assign node1148 = (inp[10]) ? node1156 : node1149;
									assign node1149 = (inp[2]) ? node1153 : node1150;
										assign node1150 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1153 = (inp[5]) ? 3'b001 : 3'b001;
									assign node1156 = (inp[2]) ? node1160 : node1157;
										assign node1157 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1160 = (inp[5]) ? 3'b010 : 3'b110;
							assign node1163 = (inp[5]) ? node1179 : node1164;
								assign node1164 = (inp[1]) ? node1172 : node1165;
									assign node1165 = (inp[8]) ? node1169 : node1166;
										assign node1166 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1169 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1172 = (inp[2]) ? node1176 : node1173;
										assign node1173 = (inp[10]) ? 3'b110 : 3'b001;
										assign node1176 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1179 = (inp[10]) ? node1187 : node1180;
									assign node1180 = (inp[2]) ? node1184 : node1181;
										assign node1181 = (inp[1]) ? 3'b110 : 3'b000;
										assign node1184 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1187 = (inp[1]) ? node1191 : node1188;
										assign node1188 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1191 = (inp[8]) ? 3'b010 : 3'b100;
						assign node1194 = (inp[4]) ? node1222 : node1195;
							assign node1195 = (inp[1]) ? node1209 : node1196;
								assign node1196 = (inp[10]) ? node1202 : node1197;
									assign node1197 = (inp[8]) ? 3'b111 : node1198;
										assign node1198 = (inp[2]) ? 3'b011 : 3'b011;
									assign node1202 = (inp[8]) ? node1206 : node1203;
										assign node1203 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1206 = (inp[5]) ? 3'b011 : 3'b011;
								assign node1209 = (inp[11]) ? node1217 : node1210;
									assign node1210 = (inp[8]) ? node1214 : node1211;
										assign node1211 = (inp[10]) ? 3'b101 : 3'b001;
										assign node1214 = (inp[10]) ? 3'b001 : 3'b011;
									assign node1217 = (inp[10]) ? node1219 : 3'b101;
										assign node1219 = (inp[8]) ? 3'b101 : 3'b001;
							assign node1222 = (inp[10]) ? node1238 : node1223;
								assign node1223 = (inp[11]) ? node1231 : node1224;
									assign node1224 = (inp[1]) ? node1228 : node1225;
										assign node1225 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1228 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1231 = (inp[1]) ? node1235 : node1232;
										assign node1232 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1235 = (inp[5]) ? 3'b001 : 3'b001;
								assign node1238 = (inp[1]) ? node1246 : node1239;
									assign node1239 = (inp[8]) ? node1243 : node1240;
										assign node1240 = (inp[11]) ? 3'b000 : 3'b001;
										assign node1243 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1246 = (inp[8]) ? node1250 : node1247;
										assign node1247 = (inp[2]) ? 3'b110 : 3'b000;
										assign node1250 = (inp[5]) ? 3'b110 : 3'b001;
					assign node1253 = (inp[4]) ? node1313 : node1254;
						assign node1254 = (inp[7]) ? node1286 : node1255;
							assign node1255 = (inp[2]) ? node1271 : node1256;
								assign node1256 = (inp[11]) ? node1264 : node1257;
									assign node1257 = (inp[5]) ? node1261 : node1258;
										assign node1258 = (inp[1]) ? 3'b000 : 3'b001;
										assign node1261 = (inp[10]) ? 3'b010 : 3'b000;
									assign node1264 = (inp[10]) ? node1268 : node1265;
										assign node1265 = (inp[1]) ? 3'b110 : 3'b000;
										assign node1268 = (inp[5]) ? 3'b010 : 3'b010;
								assign node1271 = (inp[10]) ? node1279 : node1272;
									assign node1272 = (inp[5]) ? node1276 : node1273;
										assign node1273 = (inp[8]) ? 3'b110 : 3'b110;
										assign node1276 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1279 = (inp[11]) ? node1283 : node1280;
										assign node1280 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1283 = (inp[1]) ? 3'b000 : 3'b010;
							assign node1286 = (inp[5]) ? node1300 : node1287;
								assign node1287 = (inp[8]) ? node1293 : node1288;
									assign node1288 = (inp[11]) ? node1290 : 3'b001;
										assign node1290 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1293 = (inp[10]) ? node1297 : node1294;
										assign node1294 = (inp[1]) ? 3'b101 : 3'b011;
										assign node1297 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1300 = (inp[2]) ? node1308 : node1301;
									assign node1301 = (inp[1]) ? node1305 : node1302;
										assign node1302 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1305 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1308 = (inp[10]) ? 3'b110 : node1309;
										assign node1309 = (inp[1]) ? 3'b110 : 3'b001;
						assign node1313 = (inp[7]) ? node1343 : node1314;
							assign node1314 = (inp[10]) ? node1328 : node1315;
								assign node1315 = (inp[1]) ? node1321 : node1316;
									assign node1316 = (inp[8]) ? 3'b010 : node1317;
										assign node1317 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1321 = (inp[5]) ? node1325 : node1322;
										assign node1322 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1325 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1328 = (inp[8]) ? node1336 : node1329;
									assign node1329 = (inp[5]) ? node1333 : node1330;
										assign node1330 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1333 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1336 = (inp[1]) ? node1340 : node1337;
										assign node1337 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1340 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1343 = (inp[11]) ? node1359 : node1344;
								assign node1344 = (inp[8]) ? node1352 : node1345;
									assign node1345 = (inp[5]) ? node1349 : node1346;
										assign node1346 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1349 = (inp[10]) ? 3'b100 : 3'b010;
									assign node1352 = (inp[1]) ? node1356 : node1353;
										assign node1353 = (inp[2]) ? 3'b010 : 3'b001;
										assign node1356 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1359 = (inp[2]) ? node1367 : node1360;
									assign node1360 = (inp[10]) ? node1364 : node1361;
										assign node1361 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1364 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1367 = (inp[10]) ? node1371 : node1368;
										assign node1368 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1371 = (inp[1]) ? 3'b100 : 3'b110;
				assign node1374 = (inp[0]) ? node1492 : node1375;
					assign node1375 = (inp[7]) ? node1435 : node1376;
						assign node1376 = (inp[4]) ? node1406 : node1377;
							assign node1377 = (inp[1]) ? node1391 : node1378;
								assign node1378 = (inp[11]) ? node1384 : node1379;
									assign node1379 = (inp[8]) ? 3'b110 : node1380;
										assign node1380 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1384 = (inp[10]) ? node1388 : node1385;
										assign node1385 = (inp[5]) ? 3'b110 : 3'b000;
										assign node1388 = (inp[5]) ? 3'b010 : 3'b010;
								assign node1391 = (inp[10]) ? node1399 : node1392;
									assign node1392 = (inp[11]) ? node1396 : node1393;
										assign node1393 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1396 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1399 = (inp[8]) ? node1403 : node1400;
										assign node1400 = (inp[2]) ? 3'b100 : 3'b100;
										assign node1403 = (inp[5]) ? 3'b100 : 3'b010;
							assign node1406 = (inp[10]) ? node1422 : node1407;
								assign node1407 = (inp[5]) ? node1415 : node1408;
									assign node1408 = (inp[1]) ? node1412 : node1409;
										assign node1409 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1412 = (inp[8]) ? 3'b010 : 3'b100;
									assign node1415 = (inp[2]) ? node1419 : node1416;
										assign node1416 = (inp[1]) ? 3'b000 : 3'b010;
										assign node1419 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1422 = (inp[5]) ? node1430 : node1423;
									assign node1423 = (inp[8]) ? node1427 : node1424;
										assign node1424 = (inp[1]) ? 3'b000 : 3'b100;
										assign node1427 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1430 = (inp[11]) ? 3'b000 : node1431;
										assign node1431 = (inp[1]) ? 3'b000 : 3'b100;
						assign node1435 = (inp[4]) ? node1463 : node1436;
							assign node1436 = (inp[5]) ? node1450 : node1437;
								assign node1437 = (inp[10]) ? node1445 : node1438;
									assign node1438 = (inp[1]) ? node1442 : node1439;
										assign node1439 = (inp[8]) ? 3'b101 : 3'b101;
										assign node1442 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1445 = (inp[1]) ? node1447 : 3'b001;
										assign node1447 = (inp[8]) ? 3'b001 : 3'b010;
								assign node1450 = (inp[10]) ? node1456 : node1451;
									assign node1451 = (inp[2]) ? node1453 : 3'b001;
										assign node1453 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1456 = (inp[1]) ? node1460 : node1457;
										assign node1457 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1460 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1463 = (inp[10]) ? node1477 : node1464;
								assign node1464 = (inp[1]) ? node1472 : node1465;
									assign node1465 = (inp[5]) ? node1469 : node1466;
										assign node1466 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1469 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1472 = (inp[5]) ? 3'b010 : node1473;
										assign node1473 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1477 = (inp[1]) ? node1485 : node1478;
									assign node1478 = (inp[2]) ? node1482 : node1479;
										assign node1479 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1482 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1485 = (inp[8]) ? node1489 : node1486;
										assign node1486 = (inp[5]) ? 3'b100 : 3'b100;
										assign node1489 = (inp[5]) ? 3'b100 : 3'b010;
					assign node1492 = (inp[7]) ? node1526 : node1493;
						assign node1493 = (inp[4]) ? node1517 : node1494;
							assign node1494 = (inp[10]) ? node1508 : node1495;
								assign node1495 = (inp[8]) ? node1501 : node1496;
									assign node1496 = (inp[2]) ? node1498 : 3'b100;
										assign node1498 = (inp[1]) ? 3'b000 : 3'b000;
									assign node1501 = (inp[5]) ? node1505 : node1502;
										assign node1502 = (inp[11]) ? 3'b010 : 3'b000;
										assign node1505 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1508 = (inp[1]) ? 3'b000 : node1509;
									assign node1509 = (inp[11]) ? node1513 : node1510;
										assign node1510 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1513 = (inp[5]) ? 3'b000 : 3'b100;
							assign node1517 = (inp[10]) ? 3'b000 : node1518;
								assign node1518 = (inp[8]) ? node1520 : 3'b000;
									assign node1520 = (inp[2]) ? 3'b000 : node1521;
										assign node1521 = (inp[1]) ? 3'b000 : 3'b100;
						assign node1526 = (inp[4]) ? node1556 : node1527;
							assign node1527 = (inp[10]) ? node1541 : node1528;
								assign node1528 = (inp[11]) ? node1536 : node1529;
									assign node1529 = (inp[8]) ? node1533 : node1530;
										assign node1530 = (inp[5]) ? 3'b000 : 3'b110;
										assign node1533 = (inp[1]) ? 3'b010 : 3'b001;
									assign node1536 = (inp[2]) ? 3'b010 : node1537;
										assign node1537 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1541 = (inp[8]) ? node1549 : node1542;
									assign node1542 = (inp[11]) ? node1546 : node1543;
										assign node1543 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1546 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1549 = (inp[5]) ? node1553 : node1550;
										assign node1550 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1553 = (inp[2]) ? 3'b100 : 3'b010;
							assign node1556 = (inp[10]) ? node1572 : node1557;
								assign node1557 = (inp[11]) ? node1565 : node1558;
									assign node1558 = (inp[2]) ? node1562 : node1559;
										assign node1559 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1562 = (inp[5]) ? 3'b100 : 3'b000;
									assign node1565 = (inp[1]) ? node1569 : node1566;
										assign node1566 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1569 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1572 = (inp[1]) ? node1580 : node1573;
									assign node1573 = (inp[11]) ? node1577 : node1574;
										assign node1574 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1577 = (inp[5]) ? 3'b000 : 3'b000;
									assign node1580 = (inp[2]) ? 3'b000 : node1581;
										assign node1581 = (inp[8]) ? 3'b100 : 3'b000;

endmodule