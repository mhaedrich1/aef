module dtc_split66_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node6;
	wire [2-1:0] node10;
	wire [2-1:0] node11;
	wire [2-1:0] node12;
	wire [2-1:0] node16;
	wire [2-1:0] node17;
	wire [2-1:0] node21;
	wire [2-1:0] node22;
	wire [2-1:0] node25;
	wire [2-1:0] node27;
	wire [2-1:0] node30;
	wire [2-1:0] node31;
	wire [2-1:0] node32;
	wire [2-1:0] node34;
	wire [2-1:0] node37;
	wire [2-1:0] node39;
	wire [2-1:0] node42;
	wire [2-1:0] node43;
	wire [2-1:0] node45;
	wire [2-1:0] node48;
	wire [2-1:0] node50;
	wire [2-1:0] node53;
	wire [2-1:0] node54;
	wire [2-1:0] node55;
	wire [2-1:0] node56;
	wire [2-1:0] node58;
	wire [2-1:0] node61;
	wire [2-1:0] node62;
	wire [2-1:0] node64;
	wire [2-1:0] node67;
	wire [2-1:0] node69;
	wire [2-1:0] node72;
	wire [2-1:0] node73;
	wire [2-1:0] node77;
	wire [2-1:0] node78;
	wire [2-1:0] node79;
	wire [2-1:0] node81;
	wire [2-1:0] node82;
	wire [2-1:0] node86;
	wire [2-1:0] node87;
	wire [2-1:0] node90;
	wire [2-1:0] node93;
	wire [2-1:0] node94;
	wire [2-1:0] node95;
	wire [2-1:0] node99;
	wire [2-1:0] node100;
	wire [2-1:0] node101;
	wire [2-1:0] node104;
	wire [2-1:0] node107;
	wire [2-1:0] node109;
	wire [2-1:0] node112;
	wire [2-1:0] node113;
	wire [2-1:0] node114;
	wire [2-1:0] node115;
	wire [2-1:0] node116;
	wire [2-1:0] node118;
	wire [2-1:0] node121;
	wire [2-1:0] node123;
	wire [2-1:0] node124;
	wire [2-1:0] node127;
	wire [2-1:0] node130;
	wire [2-1:0] node131;
	wire [2-1:0] node132;
	wire [2-1:0] node133;
	wire [2-1:0] node136;
	wire [2-1:0] node140;
	wire [2-1:0] node142;
	wire [2-1:0] node143;
	wire [2-1:0] node146;
	wire [2-1:0] node149;
	wire [2-1:0] node150;
	wire [2-1:0] node151;
	wire [2-1:0] node152;
	wire [2-1:0] node155;
	wire [2-1:0] node156;
	wire [2-1:0] node160;
	wire [2-1:0] node161;
	wire [2-1:0] node164;
	wire [2-1:0] node165;
	wire [2-1:0] node169;
	wire [2-1:0] node170;
	wire [2-1:0] node172;
	wire [2-1:0] node173;
	wire [2-1:0] node176;
	wire [2-1:0] node179;
	wire [2-1:0] node180;
	wire [2-1:0] node183;
	wire [2-1:0] node186;
	wire [2-1:0] node187;
	wire [2-1:0] node188;
	wire [2-1:0] node189;
	wire [2-1:0] node190;
	wire [2-1:0] node193;
	wire [2-1:0] node194;
	wire [2-1:0] node199;
	wire [2-1:0] node200;
	wire [2-1:0] node202;
	wire [2-1:0] node206;
	wire [2-1:0] node207;
	wire [2-1:0] node208;
	wire [2-1:0] node209;
	wire [2-1:0] node212;
	wire [2-1:0] node215;
	wire [2-1:0] node216;
	wire [2-1:0] node217;
	wire [2-1:0] node220;
	wire [2-1:0] node224;
	wire [2-1:0] node225;
	wire [2-1:0] node227;
	wire [2-1:0] node230;
	wire [2-1:0] node231;
	wire [2-1:0] node234;

	assign outp = (inp[0]) ? node112 : node1;
		assign node1 = (inp[7]) ? node53 : node2;
			assign node2 = (inp[2]) ? node30 : node3;
				assign node3 = (inp[6]) ? node21 : node4;
					assign node4 = (inp[4]) ? node10 : node5;
						assign node5 = (inp[1]) ? 2'b01 : node6;
							assign node6 = (inp[5]) ? 2'b01 : 2'b11;
						assign node10 = (inp[1]) ? node16 : node11;
							assign node11 = (inp[3]) ? 2'b01 : node12;
								assign node12 = (inp[5]) ? 2'b01 : 2'b11;
							assign node16 = (inp[3]) ? 2'b11 : node17;
								assign node17 = (inp[5]) ? 2'b11 : 2'b01;
					assign node21 = (inp[5]) ? node25 : node22;
						assign node22 = (inp[1]) ? 2'b00 : 2'b10;
						assign node25 = (inp[1]) ? node27 : 2'b00;
							assign node27 = (inp[4]) ? 2'b00 : 2'b10;
				assign node30 = (inp[1]) ? node42 : node31;
					assign node31 = (inp[5]) ? node37 : node32;
						assign node32 = (inp[4]) ? node34 : 2'b10;
							assign node34 = (inp[3]) ? 2'b00 : 2'b10;
						assign node37 = (inp[3]) ? node39 : 2'b00;
							assign node39 = (inp[4]) ? 2'b10 : 2'b00;
					assign node42 = (inp[5]) ? node48 : node43;
						assign node43 = (inp[3]) ? node45 : 2'b00;
							assign node45 = (inp[6]) ? 2'b00 : 2'b10;
						assign node48 = (inp[3]) ? node50 : 2'b10;
							assign node50 = (inp[4]) ? 2'b00 : 2'b10;
			assign node53 = (inp[2]) ? node77 : node54;
				assign node54 = (inp[6]) ? node72 : node55;
					assign node55 = (inp[4]) ? node61 : node56;
						assign node56 = (inp[5]) ? node58 : 2'b10;
							assign node58 = (inp[1]) ? 2'b10 : 2'b00;
						assign node61 = (inp[1]) ? node67 : node62;
							assign node62 = (inp[3]) ? node64 : 2'b10;
								assign node64 = (inp[5]) ? 2'b10 : 2'b00;
							assign node67 = (inp[3]) ? node69 : 2'b00;
								assign node69 = (inp[5]) ? 2'b00 : 2'b10;
					assign node72 = (inp[1]) ? 2'b01 : node73;
						assign node73 = (inp[4]) ? 2'b01 : 2'b11;
				assign node77 = (inp[4]) ? node93 : node78;
					assign node78 = (inp[3]) ? node86 : node79;
						assign node79 = (inp[6]) ? node81 : 2'b01;
							assign node81 = (inp[1]) ? 2'b01 : node82;
								assign node82 = (inp[5]) ? 2'b01 : 2'b11;
						assign node86 = (inp[1]) ? node90 : node87;
							assign node87 = (inp[5]) ? 2'b11 : 2'b01;
							assign node90 = (inp[5]) ? 2'b01 : 2'b11;
					assign node93 = (inp[3]) ? node99 : node94;
						assign node94 = (inp[5]) ? 2'b11 : node95;
							assign node95 = (inp[1]) ? 2'b11 : 2'b01;
						assign node99 = (inp[6]) ? node107 : node100;
							assign node100 = (inp[5]) ? node104 : node101;
								assign node101 = (inp[1]) ? 2'b11 : 2'b01;
								assign node104 = (inp[1]) ? 2'b01 : 2'b11;
							assign node107 = (inp[5]) ? node109 : 2'b01;
								assign node109 = (inp[1]) ? 2'b01 : 2'b11;
		assign node112 = (inp[7]) ? node186 : node113;
			assign node113 = (inp[2]) ? node149 : node114;
				assign node114 = (inp[6]) ? node130 : node115;
					assign node115 = (inp[4]) ? node121 : node116;
						assign node116 = (inp[1]) ? node118 : 2'b10;
							assign node118 = (inp[5]) ? 2'b10 : 2'b00;
						assign node121 = (inp[3]) ? node123 : 2'b00;
							assign node123 = (inp[1]) ? node127 : node124;
								assign node124 = (inp[5]) ? 2'b10 : 2'b00;
								assign node127 = (inp[5]) ? 2'b00 : 2'b10;
					assign node130 = (inp[3]) ? node140 : node131;
						assign node131 = (inp[1]) ? 2'b01 : node132;
							assign node132 = (inp[5]) ? node136 : node133;
								assign node133 = (inp[4]) ? 2'b01 : 2'b11;
								assign node136 = (inp[4]) ? 2'b11 : 2'b01;
						assign node140 = (inp[4]) ? node142 : 2'b11;
							assign node142 = (inp[1]) ? node146 : node143;
								assign node143 = (inp[5]) ? 2'b11 : 2'b01;
								assign node146 = (inp[5]) ? 2'b01 : 2'b11;
				assign node149 = (inp[6]) ? node169 : node150;
					assign node150 = (inp[5]) ? node160 : node151;
						assign node151 = (inp[1]) ? node155 : node152;
							assign node152 = (inp[4]) ? 2'b01 : 2'b11;
							assign node155 = (inp[3]) ? 2'b11 : node156;
								assign node156 = (inp[4]) ? 2'b11 : 2'b01;
						assign node160 = (inp[1]) ? node164 : node161;
							assign node161 = (inp[4]) ? 2'b11 : 2'b01;
							assign node164 = (inp[3]) ? 2'b01 : node165;
								assign node165 = (inp[4]) ? 2'b01 : 2'b11;
					assign node169 = (inp[3]) ? node179 : node170;
						assign node170 = (inp[1]) ? node172 : 2'b11;
							assign node172 = (inp[4]) ? node176 : node173;
								assign node173 = (inp[5]) ? 2'b11 : 2'b01;
								assign node176 = (inp[5]) ? 2'b01 : 2'b11;
						assign node179 = (inp[1]) ? node183 : node180;
							assign node180 = (inp[5]) ? 2'b11 : 2'b01;
							assign node183 = (inp[5]) ? 2'b01 : 2'b11;
			assign node186 = (inp[6]) ? node206 : node187;
				assign node187 = (inp[2]) ? node199 : node188;
					assign node188 = (inp[5]) ? 2'b11 : node189;
						assign node189 = (inp[1]) ? node193 : node190;
							assign node190 = (inp[3]) ? 2'b01 : 2'b11;
							assign node193 = (inp[4]) ? 2'b11 : node194;
								assign node194 = (inp[3]) ? 2'b11 : 2'b01;
					assign node199 = (inp[4]) ? 2'b00 : node200;
						assign node200 = (inp[1]) ? node202 : 2'b00;
							assign node202 = (inp[5]) ? 2'b10 : 2'b00;
				assign node206 = (inp[3]) ? node224 : node207;
					assign node207 = (inp[5]) ? node215 : node208;
						assign node208 = (inp[4]) ? node212 : node209;
							assign node209 = (inp[1]) ? 2'b00 : 2'b10;
							assign node212 = (inp[1]) ? 2'b10 : 2'b00;
						assign node215 = (inp[2]) ? 2'b10 : node216;
							assign node216 = (inp[1]) ? node220 : node217;
								assign node217 = (inp[4]) ? 2'b10 : 2'b00;
								assign node220 = (inp[4]) ? 2'b00 : 2'b10;
					assign node224 = (inp[4]) ? node230 : node225;
						assign node225 = (inp[1]) ? node227 : 2'b00;
							assign node227 = (inp[5]) ? 2'b00 : 2'b10;
						assign node230 = (inp[1]) ? node234 : node231;
							assign node231 = (inp[5]) ? 2'b10 : 2'b00;
							assign node234 = (inp[5]) ? 2'b00 : 2'b10;

endmodule