module dtc_split33_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node16;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node22;
	wire [4-1:0] node26;
	wire [4-1:0] node27;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node59;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node69;
	wire [4-1:0] node72;
	wire [4-1:0] node74;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node86;
	wire [4-1:0] node90;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node98;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node109;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node127;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node136;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node146;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node152;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node175;
	wire [4-1:0] node176;
	wire [4-1:0] node179;
	wire [4-1:0] node181;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node200;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node211;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node218;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node227;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node254;
	wire [4-1:0] node257;
	wire [4-1:0] node260;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node277;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node301;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node307;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node331;
	wire [4-1:0] node332;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node339;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node367;
	wire [4-1:0] node371;
	wire [4-1:0] node373;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node381;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node387;
	wire [4-1:0] node390;
	wire [4-1:0] node394;
	wire [4-1:0] node395;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node423;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node430;
	wire [4-1:0] node431;
	wire [4-1:0] node434;
	wire [4-1:0] node436;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node461;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node477;
	wire [4-1:0] node479;
	wire [4-1:0] node481;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node488;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node496;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node512;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node518;
	wire [4-1:0] node521;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node528;
	wire [4-1:0] node530;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node549;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node562;
	wire [4-1:0] node563;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node571;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node599;
	wire [4-1:0] node601;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node620;
	wire [4-1:0] node622;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node631;
	wire [4-1:0] node634;
	wire [4-1:0] node636;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node643;
	wire [4-1:0] node647;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node658;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node666;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node671;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node685;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node695;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node714;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node721;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node739;
	wire [4-1:0] node742;
	wire [4-1:0] node745;
	wire [4-1:0] node746;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node761;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node775;
	wire [4-1:0] node778;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node803;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node808;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node822;
	wire [4-1:0] node825;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node847;
	wire [4-1:0] node848;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node864;
	wire [4-1:0] node868;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node876;
	wire [4-1:0] node879;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node887;
	wire [4-1:0] node890;
	wire [4-1:0] node893;
	wire [4-1:0] node896;
	wire [4-1:0] node897;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node920;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node944;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node952;
	wire [4-1:0] node954;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node964;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node977;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1005;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1028;
	wire [4-1:0] node1033;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1064;
	wire [4-1:0] node1067;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1090;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1099;
	wire [4-1:0] node1101;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1140;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1155;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1168;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1176;
	wire [4-1:0] node1178;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1197;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1234;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1265;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1286;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1306;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1330;
	wire [4-1:0] node1332;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1377;
	wire [4-1:0] node1380;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1388;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1396;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1411;
	wire [4-1:0] node1414;
	wire [4-1:0] node1415;
	wire [4-1:0] node1416;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1423;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1433;
	wire [4-1:0] node1435;
	wire [4-1:0] node1437;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1445;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1458;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1468;
	wire [4-1:0] node1471;
	wire [4-1:0] node1472;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1487;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1499;
	wire [4-1:0] node1503;
	wire [4-1:0] node1504;
	wire [4-1:0] node1506;
	wire [4-1:0] node1509;
	wire [4-1:0] node1511;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1525;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1533;
	wire [4-1:0] node1536;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1547;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1560;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1565;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1573;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1585;
	wire [4-1:0] node1588;
	wire [4-1:0] node1592;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1596;
	wire [4-1:0] node1598;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1605;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1611;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1618;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1635;
	wire [4-1:0] node1638;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1652;
	wire [4-1:0] node1653;
	wire [4-1:0] node1655;
	wire [4-1:0] node1657;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1675;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1683;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1707;
	wire [4-1:0] node1709;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1721;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1729;
	wire [4-1:0] node1732;
	wire [4-1:0] node1735;
	wire [4-1:0] node1737;
	wire [4-1:0] node1740;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1751;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1757;
	wire [4-1:0] node1760;
	wire [4-1:0] node1762;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1774;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1799;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1812;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1825;
	wire [4-1:0] node1827;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1835;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1847;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1887;
	wire [4-1:0] node1890;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1900;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1918;
	wire [4-1:0] node1921;
	wire [4-1:0] node1922;
	wire [4-1:0] node1924;
	wire [4-1:0] node1927;
	wire [4-1:0] node1929;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1939;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1945;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1958;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1967;
	wire [4-1:0] node1971;
	wire [4-1:0] node1972;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1980;
	wire [4-1:0] node1984;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1991;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2015;
	wire [4-1:0] node2016;
	wire [4-1:0] node2019;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2029;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2039;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2047;
	wire [4-1:0] node2050;
	wire [4-1:0] node2052;
	wire [4-1:0] node2054;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2065;
	wire [4-1:0] node2067;
	wire [4-1:0] node2070;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2083;
	wire [4-1:0] node2086;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2090;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2113;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2118;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2128;
	wire [4-1:0] node2131;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2147;
	wire [4-1:0] node2150;
	wire [4-1:0] node2152;
	wire [4-1:0] node2154;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2165;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2182;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2186;
	wire [4-1:0] node2188;
	wire [4-1:0] node2192;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2205;
	wire [4-1:0] node2208;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2217;
	wire [4-1:0] node2220;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2226;
	wire [4-1:0] node2229;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2250;
	wire [4-1:0] node2254;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2270;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2279;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2293;
	wire [4-1:0] node2294;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2303;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2314;
	wire [4-1:0] node2317;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2320;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2327;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2334;
	wire [4-1:0] node2335;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2343;
	wire [4-1:0] node2346;
	wire [4-1:0] node2347;
	wire [4-1:0] node2349;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2361;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2385;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2390;
	wire [4-1:0] node2394;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2400;
	wire [4-1:0] node2401;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2407;
	wire [4-1:0] node2410;
	wire [4-1:0] node2412;
	wire [4-1:0] node2415;
	wire [4-1:0] node2417;
	wire [4-1:0] node2421;
	wire [4-1:0] node2422;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2426;
	wire [4-1:0] node2427;
	wire [4-1:0] node2428;
	wire [4-1:0] node2430;
	wire [4-1:0] node2431;
	wire [4-1:0] node2437;
	wire [4-1:0] node2438;
	wire [4-1:0] node2441;
	wire [4-1:0] node2443;
	wire [4-1:0] node2446;
	wire [4-1:0] node2447;
	wire [4-1:0] node2449;
	wire [4-1:0] node2451;
	wire [4-1:0] node2453;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2462;
	wire [4-1:0] node2464;
	wire [4-1:0] node2467;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2477;
	wire [4-1:0] node2479;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2484;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2500;
	wire [4-1:0] node2503;
	wire [4-1:0] node2504;
	wire [4-1:0] node2508;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2514;
	wire [4-1:0] node2515;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2524;
	wire [4-1:0] node2525;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2532;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2541;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2549;
	wire [4-1:0] node2550;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2558;
	wire [4-1:0] node2561;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2566;
	wire [4-1:0] node2569;
	wire [4-1:0] node2572;
	wire [4-1:0] node2573;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2584;
	wire [4-1:0] node2587;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2593;
	wire [4-1:0] node2594;
	wire [4-1:0] node2597;
	wire [4-1:0] node2599;
	wire [4-1:0] node2603;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2612;
	wire [4-1:0] node2616;
	wire [4-1:0] node2617;
	wire [4-1:0] node2618;
	wire [4-1:0] node2621;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2627;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2633;
	wire [4-1:0] node2635;
	wire [4-1:0] node2637;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2644;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2664;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2670;
	wire [4-1:0] node2675;
	wire [4-1:0] node2677;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2684;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2692;
	wire [4-1:0] node2694;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2706;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2715;
	wire [4-1:0] node2716;
	wire [4-1:0] node2717;
	wire [4-1:0] node2721;
	wire [4-1:0] node2724;
	wire [4-1:0] node2725;
	wire [4-1:0] node2726;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2733;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2738;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2747;
	wire [4-1:0] node2750;
	wire [4-1:0] node2751;
	wire [4-1:0] node2752;
	wire [4-1:0] node2755;
	wire [4-1:0] node2758;
	wire [4-1:0] node2759;
	wire [4-1:0] node2764;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2770;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2790;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2795;
	wire [4-1:0] node2798;
	wire [4-1:0] node2801;
	wire [4-1:0] node2802;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2811;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2817;
	wire [4-1:0] node2820;
	wire [4-1:0] node2822;
	wire [4-1:0] node2824;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2833;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2840;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2853;
	wire [4-1:0] node2854;
	wire [4-1:0] node2858;
	wire [4-1:0] node2861;
	wire [4-1:0] node2862;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2868;
	wire [4-1:0] node2871;
	wire [4-1:0] node2874;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2880;
	wire [4-1:0] node2882;
	wire [4-1:0] node2886;
	wire [4-1:0] node2887;
	wire [4-1:0] node2888;
	wire [4-1:0] node2889;
	wire [4-1:0] node2890;
	wire [4-1:0] node2892;
	wire [4-1:0] node2894;
	wire [4-1:0] node2896;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2906;
	wire [4-1:0] node2907;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2914;
	wire [4-1:0] node2917;
	wire [4-1:0] node2919;
	wire [4-1:0] node2920;
	wire [4-1:0] node2924;
	wire [4-1:0] node2926;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2937;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2948;
	wire [4-1:0] node2949;
	wire [4-1:0] node2952;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2958;
	wire [4-1:0] node2960;
	wire [4-1:0] node2961;
	wire [4-1:0] node2965;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2975;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2981;
	wire [4-1:0] node2982;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2992;
	wire [4-1:0] node2994;
	wire [4-1:0] node2997;
	wire [4-1:0] node2999;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3009;
	wire [4-1:0] node3012;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3030;
	wire [4-1:0] node3031;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3038;
	wire [4-1:0] node3039;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3054;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3062;
	wire [4-1:0] node3063;
	wire [4-1:0] node3066;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3073;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3086;
	wire [4-1:0] node3087;
	wire [4-1:0] node3090;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3096;
	wire [4-1:0] node3098;
	wire [4-1:0] node3102;
	wire [4-1:0] node3105;
	wire [4-1:0] node3106;
	wire [4-1:0] node3107;
	wire [4-1:0] node3108;
	wire [4-1:0] node3109;
	wire [4-1:0] node3111;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3117;
	wire [4-1:0] node3120;
	wire [4-1:0] node3123;
	wire [4-1:0] node3124;
	wire [4-1:0] node3125;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3151;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3158;
	wire [4-1:0] node3160;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3172;
	wire [4-1:0] node3173;
	wire [4-1:0] node3175;
	wire [4-1:0] node3178;
	wire [4-1:0] node3180;
	wire [4-1:0] node3182;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3191;
	wire [4-1:0] node3192;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3200;
	wire [4-1:0] node3202;
	wire [4-1:0] node3203;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3210;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3215;
	wire [4-1:0] node3219;
	wire [4-1:0] node3221;
	wire [4-1:0] node3222;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3235;
	wire [4-1:0] node3237;
	wire [4-1:0] node3240;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3246;
	wire [4-1:0] node3248;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3255;
	wire [4-1:0] node3259;
	wire [4-1:0] node3261;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3268;
	wire [4-1:0] node3271;
	wire [4-1:0] node3273;
	wire [4-1:0] node3275;
	wire [4-1:0] node3278;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3282;
	wire [4-1:0] node3284;
	wire [4-1:0] node3287;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3300;
	wire [4-1:0] node3301;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3313;
	wire [4-1:0] node3315;
	wire [4-1:0] node3316;
	wire [4-1:0] node3318;
	wire [4-1:0] node3322;
	wire [4-1:0] node3323;
	wire [4-1:0] node3324;
	wire [4-1:0] node3325;
	wire [4-1:0] node3326;
	wire [4-1:0] node3330;
	wire [4-1:0] node3333;
	wire [4-1:0] node3334;
	wire [4-1:0] node3338;
	wire [4-1:0] node3339;
	wire [4-1:0] node3341;
	wire [4-1:0] node3343;
	wire [4-1:0] node3344;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3352;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3357;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3366;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3372;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3383;
	wire [4-1:0] node3384;
	wire [4-1:0] node3387;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3394;
	wire [4-1:0] node3395;
	wire [4-1:0] node3396;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3401;
	wire [4-1:0] node3405;
	wire [4-1:0] node3409;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3434;
	wire [4-1:0] node3437;
	wire [4-1:0] node3439;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3446;
	wire [4-1:0] node3448;
	wire [4-1:0] node3450;
	wire [4-1:0] node3453;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3463;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3474;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3486;
	wire [4-1:0] node3488;
	wire [4-1:0] node3490;
	wire [4-1:0] node3492;
	wire [4-1:0] node3497;
	wire [4-1:0] node3498;
	wire [4-1:0] node3499;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3505;
	wire [4-1:0] node3507;
	wire [4-1:0] node3508;
	wire [4-1:0] node3510;
	wire [4-1:0] node3512;
	wire [4-1:0] node3516;
	wire [4-1:0] node3517;
	wire [4-1:0] node3519;
	wire [4-1:0] node3522;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3527;
	wire [4-1:0] node3530;
	wire [4-1:0] node3532;
	wire [4-1:0] node3534;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3545;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3551;
	wire [4-1:0] node3554;
	wire [4-1:0] node3555;
	wire [4-1:0] node3556;
	wire [4-1:0] node3560;
	wire [4-1:0] node3561;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3575;
	wire [4-1:0] node3579;
	wire [4-1:0] node3582;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3587;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3596;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3613;
	wire [4-1:0] node3614;
	wire [4-1:0] node3616;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3624;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3633;
	wire [4-1:0] node3634;
	wire [4-1:0] node3638;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3647;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3658;
	wire [4-1:0] node3660;
	wire [4-1:0] node3663;
	wire [4-1:0] node3666;
	wire [4-1:0] node3667;
	wire [4-1:0] node3668;
	wire [4-1:0] node3672;
	wire [4-1:0] node3673;
	wire [4-1:0] node3674;
	wire [4-1:0] node3679;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3683;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3694;
	wire [4-1:0] node3697;
	wire [4-1:0] node3698;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3709;
	wire [4-1:0] node3711;
	wire [4-1:0] node3714;
	wire [4-1:0] node3716;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3725;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3733;
	wire [4-1:0] node3735;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3741;
	wire [4-1:0] node3744;
	wire [4-1:0] node3745;
	wire [4-1:0] node3747;
	wire [4-1:0] node3751;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3763;
	wire [4-1:0] node3765;
	wire [4-1:0] node3767;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3772;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3779;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3785;
	wire [4-1:0] node3786;
	wire [4-1:0] node3788;
	wire [4-1:0] node3792;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3801;
	wire [4-1:0] node3804;
	wire [4-1:0] node3806;
	wire [4-1:0] node3807;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3820;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3824;
	wire [4-1:0] node3825;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3830;
	wire [4-1:0] node3833;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3841;
	wire [4-1:0] node3842;
	wire [4-1:0] node3844;
	wire [4-1:0] node3847;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3856;
	wire [4-1:0] node3858;
	wire [4-1:0] node3861;
	wire [4-1:0] node3863;
	wire [4-1:0] node3865;
	wire [4-1:0] node3866;
	wire [4-1:0] node3867;
	wire [4-1:0] node3869;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3882;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3890;
	wire [4-1:0] node3892;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3900;
	wire [4-1:0] node3901;
	wire [4-1:0] node3903;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3911;
	wire [4-1:0] node3912;
	wire [4-1:0] node3913;
	wire [4-1:0] node3916;
	wire [4-1:0] node3919;
	wire [4-1:0] node3921;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3931;
	wire [4-1:0] node3933;
	wire [4-1:0] node3936;
	wire [4-1:0] node3938;
	wire [4-1:0] node3940;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3947;
	wire [4-1:0] node3951;
	wire [4-1:0] node3953;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3960;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3970;
	wire [4-1:0] node3971;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3976;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3987;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3990;
	wire [4-1:0] node3991;
	wire [4-1:0] node3994;
	wire [4-1:0] node3997;
	wire [4-1:0] node3999;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4006;
	wire [4-1:0] node4007;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4014;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4037;
	wire [4-1:0] node4038;
	wire [4-1:0] node4040;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4047;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4055;
	wire [4-1:0] node4058;
	wire [4-1:0] node4059;
	wire [4-1:0] node4063;
	wire [4-1:0] node4064;
	wire [4-1:0] node4067;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4075;
	wire [4-1:0] node4076;
	wire [4-1:0] node4077;
	wire [4-1:0] node4081;
	wire [4-1:0] node4084;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4093;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4099;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4108;
	wire [4-1:0] node4110;
	wire [4-1:0] node4114;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4123;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4141;
	wire [4-1:0] node4144;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4153;
	wire [4-1:0] node4154;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4161;
	wire [4-1:0] node4162;
	wire [4-1:0] node4163;
	wire [4-1:0] node4166;
	wire [4-1:0] node4170;
	wire [4-1:0] node4173;
	wire [4-1:0] node4174;
	wire [4-1:0] node4175;
	wire [4-1:0] node4176;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4186;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4196;
	wire [4-1:0] node4198;
	wire [4-1:0] node4201;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4211;
	wire [4-1:0] node4214;
	wire [4-1:0] node4215;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4222;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4233;
	wire [4-1:0] node4237;
	wire [4-1:0] node4238;
	wire [4-1:0] node4241;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4248;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4258;
	wire [4-1:0] node4260;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4265;
	wire [4-1:0] node4266;
	wire [4-1:0] node4268;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4275;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4283;
	wire [4-1:0] node4285;
	wire [4-1:0] node4288;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4294;
	wire [4-1:0] node4297;
	wire [4-1:0] node4300;
	wire [4-1:0] node4301;
	wire [4-1:0] node4305;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4311;
	wire [4-1:0] node4312;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4332;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4342;
	wire [4-1:0] node4343;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4369;
	wire [4-1:0] node4372;
	wire [4-1:0] node4373;
	wire [4-1:0] node4376;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4382;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4400;
	wire [4-1:0] node4401;
	wire [4-1:0] node4402;
	wire [4-1:0] node4404;
	wire [4-1:0] node4408;
	wire [4-1:0] node4410;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4415;
	wire [4-1:0] node4416;
	wire [4-1:0] node4417;
	wire [4-1:0] node4418;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4431;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4435;
	wire [4-1:0] node4437;
	wire [4-1:0] node4440;
	wire [4-1:0] node4444;
	wire [4-1:0] node4445;
	wire [4-1:0] node4449;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4455;
	wire [4-1:0] node4459;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4466;
	wire [4-1:0] node4467;
	wire [4-1:0] node4468;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4474;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4495;
	wire [4-1:0] node4499;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4528;
	wire [4-1:0] node4531;
	wire [4-1:0] node4532;
	wire [4-1:0] node4534;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4541;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4549;
	wire [4-1:0] node4552;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4562;
	wire [4-1:0] node4563;
	wire [4-1:0] node4564;
	wire [4-1:0] node4565;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4569;
	wire [4-1:0] node4573;
	wire [4-1:0] node4574;
	wire [4-1:0] node4576;
	wire [4-1:0] node4578;
	wire [4-1:0] node4581;
	wire [4-1:0] node4583;
	wire [4-1:0] node4586;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4594;
	wire [4-1:0] node4596;
	wire [4-1:0] node4598;
	wire [4-1:0] node4601;
	wire [4-1:0] node4602;
	wire [4-1:0] node4603;
	wire [4-1:0] node4604;
	wire [4-1:0] node4606;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4613;
	wire [4-1:0] node4616;
	wire [4-1:0] node4617;
	wire [4-1:0] node4618;
	wire [4-1:0] node4621;
	wire [4-1:0] node4623;
	wire [4-1:0] node4626;
	wire [4-1:0] node4629;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4634;
	wire [4-1:0] node4636;
	wire [4-1:0] node4639;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4651;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4656;
	wire [4-1:0] node4657;
	wire [4-1:0] node4662;
	wire [4-1:0] node4663;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4676;
	wire [4-1:0] node4677;
	wire [4-1:0] node4680;
	wire [4-1:0] node4684;
	wire [4-1:0] node4685;
	wire [4-1:0] node4686;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4692;
	wire [4-1:0] node4693;
	wire [4-1:0] node4697;
	wire [4-1:0] node4698;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4705;
	wire [4-1:0] node4708;
	wire [4-1:0] node4711;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4717;
	wire [4-1:0] node4718;
	wire [4-1:0] node4720;
	wire [4-1:0] node4725;
	wire [4-1:0] node4726;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4734;
	wire [4-1:0] node4736;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4747;
	wire [4-1:0] node4749;
	wire [4-1:0] node4752;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4756;
	wire [4-1:0] node4760;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4765;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4772;
	wire [4-1:0] node4773;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4782;
	wire [4-1:0] node4787;
	wire [4-1:0] node4788;
	wire [4-1:0] node4791;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4800;
	wire [4-1:0] node4803;
	wire [4-1:0] node4806;
	wire [4-1:0] node4809;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4818;
	wire [4-1:0] node4821;
	wire [4-1:0] node4822;
	wire [4-1:0] node4824;
	wire [4-1:0] node4826;
	wire [4-1:0] node4829;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4836;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4844;
	wire [4-1:0] node4846;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4852;
	wire [4-1:0] node4856;
	wire [4-1:0] node4858;
	wire [4-1:0] node4860;
	wire [4-1:0] node4863;
	wire [4-1:0] node4864;
	wire [4-1:0] node4865;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4869;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4881;
	wire [4-1:0] node4882;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4894;
	wire [4-1:0] node4897;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4904;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4918;
	wire [4-1:0] node4919;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4926;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4932;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4938;
	wire [4-1:0] node4939;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4949;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4955;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4972;
	wire [4-1:0] node4976;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4982;
	wire [4-1:0] node4983;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4994;
	wire [4-1:0] node4996;
	wire [4-1:0] node4999;
	wire [4-1:0] node5001;
	wire [4-1:0] node5002;
	wire [4-1:0] node5005;
	wire [4-1:0] node5007;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5015;
	wire [4-1:0] node5017;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5029;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5036;
	wire [4-1:0] node5037;
	wire [4-1:0] node5038;
	wire [4-1:0] node5040;
	wire [4-1:0] node5042;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5051;
	wire [4-1:0] node5052;
	wire [4-1:0] node5053;
	wire [4-1:0] node5057;
	wire [4-1:0] node5058;
	wire [4-1:0] node5061;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5066;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5078;
	wire [4-1:0] node5080;
	wire [4-1:0] node5081;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5087;
	wire [4-1:0] node5089;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5100;
	wire [4-1:0] node5101;
	wire [4-1:0] node5102;
	wire [4-1:0] node5104;
	wire [4-1:0] node5108;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5115;
	wire [4-1:0] node5118;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5126;
	wire [4-1:0] node5128;
	wire [4-1:0] node5132;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5136;
	wire [4-1:0] node5138;
	wire [4-1:0] node5140;
	wire [4-1:0] node5143;
	wire [4-1:0] node5144;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5151;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5161;
	wire [4-1:0] node5165;
	wire [4-1:0] node5167;
	wire [4-1:0] node5170;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5175;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5189;
	wire [4-1:0] node5191;
	wire [4-1:0] node5194;
	wire [4-1:0] node5195;
	wire [4-1:0] node5196;
	wire [4-1:0] node5198;
	wire [4-1:0] node5201;
	wire [4-1:0] node5204;
	wire [4-1:0] node5205;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5215;
	wire [4-1:0] node5216;
	wire [4-1:0] node5222;
	wire [4-1:0] node5223;
	wire [4-1:0] node5224;
	wire [4-1:0] node5225;
	wire [4-1:0] node5226;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5238;
	wire [4-1:0] node5242;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5252;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5265;
	wire [4-1:0] node5271;
	wire [4-1:0] node5272;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5277;
	wire [4-1:0] node5278;
	wire [4-1:0] node5279;
	wire [4-1:0] node5281;
	wire [4-1:0] node5282;
	wire [4-1:0] node5284;
	wire [4-1:0] node5286;
	wire [4-1:0] node5288;
	wire [4-1:0] node5291;
	wire [4-1:0] node5292;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5302;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5309;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5315;
	wire [4-1:0] node5318;
	wire [4-1:0] node5321;
	wire [4-1:0] node5323;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5329;
	wire [4-1:0] node5332;
	wire [4-1:0] node5334;
	wire [4-1:0] node5337;
	wire [4-1:0] node5340;
	wire [4-1:0] node5341;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5346;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5354;
	wire [4-1:0] node5356;
	wire [4-1:0] node5359;
	wire [4-1:0] node5360;
	wire [4-1:0] node5363;
	wire [4-1:0] node5365;
	wire [4-1:0] node5367;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5383;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5390;
	wire [4-1:0] node5391;
	wire [4-1:0] node5395;
	wire [4-1:0] node5397;
	wire [4-1:0] node5399;
	wire [4-1:0] node5400;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5407;
	wire [4-1:0] node5409;
	wire [4-1:0] node5412;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5418;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5427;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5433;
	wire [4-1:0] node5435;
	wire [4-1:0] node5439;
	wire [4-1:0] node5440;
	wire [4-1:0] node5441;
	wire [4-1:0] node5444;
	wire [4-1:0] node5446;
	wire [4-1:0] node5450;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5454;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5463;
	wire [4-1:0] node5466;
	wire [4-1:0] node5469;
	wire [4-1:0] node5470;
	wire [4-1:0] node5471;
	wire [4-1:0] node5473;
	wire [4-1:0] node5474;
	wire [4-1:0] node5477;
	wire [4-1:0] node5479;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5484;
	wire [4-1:0] node5487;
	wire [4-1:0] node5489;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5504;
	wire [4-1:0] node5505;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5513;
	wire [4-1:0] node5514;
	wire [4-1:0] node5516;
	wire [4-1:0] node5520;
	wire [4-1:0] node5522;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5536;
	wire [4-1:0] node5537;
	wire [4-1:0] node5540;
	wire [4-1:0] node5544;
	wire [4-1:0] node5546;
	wire [4-1:0] node5549;
	wire [4-1:0] node5551;
	wire [4-1:0] node5553;
	wire [4-1:0] node5554;
	wire [4-1:0] node5555;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5565;
	wire [4-1:0] node5568;
	wire [4-1:0] node5569;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5588;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5596;
	wire [4-1:0] node5599;
	wire [4-1:0] node5601;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5609;
	wire [4-1:0] node5611;
	wire [4-1:0] node5612;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5623;
	wire [4-1:0] node5626;
	wire [4-1:0] node5627;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5635;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5645;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5656;
	wire [4-1:0] node5659;
	wire [4-1:0] node5662;
	wire [4-1:0] node5663;
	wire [4-1:0] node5664;
	wire [4-1:0] node5667;
	wire [4-1:0] node5669;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5676;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5683;
	wire [4-1:0] node5684;
	wire [4-1:0] node5685;
	wire [4-1:0] node5686;
	wire [4-1:0] node5687;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5696;
	wire [4-1:0] node5697;
	wire [4-1:0] node5698;
	wire [4-1:0] node5700;
	wire [4-1:0] node5704;
	wire [4-1:0] node5706;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5716;
	wire [4-1:0] node5718;
	wire [4-1:0] node5721;
	wire [4-1:0] node5722;
	wire [4-1:0] node5723;
	wire [4-1:0] node5725;
	wire [4-1:0] node5729;
	wire [4-1:0] node5731;
	wire [4-1:0] node5734;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5738;
	wire [4-1:0] node5739;
	wire [4-1:0] node5742;
	wire [4-1:0] node5744;
	wire [4-1:0] node5745;
	wire [4-1:0] node5749;
	wire [4-1:0] node5750;
	wire [4-1:0] node5751;
	wire [4-1:0] node5752;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5761;
	wire [4-1:0] node5763;
	wire [4-1:0] node5765;
	wire [4-1:0] node5768;
	wire [4-1:0] node5769;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5778;
	wire [4-1:0] node5781;
	wire [4-1:0] node5785;
	wire [4-1:0] node5786;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5793;
	wire [4-1:0] node5794;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5800;
	wire [4-1:0] node5802;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5809;
	wire [4-1:0] node5811;
	wire [4-1:0] node5814;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5820;
	wire [4-1:0] node5822;
	wire [4-1:0] node5824;
	wire [4-1:0] node5827;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5833;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5842;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5847;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5853;
	wire [4-1:0] node5856;
	wire [4-1:0] node5858;
	wire [4-1:0] node5861;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5872;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5878;
	wire [4-1:0] node5883;
	wire [4-1:0] node5886;
	wire [4-1:0] node5887;
	wire [4-1:0] node5888;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5897;
	wire [4-1:0] node5898;
	wire [4-1:0] node5900;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5909;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5918;
	wire [4-1:0] node5921;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5928;
	wire [4-1:0] node5929;
	wire [4-1:0] node5930;
	wire [4-1:0] node5933;
	wire [4-1:0] node5936;
	wire [4-1:0] node5939;
	wire [4-1:0] node5940;
	wire [4-1:0] node5941;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5947;
	wire [4-1:0] node5950;
	wire [4-1:0] node5952;
	wire [4-1:0] node5954;
	wire [4-1:0] node5957;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5974;
	wire [4-1:0] node5975;
	wire [4-1:0] node5977;
	wire [4-1:0] node5979;
	wire [4-1:0] node5982;
	wire [4-1:0] node5984;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5994;
	wire [4-1:0] node5999;
	wire [4-1:0] node6000;
	wire [4-1:0] node6002;
	wire [4-1:0] node6003;
	wire [4-1:0] node6007;
	wire [4-1:0] node6008;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6015;
	wire [4-1:0] node6019;
	wire [4-1:0] node6021;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6027;
	wire [4-1:0] node6028;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6031;
	wire [4-1:0] node6034;
	wire [4-1:0] node6036;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6048;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6055;
	wire [4-1:0] node6059;
	wire [4-1:0] node6060;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6076;
	wire [4-1:0] node6080;
	wire [4-1:0] node6083;
	wire [4-1:0] node6084;
	wire [4-1:0] node6086;
	wire [4-1:0] node6087;
	wire [4-1:0] node6090;
	wire [4-1:0] node6093;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6102;
	wire [4-1:0] node6105;
	wire [4-1:0] node6107;
	wire [4-1:0] node6108;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6117;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6125;
	wire [4-1:0] node6127;
	wire [4-1:0] node6130;
	wire [4-1:0] node6131;
	wire [4-1:0] node6132;
	wire [4-1:0] node6134;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6140;
	wire [4-1:0] node6144;
	wire [4-1:0] node6145;
	wire [4-1:0] node6146;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6155;
	wire [4-1:0] node6156;
	wire [4-1:0] node6157;
	wire [4-1:0] node6158;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6164;
	wire [4-1:0] node6166;
	wire [4-1:0] node6167;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6180;
	wire [4-1:0] node6181;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6194;
	wire [4-1:0] node6197;
	wire [4-1:0] node6200;
	wire [4-1:0] node6201;
	wire [4-1:0] node6202;
	wire [4-1:0] node6205;
	wire [4-1:0] node6207;
	wire [4-1:0] node6210;
	wire [4-1:0] node6212;
	wire [4-1:0] node6214;
	wire [4-1:0] node6217;
	wire [4-1:0] node6218;
	wire [4-1:0] node6219;
	wire [4-1:0] node6220;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6227;
	wire [4-1:0] node6229;
	wire [4-1:0] node6232;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6238;
	wire [4-1:0] node6240;
	wire [4-1:0] node6243;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6249;
	wire [4-1:0] node6252;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6258;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6265;
	wire [4-1:0] node6266;
	wire [4-1:0] node6268;
	wire [4-1:0] node6269;
	wire [4-1:0] node6272;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6279;
	wire [4-1:0] node6281;
	wire [4-1:0] node6284;
	wire [4-1:0] node6285;
	wire [4-1:0] node6287;
	wire [4-1:0] node6289;
	wire [4-1:0] node6292;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6298;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6317;
	wire [4-1:0] node6322;
	wire [4-1:0] node6323;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6335;
	wire [4-1:0] node6337;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6342;
	wire [4-1:0] node6344;
	wire [4-1:0] node6347;
	wire [4-1:0] node6348;
	wire [4-1:0] node6353;
	wire [4-1:0] node6355;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6364;
	wire [4-1:0] node6365;
	wire [4-1:0] node6367;
	wire [4-1:0] node6368;
	wire [4-1:0] node6370;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6379;
	wire [4-1:0] node6380;
	wire [4-1:0] node6381;
	wire [4-1:0] node6384;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6390;
	wire [4-1:0] node6391;
	wire [4-1:0] node6396;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6401;
	wire [4-1:0] node6402;
	wire [4-1:0] node6405;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6413;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6417;
	wire [4-1:0] node6421;
	wire [4-1:0] node6423;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6429;
	wire [4-1:0] node6433;
	wire [4-1:0] node6435;
	wire [4-1:0] node6436;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6449;
	wire [4-1:0] node6450;
	wire [4-1:0] node6452;
	wire [4-1:0] node6453;
	wire [4-1:0] node6456;
	wire [4-1:0] node6458;
	wire [4-1:0] node6461;
	wire [4-1:0] node6462;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6476;
	wire [4-1:0] node6477;
	wire [4-1:0] node6480;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6494;
	wire [4-1:0] node6496;
	wire [4-1:0] node6498;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6503;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6521;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6527;
	wire [4-1:0] node6530;
	wire [4-1:0] node6533;
	wire [4-1:0] node6535;
	wire [4-1:0] node6538;
	wire [4-1:0] node6540;
	wire [4-1:0] node6541;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6548;
	wire [4-1:0] node6549;
	wire [4-1:0] node6552;
	wire [4-1:0] node6554;
	wire [4-1:0] node6557;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6563;
	wire [4-1:0] node6565;
	wire [4-1:0] node6566;
	wire [4-1:0] node6570;
	wire [4-1:0] node6571;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6591;
	wire [4-1:0] node6598;
	wire [4-1:0] node6599;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6605;
	wire [4-1:0] node6608;
	wire [4-1:0] node6611;
	wire [4-1:0] node6615;
	wire [4-1:0] node6617;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6622;
	wire [4-1:0] node6624;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6632;
	wire [4-1:0] node6634;
	wire [4-1:0] node6637;
	wire [4-1:0] node6638;
	wire [4-1:0] node6640;
	wire [4-1:0] node6643;
	wire [4-1:0] node6644;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6650;
	wire [4-1:0] node6654;
	wire [4-1:0] node6655;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6666;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6674;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6684;
	wire [4-1:0] node6687;
	wire [4-1:0] node6689;
	wire [4-1:0] node6690;
	wire [4-1:0] node6692;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6699;
	wire [4-1:0] node6700;
	wire [4-1:0] node6701;
	wire [4-1:0] node6703;
	wire [4-1:0] node6706;
	wire [4-1:0] node6709;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6721;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6726;
	wire [4-1:0] node6731;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6735;
	wire [4-1:0] node6737;
	wire [4-1:0] node6738;
	wire [4-1:0] node6741;
	wire [4-1:0] node6745;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6750;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6756;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6760;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6769;
	wire [4-1:0] node6772;
	wire [4-1:0] node6775;
	wire [4-1:0] node6776;
	wire [4-1:0] node6778;
	wire [4-1:0] node6780;
	wire [4-1:0] node6783;
	wire [4-1:0] node6785;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6791;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6800;
	wire [4-1:0] node6801;
	wire [4-1:0] node6802;
	wire [4-1:0] node6805;
	wire [4-1:0] node6808;
	wire [4-1:0] node6810;
	wire [4-1:0] node6813;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6817;
	wire [4-1:0] node6819;
	wire [4-1:0] node6822;
	wire [4-1:0] node6824;
	wire [4-1:0] node6827;
	wire [4-1:0] node6828;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6842;
	wire [4-1:0] node6843;
	wire [4-1:0] node6844;
	wire [4-1:0] node6845;
	wire [4-1:0] node6847;
	wire [4-1:0] node6848;
	wire [4-1:0] node6851;
	wire [4-1:0] node6854;
	wire [4-1:0] node6855;
	wire [4-1:0] node6856;
	wire [4-1:0] node6859;
	wire [4-1:0] node6860;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6872;
	wire [4-1:0] node6873;
	wire [4-1:0] node6876;
	wire [4-1:0] node6878;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6887;
	wire [4-1:0] node6888;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6895;
	wire [4-1:0] node6897;
	wire [4-1:0] node6901;
	wire [4-1:0] node6903;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6908;
	wire [4-1:0] node6911;
	wire [4-1:0] node6913;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6932;
	wire [4-1:0] node6936;
	wire [4-1:0] node6938;
	wire [4-1:0] node6939;
	wire [4-1:0] node6940;
	wire [4-1:0] node6944;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6949;
	wire [4-1:0] node6950;
	wire [4-1:0] node6953;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6961;
	wire [4-1:0] node6962;
	wire [4-1:0] node6964;
	wire [4-1:0] node6967;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6972;
	wire [4-1:0] node6974;
	wire [4-1:0] node6977;
	wire [4-1:0] node6979;
	wire [4-1:0] node6981;
	wire [4-1:0] node6983;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6993;
	wire [4-1:0] node6994;
	wire [4-1:0] node6998;
	wire [4-1:0] node6999;
	wire [4-1:0] node7001;
	wire [4-1:0] node7002;
	wire [4-1:0] node7005;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7011;
	wire [4-1:0] node7012;
	wire [4-1:0] node7013;
	wire [4-1:0] node7014;
	wire [4-1:0] node7015;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7025;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7034;
	wire [4-1:0] node7035;
	wire [4-1:0] node7038;
	wire [4-1:0] node7039;
	wire [4-1:0] node7042;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7059;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7067;
	wire [4-1:0] node7068;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7079;
	wire [4-1:0] node7081;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7088;
	wire [4-1:0] node7091;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7096;
	wire [4-1:0] node7099;
	wire [4-1:0] node7101;
	wire [4-1:0] node7104;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7108;
	wire [4-1:0] node7112;
	wire [4-1:0] node7113;
	wire [4-1:0] node7114;
	wire [4-1:0] node7119;
	wire [4-1:0] node7120;
	wire [4-1:0] node7121;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7127;
	wire [4-1:0] node7128;
	wire [4-1:0] node7132;
	wire [4-1:0] node7134;
	wire [4-1:0] node7135;
	wire [4-1:0] node7137;
	wire [4-1:0] node7140;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7145;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7152;
	wire [4-1:0] node7154;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7163;
	wire [4-1:0] node7165;
	wire [4-1:0] node7168;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7173;
	wire [4-1:0] node7175;
	wire [4-1:0] node7179;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7187;
	wire [4-1:0] node7188;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7201;
	wire [4-1:0] node7203;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7210;
	wire [4-1:0] node7213;
	wire [4-1:0] node7215;
	wire [4-1:0] node7218;
	wire [4-1:0] node7220;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7236;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7244;
	wire [4-1:0] node7245;
	wire [4-1:0] node7246;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7258;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7276;
	wire [4-1:0] node7278;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7286;
	wire [4-1:0] node7287;
	wire [4-1:0] node7291;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7299;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7308;
	wire [4-1:0] node7310;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7317;
	wire [4-1:0] node7319;
	wire [4-1:0] node7322;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7326;
	wire [4-1:0] node7328;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7339;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7351;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7362;
	wire [4-1:0] node7364;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7371;
	wire [4-1:0] node7372;
	wire [4-1:0] node7375;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7385;
	wire [4-1:0] node7386;
	wire [4-1:0] node7390;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7404;
	wire [4-1:0] node7408;
	wire [4-1:0] node7409;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7419;
	wire [4-1:0] node7422;
	wire [4-1:0] node7423;
	wire [4-1:0] node7427;
	wire [4-1:0] node7429;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7434;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7445;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7450;
	wire [4-1:0] node7455;
	wire [4-1:0] node7457;
	wire [4-1:0] node7459;
	wire [4-1:0] node7462;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7468;
	wire [4-1:0] node7471;
	wire [4-1:0] node7474;
	wire [4-1:0] node7475;
	wire [4-1:0] node7476;
	wire [4-1:0] node7480;
	wire [4-1:0] node7481;
	wire [4-1:0] node7483;
	wire [4-1:0] node7486;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7497;
	wire [4-1:0] node7499;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7504;
	wire [4-1:0] node7508;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7513;
	wire [4-1:0] node7514;
	wire [4-1:0] node7518;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7525;
	wire [4-1:0] node7526;
	wire [4-1:0] node7527;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7533;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7541;
	wire [4-1:0] node7544;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7547;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7557;
	wire [4-1:0] node7560;
	wire [4-1:0] node7561;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7568;
	wire [4-1:0] node7571;
	wire [4-1:0] node7572;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7586;
	wire [4-1:0] node7590;
	wire [4-1:0] node7591;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7600;
	wire [4-1:0] node7603;
	wire [4-1:0] node7604;
	wire [4-1:0] node7605;
	wire [4-1:0] node7607;
	wire [4-1:0] node7609;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7616;
	wire [4-1:0] node7617;
	wire [4-1:0] node7620;
	wire [4-1:0] node7623;
	wire [4-1:0] node7625;
	wire [4-1:0] node7627;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7642;
	wire [4-1:0] node7646;
	wire [4-1:0] node7648;
	wire [4-1:0] node7651;
	wire [4-1:0] node7653;
	wire [4-1:0] node7655;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7661;
	wire [4-1:0] node7662;
	wire [4-1:0] node7666;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7671;
	wire [4-1:0] node7673;
	wire [4-1:0] node7676;
	wire [4-1:0] node7679;
	wire [4-1:0] node7680;
	wire [4-1:0] node7681;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7687;
	wire [4-1:0] node7690;
	wire [4-1:0] node7692;
	wire [4-1:0] node7693;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7703;
	wire [4-1:0] node7706;
	wire [4-1:0] node7708;
	wire [4-1:0] node7709;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7716;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7723;
	wire [4-1:0] node7725;
	wire [4-1:0] node7728;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7742;
	wire [4-1:0] node7746;
	wire [4-1:0] node7747;
	wire [4-1:0] node7751;
	wire [4-1:0] node7752;
	wire [4-1:0] node7754;
	wire [4-1:0] node7757;
	wire [4-1:0] node7760;
	wire [4-1:0] node7761;
	wire [4-1:0] node7762;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7768;
	wire [4-1:0] node7770;
	wire [4-1:0] node7772;
	wire [4-1:0] node7775;
	wire [4-1:0] node7777;
	wire [4-1:0] node7779;
	wire [4-1:0] node7782;
	wire [4-1:0] node7783;
	wire [4-1:0] node7784;
	wire [4-1:0] node7787;
	wire [4-1:0] node7788;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7795;
	wire [4-1:0] node7796;
	wire [4-1:0] node7799;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7807;
	wire [4-1:0] node7810;
	wire [4-1:0] node7811;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7818;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7822;
	wire [4-1:0] node7824;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7830;
	wire [4-1:0] node7833;
	wire [4-1:0] node7835;
	wire [4-1:0] node7838;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7841;
	wire [4-1:0] node7844;
	wire [4-1:0] node7845;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7860;
	wire [4-1:0] node7863;
	wire [4-1:0] node7864;
	wire [4-1:0] node7865;
	wire [4-1:0] node7866;
	wire [4-1:0] node7867;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7879;
	wire [4-1:0] node7881;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7894;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7913;
	wire [4-1:0] node7915;
	wire [4-1:0] node7917;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7926;
	wire [4-1:0] node7929;
	wire [4-1:0] node7931;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7940;
	wire [4-1:0] node7945;
	wire [4-1:0] node7946;
	wire [4-1:0] node7947;
	wire [4-1:0] node7949;
	wire [4-1:0] node7951;
	wire [4-1:0] node7954;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7959;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7964;
	wire [4-1:0] node7968;
	wire [4-1:0] node7971;
	wire [4-1:0] node7974;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7980;
	wire [4-1:0] node7985;
	wire [4-1:0] node7986;
	wire [4-1:0] node7988;
	wire [4-1:0] node7991;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node7997;
	wire [4-1:0] node7998;
	wire [4-1:0] node7999;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8005;
	wire [4-1:0] node8007;
	wire [4-1:0] node8009;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8016;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8024;
	wire [4-1:0] node8025;
	wire [4-1:0] node8029;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8034;
	wire [4-1:0] node8035;
	wire [4-1:0] node8037;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8051;
	wire [4-1:0] node8053;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8061;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8069;
	wire [4-1:0] node8071;
	wire [4-1:0] node8074;
	wire [4-1:0] node8075;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8083;
	wire [4-1:0] node8085;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8100;
	wire [4-1:0] node8102;
	wire [4-1:0] node8105;
	wire [4-1:0] node8106;
	wire [4-1:0] node8109;
	wire [4-1:0] node8112;
	wire [4-1:0] node8114;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8120;
	wire [4-1:0] node8123;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8127;
	wire [4-1:0] node8128;
	wire [4-1:0] node8132;
	wire [4-1:0] node8133;
	wire [4-1:0] node8134;
	wire [4-1:0] node8137;
	wire [4-1:0] node8141;
	wire [4-1:0] node8142;
	wire [4-1:0] node8143;
	wire [4-1:0] node8146;
	wire [4-1:0] node8150;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8156;
	wire [4-1:0] node8160;
	wire [4-1:0] node8161;
	wire [4-1:0] node8163;
	wire [4-1:0] node8167;
	wire [4-1:0] node8168;
	wire [4-1:0] node8169;
	wire [4-1:0] node8170;
	wire [4-1:0] node8171;
	wire [4-1:0] node8176;
	wire [4-1:0] node8177;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8185;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8198;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8201;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8207;
	wire [4-1:0] node8209;
	wire [4-1:0] node8212;
	wire [4-1:0] node8213;
	wire [4-1:0] node8217;
	wire [4-1:0] node8218;
	wire [4-1:0] node8219;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8226;
	wire [4-1:0] node8227;
	wire [4-1:0] node8230;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8236;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8247;
	wire [4-1:0] node8250;
	wire [4-1:0] node8251;
	wire [4-1:0] node8252;
	wire [4-1:0] node8253;
	wire [4-1:0] node8255;
	wire [4-1:0] node8258;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8265;
	wire [4-1:0] node8268;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8275;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8282;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8289;
	wire [4-1:0] node8292;
	wire [4-1:0] node8293;
	wire [4-1:0] node8294;
	wire [4-1:0] node8297;
	wire [4-1:0] node8299;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8308;
	wire [4-1:0] node8312;
	wire [4-1:0] node8313;
	wire [4-1:0] node8315;
	wire [4-1:0] node8318;
	wire [4-1:0] node8321;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8327;
	wire [4-1:0] node8328;
	wire [4-1:0] node8332;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8336;
	wire [4-1:0] node8339;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8352;
	wire [4-1:0] node8354;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8362;
	wire [4-1:0] node8367;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8380;
	wire [4-1:0] node8381;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8386;
	wire [4-1:0] node8390;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8396;
	wire [4-1:0] node8398;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8404;
	wire [4-1:0] node8408;
	wire [4-1:0] node8410;
	wire [4-1:0] node8411;
	wire [4-1:0] node8412;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8419;
	wire [4-1:0] node8422;
	wire [4-1:0] node8424;
	wire [4-1:0] node8427;
	wire [4-1:0] node8428;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8432;
	wire [4-1:0] node8435;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8440;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8450;
	wire [4-1:0] node8452;
	wire [4-1:0] node8455;
	wire [4-1:0] node8459;
	wire [4-1:0] node8460;
	wire [4-1:0] node8461;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8474;
	wire [4-1:0] node8475;
	wire [4-1:0] node8476;
	wire [4-1:0] node8477;
	wire [4-1:0] node8478;
	wire [4-1:0] node8479;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8490;
	wire [4-1:0] node8494;
	wire [4-1:0] node8496;
	wire [4-1:0] node8498;
	wire [4-1:0] node8500;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8507;
	wire [4-1:0] node8509;
	wire [4-1:0] node8512;
	wire [4-1:0] node8513;
	wire [4-1:0] node8515;
	wire [4-1:0] node8520;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8524;
	wire [4-1:0] node8525;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8540;
	wire [4-1:0] node8541;
	wire [4-1:0] node8543;
	wire [4-1:0] node8547;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8552;
	wire [4-1:0] node8554;
	wire [4-1:0] node8555;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8565;
	wire [4-1:0] node8567;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8573;
	wire [4-1:0] node8577;
	wire [4-1:0] node8581;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8587;
	wire [4-1:0] node8589;
	wire [4-1:0] node8593;
	wire [4-1:0] node8594;
	wire [4-1:0] node8595;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8602;
	wire [4-1:0] node8605;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8611;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8614;
	wire [4-1:0] node8616;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8627;
	wire [4-1:0] node8630;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8637;
	wire [4-1:0] node8639;
	wire [4-1:0] node8642;
	wire [4-1:0] node8643;
	wire [4-1:0] node8646;
	wire [4-1:0] node8648;
	wire [4-1:0] node8651;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8661;
	wire [4-1:0] node8663;
	wire [4-1:0] node8665;
	wire [4-1:0] node8668;
	wire [4-1:0] node8670;
	wire [4-1:0] node8672;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8677;
	wire [4-1:0] node8680;
	wire [4-1:0] node8681;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8689;
	wire [4-1:0] node8694;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8699;
	wire [4-1:0] node8703;
	wire [4-1:0] node8706;
	wire [4-1:0] node8707;
	wire [4-1:0] node8708;
	wire [4-1:0] node8709;
	wire [4-1:0] node8712;
	wire [4-1:0] node8715;
	wire [4-1:0] node8716;
	wire [4-1:0] node8720;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8727;
	wire [4-1:0] node8728;
	wire [4-1:0] node8729;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8736;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8741;
	wire [4-1:0] node8744;
	wire [4-1:0] node8748;
	wire [4-1:0] node8749;
	wire [4-1:0] node8750;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8756;
	wire [4-1:0] node8757;
	wire [4-1:0] node8761;
	wire [4-1:0] node8762;
	wire [4-1:0] node8763;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8770;
	wire [4-1:0] node8774;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8778;
	wire [4-1:0] node8781;
	wire [4-1:0] node8784;
	wire [4-1:0] node8787;
	wire [4-1:0] node8789;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8798;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8811;
	wire [4-1:0] node8813;
	wire [4-1:0] node8815;
	wire [4-1:0] node8819;
	wire [4-1:0] node8820;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8823;
	wire [4-1:0] node8826;
	wire [4-1:0] node8829;
	wire [4-1:0] node8830;
	wire [4-1:0] node8832;
	wire [4-1:0] node8836;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8850;
	wire [4-1:0] node8853;
	wire [4-1:0] node8856;
	wire [4-1:0] node8857;
	wire [4-1:0] node8860;
	wire [4-1:0] node8861;
	wire [4-1:0] node8865;
	wire [4-1:0] node8866;
	wire [4-1:0] node8868;
	wire [4-1:0] node8871;
	wire [4-1:0] node8873;
	wire [4-1:0] node8876;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8880;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8885;
	wire [4-1:0] node8888;
	wire [4-1:0] node8890;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8898;
	wire [4-1:0] node8899;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8907;
	wire [4-1:0] node8909;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8916;
	wire [4-1:0] node8920;
	wire [4-1:0] node8921;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8931;
	wire [4-1:0] node8932;
	wire [4-1:0] node8933;
	wire [4-1:0] node8934;
	wire [4-1:0] node8935;
	wire [4-1:0] node8936;
	wire [4-1:0] node8940;
	wire [4-1:0] node8941;
	wire [4-1:0] node8942;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8958;
	wire [4-1:0] node8960;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8977;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8985;
	wire [4-1:0] node8986;
	wire [4-1:0] node8987;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8995;
	wire [4-1:0] node8996;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9007;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9015;
	wire [4-1:0] node9018;
	wire [4-1:0] node9020;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9027;
	wire [4-1:0] node9028;
	wire [4-1:0] node9029;
	wire [4-1:0] node9034;
	wire [4-1:0] node9036;
	wire [4-1:0] node9037;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9045;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9050;
	wire [4-1:0] node9051;
	wire [4-1:0] node9052;
	wire [4-1:0] node9054;
	wire [4-1:0] node9058;
	wire [4-1:0] node9059;
	wire [4-1:0] node9060;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9068;
	wire [4-1:0] node9070;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9078;
	wire [4-1:0] node9079;
	wire [4-1:0] node9080;
	wire [4-1:0] node9081;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9089;
	wire [4-1:0] node9092;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9098;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9106;
	wire [4-1:0] node9109;
	wire [4-1:0] node9110;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9113;
	wire [4-1:0] node9115;
	wire [4-1:0] node9116;
	wire [4-1:0] node9120;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9129;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9138;
	wire [4-1:0] node9142;
	wire [4-1:0] node9144;
	wire [4-1:0] node9147;
	wire [4-1:0] node9149;
	wire [4-1:0] node9150;
	wire [4-1:0] node9154;
	wire [4-1:0] node9155;
	wire [4-1:0] node9156;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9163;
	wire [4-1:0] node9165;
	wire [4-1:0] node9168;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9175;
	wire [4-1:0] node9177;
	wire [4-1:0] node9179;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9184;
	wire [4-1:0] node9185;
	wire [4-1:0] node9189;
	wire [4-1:0] node9191;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9199;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9207;
	wire [4-1:0] node9210;
	wire [4-1:0] node9211;
	wire [4-1:0] node9214;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9221;
	wire [4-1:0] node9222;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9235;
	wire [4-1:0] node9237;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9242;
	wire [4-1:0] node9244;
	wire [4-1:0] node9247;
	wire [4-1:0] node9248;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9255;
	wire [4-1:0] node9256;
	wire [4-1:0] node9260;
	wire [4-1:0] node9262;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9268;
	wire [4-1:0] node9272;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9275;
	wire [4-1:0] node9279;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9287;
	wire [4-1:0] node9288;
	wire [4-1:0] node9289;
	wire [4-1:0] node9292;
	wire [4-1:0] node9295;
	wire [4-1:0] node9297;
	wire [4-1:0] node9300;
	wire [4-1:0] node9301;
	wire [4-1:0] node9302;
	wire [4-1:0] node9303;
	wire [4-1:0] node9304;
	wire [4-1:0] node9305;
	wire [4-1:0] node9306;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9310;
	wire [4-1:0] node9314;
	wire [4-1:0] node9317;
	wire [4-1:0] node9318;
	wire [4-1:0] node9322;
	wire [4-1:0] node9323;
	wire [4-1:0] node9324;
	wire [4-1:0] node9326;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9334;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9342;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9364;
	wire [4-1:0] node9365;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9372;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9384;
	wire [4-1:0] node9387;
	wire [4-1:0] node9388;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9397;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9407;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9414;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9425;
	wire [4-1:0] node9428;
	wire [4-1:0] node9429;
	wire [4-1:0] node9433;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9439;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9447;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9456;
	wire [4-1:0] node9457;
	wire [4-1:0] node9458;
	wire [4-1:0] node9460;
	wire [4-1:0] node9463;
	wire [4-1:0] node9465;
	wire [4-1:0] node9468;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9474;
	wire [4-1:0] node9477;
	wire [4-1:0] node9479;
	wire [4-1:0] node9480;
	wire [4-1:0] node9484;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9491;
	wire [4-1:0] node9494;
	wire [4-1:0] node9497;
	wire [4-1:0] node9498;
	wire [4-1:0] node9499;
	wire [4-1:0] node9501;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9508;
	wire [4-1:0] node9511;
	wire [4-1:0] node9512;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9520;
	wire [4-1:0] node9521;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9534;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9546;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9553;
	wire [4-1:0] node9555;
	wire [4-1:0] node9558;
	wire [4-1:0] node9560;
	wire [4-1:0] node9561;
	wire [4-1:0] node9563;
	wire [4-1:0] node9565;
	wire [4-1:0] node9568;
	wire [4-1:0] node9570;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9582;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9589;
	wire [4-1:0] node9591;
	wire [4-1:0] node9593;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9600;
	wire [4-1:0] node9601;
	wire [4-1:0] node9603;
	wire [4-1:0] node9607;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9614;
	wire [4-1:0] node9616;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9632;
	wire [4-1:0] node9635;
	wire [4-1:0] node9636;
	wire [4-1:0] node9637;
	wire [4-1:0] node9641;
	wire [4-1:0] node9643;
	wire [4-1:0] node9646;
	wire [4-1:0] node9647;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9655;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9664;
	wire [4-1:0] node9666;
	wire [4-1:0] node9669;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9681;
	wire [4-1:0] node9682;
	wire [4-1:0] node9683;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9690;
	wire [4-1:0] node9692;
	wire [4-1:0] node9697;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9702;
	wire [4-1:0] node9703;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9711;
	wire [4-1:0] node9714;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9723;
	wire [4-1:0] node9726;
	wire [4-1:0] node9729;
	wire [4-1:0] node9730;
	wire [4-1:0] node9733;
	wire [4-1:0] node9735;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9741;
	wire [4-1:0] node9744;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9749;
	wire [4-1:0] node9753;
	wire [4-1:0] node9754;
	wire [4-1:0] node9755;
	wire [4-1:0] node9758;
	wire [4-1:0] node9760;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9765;
	wire [4-1:0] node9768;
	wire [4-1:0] node9769;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9777;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9787;
	wire [4-1:0] node9789;
	wire [4-1:0] node9792;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9804;
	wire [4-1:0] node9805;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9813;
	wire [4-1:0] node9816;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9820;
	wire [4-1:0] node9824;
	wire [4-1:0] node9826;
	wire [4-1:0] node9827;
	wire [4-1:0] node9831;
	wire [4-1:0] node9833;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9844;
	wire [4-1:0] node9845;
	wire [4-1:0] node9846;
	wire [4-1:0] node9851;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9856;
	wire [4-1:0] node9859;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9868;
	wire [4-1:0] node9869;
	wire [4-1:0] node9872;
	wire [4-1:0] node9874;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9884;
	wire [4-1:0] node9887;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9893;
	wire [4-1:0] node9896;
	wire [4-1:0] node9897;
	wire [4-1:0] node9898;
	wire [4-1:0] node9899;
	wire [4-1:0] node9900;
	wire [4-1:0] node9901;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9907;
	wire [4-1:0] node9910;
	wire [4-1:0] node9913;
	wire [4-1:0] node9914;
	wire [4-1:0] node9917;
	wire [4-1:0] node9919;
	wire [4-1:0] node9922;
	wire [4-1:0] node9923;
	wire [4-1:0] node9925;
	wire [4-1:0] node9926;
	wire [4-1:0] node9930;
	wire [4-1:0] node9933;
	wire [4-1:0] node9934;
	wire [4-1:0] node9935;
	wire [4-1:0] node9936;
	wire [4-1:0] node9937;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9956;
	wire [4-1:0] node9957;
	wire [4-1:0] node9958;
	wire [4-1:0] node9959;
	wire [4-1:0] node9960;
	wire [4-1:0] node9961;
	wire [4-1:0] node9966;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9973;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9982;
	wire [4-1:0] node9985;
	wire [4-1:0] node9988;
	wire [4-1:0] node9990;
	wire [4-1:0] node9995;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10002;
	wire [4-1:0] node10004;
	wire [4-1:0] node10008;
	wire [4-1:0] node10011;
	wire [4-1:0] node10013;
	wire [4-1:0] node10017;
	wire [4-1:0] node10018;
	wire [4-1:0] node10019;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10025;
	wire [4-1:0] node10027;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10033;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10042;
	wire [4-1:0] node10043;
	wire [4-1:0] node10046;
	wire [4-1:0] node10049;
	wire [4-1:0] node10050;
	wire [4-1:0] node10052;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10056;
	wire [4-1:0] node10061;
	wire [4-1:0] node10062;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10070;
	wire [4-1:0] node10071;
	wire [4-1:0] node10072;
	wire [4-1:0] node10073;
	wire [4-1:0] node10074;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10080;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10084;
	wire [4-1:0] node10087;
	wire [4-1:0] node10090;
	wire [4-1:0] node10092;
	wire [4-1:0] node10094;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10104;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10114;
	wire [4-1:0] node10116;
	wire [4-1:0] node10119;
	wire [4-1:0] node10120;
	wire [4-1:0] node10122;
	wire [4-1:0] node10126;
	wire [4-1:0] node10128;
	wire [4-1:0] node10130;
	wire [4-1:0] node10132;
	wire [4-1:0] node10134;
	wire [4-1:0] node10137;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10146;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10152;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10159;
	wire [4-1:0] node10160;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10169;
	wire [4-1:0] node10170;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10182;
	wire [4-1:0] node10184;
	wire [4-1:0] node10187;
	wire [4-1:0] node10189;
	wire [4-1:0] node10192;
	wire [4-1:0] node10193;
	wire [4-1:0] node10196;
	wire [4-1:0] node10197;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10208;
	wire [4-1:0] node10209;
	wire [4-1:0] node10212;
	wire [4-1:0] node10215;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10219;
	wire [4-1:0] node10223;
	wire [4-1:0] node10224;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10234;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10240;
	wire [4-1:0] node10244;
	wire [4-1:0] node10245;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10251;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10261;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10267;
	wire [4-1:0] node10268;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10276;
	wire [4-1:0] node10278;
	wire [4-1:0] node10280;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10286;
	wire [4-1:0] node10288;
	wire [4-1:0] node10291;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10301;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10305;
	wire [4-1:0] node10307;
	wire [4-1:0] node10310;
	wire [4-1:0] node10311;
	wire [4-1:0] node10312;
	wire [4-1:0] node10316;
	wire [4-1:0] node10318;
	wire [4-1:0] node10320;
	wire [4-1:0] node10323;
	wire [4-1:0] node10324;
	wire [4-1:0] node10325;
	wire [4-1:0] node10327;
	wire [4-1:0] node10330;
	wire [4-1:0] node10333;
	wire [4-1:0] node10334;
	wire [4-1:0] node10337;
	wire [4-1:0] node10338;
	wire [4-1:0] node10340;
	wire [4-1:0] node10341;
	wire [4-1:0] node10346;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10350;
	wire [4-1:0] node10351;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10358;
	wire [4-1:0] node10362;
	wire [4-1:0] node10365;
	wire [4-1:0] node10366;
	wire [4-1:0] node10368;
	wire [4-1:0] node10372;
	wire [4-1:0] node10373;
	wire [4-1:0] node10374;
	wire [4-1:0] node10376;
	wire [4-1:0] node10380;
	wire [4-1:0] node10383;
	wire [4-1:0] node10385;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10389;
	wire [4-1:0] node10390;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10395;
	wire [4-1:0] node10399;
	wire [4-1:0] node10401;
	wire [4-1:0] node10403;
	wire [4-1:0] node10404;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10410;
	wire [4-1:0] node10411;
	wire [4-1:0] node10412;
	wire [4-1:0] node10414;
	wire [4-1:0] node10418;
	wire [4-1:0] node10419;
	wire [4-1:0] node10423;
	wire [4-1:0] node10424;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10430;
	wire [4-1:0] node10433;
	wire [4-1:0] node10436;
	wire [4-1:0] node10438;
	wire [4-1:0] node10440;
	wire [4-1:0] node10441;
	wire [4-1:0] node10444;
	wire [4-1:0] node10447;
	wire [4-1:0] node10448;
	wire [4-1:0] node10449;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10459;
	wire [4-1:0] node10460;
	wire [4-1:0] node10464;
	wire [4-1:0] node10465;
	wire [4-1:0] node10467;
	wire [4-1:0] node10468;
	wire [4-1:0] node10472;
	wire [4-1:0] node10473;
	wire [4-1:0] node10474;
	wire [4-1:0] node10476;
	wire [4-1:0] node10479;
	wire [4-1:0] node10482;
	wire [4-1:0] node10484;
	wire [4-1:0] node10487;
	wire [4-1:0] node10488;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10498;
	wire [4-1:0] node10502;
	wire [4-1:0] node10503;
	wire [4-1:0] node10504;
	wire [4-1:0] node10508;
	wire [4-1:0] node10509;
	wire [4-1:0] node10512;
	wire [4-1:0] node10515;
	wire [4-1:0] node10516;
	wire [4-1:0] node10518;
	wire [4-1:0] node10520;
	wire [4-1:0] node10523;
	wire [4-1:0] node10524;
	wire [4-1:0] node10529;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10534;
	wire [4-1:0] node10535;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10540;
	wire [4-1:0] node10543;
	wire [4-1:0] node10546;
	wire [4-1:0] node10548;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10558;
	wire [4-1:0] node10560;
	wire [4-1:0] node10563;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10569;
	wire [4-1:0] node10571;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10577;
	wire [4-1:0] node10578;
	wire [4-1:0] node10582;
	wire [4-1:0] node10583;
	wire [4-1:0] node10586;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10598;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10605;
	wire [4-1:0] node10608;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10615;
	wire [4-1:0] node10619;
	wire [4-1:0] node10620;
	wire [4-1:0] node10621;
	wire [4-1:0] node10622;
	wire [4-1:0] node10624;
	wire [4-1:0] node10627;
	wire [4-1:0] node10630;
	wire [4-1:0] node10631;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10644;
	wire [4-1:0] node10645;
	wire [4-1:0] node10647;
	wire [4-1:0] node10650;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10657;
	wire [4-1:0] node10660;
	wire [4-1:0] node10662;
	wire [4-1:0] node10665;
	wire [4-1:0] node10666;
	wire [4-1:0] node10669;
	wire [4-1:0] node10671;
	wire [4-1:0] node10674;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10681;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10686;
	wire [4-1:0] node10689;
	wire [4-1:0] node10692;
	wire [4-1:0] node10694;
	wire [4-1:0] node10695;
	wire [4-1:0] node10699;
	wire [4-1:0] node10700;
	wire [4-1:0] node10702;
	wire [4-1:0] node10704;
	wire [4-1:0] node10707;
	wire [4-1:0] node10708;
	wire [4-1:0] node10709;
	wire [4-1:0] node10710;
	wire [4-1:0] node10714;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10724;
	wire [4-1:0] node10725;
	wire [4-1:0] node10730;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10736;
	wire [4-1:0] node10739;
	wire [4-1:0] node10740;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10746;
	wire [4-1:0] node10749;
	wire [4-1:0] node10751;
	wire [4-1:0] node10754;
	wire [4-1:0] node10755;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10760;
	wire [4-1:0] node10763;
	wire [4-1:0] node10764;
	wire [4-1:0] node10766;
	wire [4-1:0] node10769;
	wire [4-1:0] node10772;
	wire [4-1:0] node10774;
	wire [4-1:0] node10775;
	wire [4-1:0] node10777;
	wire [4-1:0] node10780;
	wire [4-1:0] node10781;
	wire [4-1:0] node10784;
	wire [4-1:0] node10785;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10796;
	wire [4-1:0] node10797;
	wire [4-1:0] node10800;
	wire [4-1:0] node10803;
	wire [4-1:0] node10805;
	wire [4-1:0] node10807;
	wire [4-1:0] node10810;
	wire [4-1:0] node10811;
	wire [4-1:0] node10815;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10819;
	wire [4-1:0] node10822;
	wire [4-1:0] node10824;
	wire [4-1:0] node10826;
	wire [4-1:0] node10829;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10834;
	wire [4-1:0] node10837;
	wire [4-1:0] node10840;
	wire [4-1:0] node10841;
	wire [4-1:0] node10842;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10848;
	wire [4-1:0] node10850;
	wire [4-1:0] node10854;
	wire [4-1:0] node10855;
	wire [4-1:0] node10858;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10867;
	wire [4-1:0] node10871;
	wire [4-1:0] node10872;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10880;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10883;
	wire [4-1:0] node10886;
	wire [4-1:0] node10888;
	wire [4-1:0] node10889;
	wire [4-1:0] node10892;
	wire [4-1:0] node10895;
	wire [4-1:0] node10897;
	wire [4-1:0] node10899;
	wire [4-1:0] node10902;
	wire [4-1:0] node10903;
	wire [4-1:0] node10905;
	wire [4-1:0] node10908;
	wire [4-1:0] node10910;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10915;
	wire [4-1:0] node10916;
	wire [4-1:0] node10918;
	wire [4-1:0] node10919;
	wire [4-1:0] node10923;
	wire [4-1:0] node10924;
	wire [4-1:0] node10926;
	wire [4-1:0] node10929;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10940;
	wire [4-1:0] node10941;
	wire [4-1:0] node10943;
	wire [4-1:0] node10944;
	wire [4-1:0] node10948;
	wire [4-1:0] node10951;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10954;
	wire [4-1:0] node10955;
	wire [4-1:0] node10959;
	wire [4-1:0] node10961;
	wire [4-1:0] node10964;
	wire [4-1:0] node10966;
	wire [4-1:0] node10968;
	wire [4-1:0] node10970;
	wire [4-1:0] node10973;
	wire [4-1:0] node10974;
	wire [4-1:0] node10976;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10984;
	wire [4-1:0] node10985;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10989;
	wire [4-1:0] node10990;
	wire [4-1:0] node10991;
	wire [4-1:0] node10996;
	wire [4-1:0] node10997;
	wire [4-1:0] node10998;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11003;
	wire [4-1:0] node11005;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11011;
	wire [4-1:0] node11012;
	wire [4-1:0] node11017;
	wire [4-1:0] node11019;
	wire [4-1:0] node11020;
	wire [4-1:0] node11024;
	wire [4-1:0] node11026;
	wire [4-1:0] node11028;
	wire [4-1:0] node11029;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11035;
	wire [4-1:0] node11036;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11047;
	wire [4-1:0] node11048;
	wire [4-1:0] node11050;
	wire [4-1:0] node11052;
	wire [4-1:0] node11055;
	wire [4-1:0] node11058;
	wire [4-1:0] node11059;
	wire [4-1:0] node11060;
	wire [4-1:0] node11063;
	wire [4-1:0] node11064;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11071;
	wire [4-1:0] node11074;
	wire [4-1:0] node11075;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11082;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11087;
	wire [4-1:0] node11088;
	wire [4-1:0] node11089;
	wire [4-1:0] node11093;
	wire [4-1:0] node11096;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11102;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11114;
	wire [4-1:0] node11115;
	wire [4-1:0] node11118;
	wire [4-1:0] node11121;
	wire [4-1:0] node11122;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11131;
	wire [4-1:0] node11132;
	wire [4-1:0] node11133;
	wire [4-1:0] node11134;
	wire [4-1:0] node11135;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11140;
	wire [4-1:0] node11142;
	wire [4-1:0] node11145;
	wire [4-1:0] node11146;
	wire [4-1:0] node11148;
	wire [4-1:0] node11152;
	wire [4-1:0] node11154;
	wire [4-1:0] node11156;
	wire [4-1:0] node11159;
	wire [4-1:0] node11160;
	wire [4-1:0] node11162;
	wire [4-1:0] node11164;
	wire [4-1:0] node11167;
	wire [4-1:0] node11168;
	wire [4-1:0] node11171;
	wire [4-1:0] node11172;
	wire [4-1:0] node11175;
	wire [4-1:0] node11176;
	wire [4-1:0] node11180;
	wire [4-1:0] node11181;
	wire [4-1:0] node11182;
	wire [4-1:0] node11183;
	wire [4-1:0] node11184;
	wire [4-1:0] node11188;
	wire [4-1:0] node11190;
	wire [4-1:0] node11193;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11199;
	wire [4-1:0] node11201;
	wire [4-1:0] node11205;
	wire [4-1:0] node11206;
	wire [4-1:0] node11207;
	wire [4-1:0] node11208;
	wire [4-1:0] node11209;
	wire [4-1:0] node11211;
	wire [4-1:0] node11213;
	wire [4-1:0] node11216;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11221;
	wire [4-1:0] node11223;
	wire [4-1:0] node11227;
	wire [4-1:0] node11228;
	wire [4-1:0] node11232;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11238;
	wire [4-1:0] node11240;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11248;
	wire [4-1:0] node11250;
	wire [4-1:0] node11252;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11259;
	wire [4-1:0] node11261;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11266;
	wire [4-1:0] node11267;
	wire [4-1:0] node11272;
	wire [4-1:0] node11273;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11285;
	wire [4-1:0] node11286;
	wire [4-1:0] node11289;
	wire [4-1:0] node11292;
	wire [4-1:0] node11293;
	wire [4-1:0] node11296;
	wire [4-1:0] node11299;
	wire [4-1:0] node11300;
	wire [4-1:0] node11301;
	wire [4-1:0] node11306;
	wire [4-1:0] node11307;
	wire [4-1:0] node11308;
	wire [4-1:0] node11309;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11312;
	wire [4-1:0] node11315;
	wire [4-1:0] node11317;
	wire [4-1:0] node11320;
	wire [4-1:0] node11323;
	wire [4-1:0] node11324;
	wire [4-1:0] node11325;
	wire [4-1:0] node11326;
	wire [4-1:0] node11331;
	wire [4-1:0] node11334;
	wire [4-1:0] node11335;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11345;
	wire [4-1:0] node11347;
	wire [4-1:0] node11349;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11355;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11363;
	wire [4-1:0] node11365;
	wire [4-1:0] node11368;
	wire [4-1:0] node11370;
	wire [4-1:0] node11373;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11376;
	wire [4-1:0] node11379;
	wire [4-1:0] node11380;
	wire [4-1:0] node11383;
	wire [4-1:0] node11385;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11395;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11401;
	wire [4-1:0] node11402;
	wire [4-1:0] node11405;
	wire [4-1:0] node11406;
	wire [4-1:0] node11410;
	wire [4-1:0] node11411;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11420;
	wire [4-1:0] node11421;
	wire [4-1:0] node11425;
	wire [4-1:0] node11427;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11437;
	wire [4-1:0] node11439;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11448;
	wire [4-1:0] node11449;
	wire [4-1:0] node11452;
	wire [4-1:0] node11454;
	wire [4-1:0] node11457;
	wire [4-1:0] node11458;
	wire [4-1:0] node11460;
	wire [4-1:0] node11461;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11468;
	wire [4-1:0] node11472;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11483;
	wire [4-1:0] node11485;
	wire [4-1:0] node11487;
	wire [4-1:0] node11490;
	wire [4-1:0] node11491;
	wire [4-1:0] node11495;
	wire [4-1:0] node11496;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11501;
	wire [4-1:0] node11503;
	wire [4-1:0] node11504;
	wire [4-1:0] node11508;
	wire [4-1:0] node11509;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11517;
	wire [4-1:0] node11518;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11523;
	wire [4-1:0] node11528;
	wire [4-1:0] node11529;
	wire [4-1:0] node11530;
	wire [4-1:0] node11532;
	wire [4-1:0] node11536;
	wire [4-1:0] node11537;
	wire [4-1:0] node11538;
	wire [4-1:0] node11540;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11549;
	wire [4-1:0] node11550;
	wire [4-1:0] node11551;
	wire [4-1:0] node11553;
	wire [4-1:0] node11554;
	wire [4-1:0] node11557;
	wire [4-1:0] node11560;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11565;
	wire [4-1:0] node11566;
	wire [4-1:0] node11569;
	wire [4-1:0] node11570;
	wire [4-1:0] node11574;
	wire [4-1:0] node11575;
	wire [4-1:0] node11579;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11583;
	wire [4-1:0] node11584;
	wire [4-1:0] node11587;
	wire [4-1:0] node11590;
	wire [4-1:0] node11591;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11599;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11603;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11609;
	wire [4-1:0] node11613;
	wire [4-1:0] node11615;
	wire [4-1:0] node11616;
	wire [4-1:0] node11620;
	wire [4-1:0] node11621;
	wire [4-1:0] node11622;
	wire [4-1:0] node11623;
	wire [4-1:0] node11624;
	wire [4-1:0] node11627;
	wire [4-1:0] node11629;
	wire [4-1:0] node11632;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11637;
	wire [4-1:0] node11639;
	wire [4-1:0] node11642;
	wire [4-1:0] node11645;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11649;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11656;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11669;
	wire [4-1:0] node11670;
	wire [4-1:0] node11672;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11680;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11686;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11696;
	wire [4-1:0] node11697;
	wire [4-1:0] node11701;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11704;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11707;
	wire [4-1:0] node11710;
	wire [4-1:0] node11712;
	wire [4-1:0] node11715;
	wire [4-1:0] node11718;
	wire [4-1:0] node11719;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11726;
	wire [4-1:0] node11729;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11733;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11740;
	wire [4-1:0] node11742;
	wire [4-1:0] node11745;
	wire [4-1:0] node11747;
	wire [4-1:0] node11748;
	wire [4-1:0] node11749;
	wire [4-1:0] node11753;
	wire [4-1:0] node11754;
	wire [4-1:0] node11755;
	wire [4-1:0] node11760;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11764;
	wire [4-1:0] node11765;
	wire [4-1:0] node11767;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11773;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11779;
	wire [4-1:0] node11783;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11789;
	wire [4-1:0] node11791;
	wire [4-1:0] node11794;
	wire [4-1:0] node11795;
	wire [4-1:0] node11796;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11803;
	wire [4-1:0] node11804;
	wire [4-1:0] node11805;
	wire [4-1:0] node11807;
	wire [4-1:0] node11809;
	wire [4-1:0] node11812;
	wire [4-1:0] node11813;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11821;
	wire [4-1:0] node11822;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11829;
	wire [4-1:0] node11830;
	wire [4-1:0] node11832;
	wire [4-1:0] node11835;
	wire [4-1:0] node11837;
	wire [4-1:0] node11840;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11845;
	wire [4-1:0] node11846;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11853;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11862;
	wire [4-1:0] node11863;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11866;
	wire [4-1:0] node11868;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11872;
	wire [4-1:0] node11873;
	wire [4-1:0] node11875;
	wire [4-1:0] node11878;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11886;
	wire [4-1:0] node11887;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11891;
	wire [4-1:0] node11893;
	wire [4-1:0] node11896;
	wire [4-1:0] node11898;
	wire [4-1:0] node11900;
	wire [4-1:0] node11901;
	wire [4-1:0] node11905;
	wire [4-1:0] node11906;
	wire [4-1:0] node11907;
	wire [4-1:0] node11909;
	wire [4-1:0] node11912;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11920;
	wire [4-1:0] node11921;
	wire [4-1:0] node11924;
	wire [4-1:0] node11926;
	wire [4-1:0] node11928;
	wire [4-1:0] node11931;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11936;
	wire [4-1:0] node11938;
	wire [4-1:0] node11940;
	wire [4-1:0] node11943;
	wire [4-1:0] node11945;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11950;
	wire [4-1:0] node11953;
	wire [4-1:0] node11954;
	wire [4-1:0] node11958;
	wire [4-1:0] node11959;
	wire [4-1:0] node11962;
	wire [4-1:0] node11963;
	wire [4-1:0] node11967;
	wire [4-1:0] node11968;
	wire [4-1:0] node11969;
	wire [4-1:0] node11970;
	wire [4-1:0] node11972;
	wire [4-1:0] node11976;
	wire [4-1:0] node11977;
	wire [4-1:0] node11981;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11992;
	wire [4-1:0] node11993;
	wire [4-1:0] node11994;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node12000;
	wire [4-1:0] node12001;
	wire [4-1:0] node12005;
	wire [4-1:0] node12006;
	wire [4-1:0] node12008;
	wire [4-1:0] node12011;
	wire [4-1:0] node12014;
	wire [4-1:0] node12015;
	wire [4-1:0] node12017;
	wire [4-1:0] node12018;
	wire [4-1:0] node12022;
	wire [4-1:0] node12023;
	wire [4-1:0] node12025;
	wire [4-1:0] node12027;
	wire [4-1:0] node12028;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12035;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12043;
	wire [4-1:0] node12044;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12057;
	wire [4-1:0] node12058;
	wire [4-1:0] node12062;
	wire [4-1:0] node12063;
	wire [4-1:0] node12064;
	wire [4-1:0] node12066;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12075;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12089;
	wire [4-1:0] node12091;
	wire [4-1:0] node12094;
	wire [4-1:0] node12095;
	wire [4-1:0] node12097;
	wire [4-1:0] node12099;
	wire [4-1:0] node12103;
	wire [4-1:0] node12104;
	wire [4-1:0] node12105;
	wire [4-1:0] node12107;
	wire [4-1:0] node12110;
	wire [4-1:0] node12111;
	wire [4-1:0] node12113;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12119;
	wire [4-1:0] node12120;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12130;
	wire [4-1:0] node12134;
	wire [4-1:0] node12136;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12142;
	wire [4-1:0] node12145;
	wire [4-1:0] node12146;
	wire [4-1:0] node12149;
	wire [4-1:0] node12150;
	wire [4-1:0] node12153;
	wire [4-1:0] node12156;
	wire [4-1:0] node12158;
	wire [4-1:0] node12160;
	wire [4-1:0] node12162;
	wire [4-1:0] node12163;
	wire [4-1:0] node12167;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12170;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12173;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12180;
	wire [4-1:0] node12182;
	wire [4-1:0] node12184;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12191;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12198;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12210;
	wire [4-1:0] node12211;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12217;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12224;
	wire [4-1:0] node12227;
	wire [4-1:0] node12228;
	wire [4-1:0] node12230;
	wire [4-1:0] node12233;
	wire [4-1:0] node12234;
	wire [4-1:0] node12237;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12244;
	wire [4-1:0] node12246;
	wire [4-1:0] node12249;
	wire [4-1:0] node12252;
	wire [4-1:0] node12253;
	wire [4-1:0] node12255;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12263;
	wire [4-1:0] node12266;
	wire [4-1:0] node12269;
	wire [4-1:0] node12270;
	wire [4-1:0] node12271;
	wire [4-1:0] node12272;
	wire [4-1:0] node12273;
	wire [4-1:0] node12276;
	wire [4-1:0] node12278;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12284;
	wire [4-1:0] node12285;
	wire [4-1:0] node12286;
	wire [4-1:0] node12290;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12298;
	wire [4-1:0] node12299;
	wire [4-1:0] node12301;
	wire [4-1:0] node12304;
	wire [4-1:0] node12306;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12313;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12323;
	wire [4-1:0] node12324;
	wire [4-1:0] node12328;
	wire [4-1:0] node12331;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12334;
	wire [4-1:0] node12336;
	wire [4-1:0] node12339;
	wire [4-1:0] node12342;
	wire [4-1:0] node12343;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12349;
	wire [4-1:0] node12350;
	wire [4-1:0] node12354;
	wire [4-1:0] node12357;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12369;
	wire [4-1:0] node12372;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12375;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12387;
	wire [4-1:0] node12388;
	wire [4-1:0] node12392;
	wire [4-1:0] node12393;
	wire [4-1:0] node12396;
	wire [4-1:0] node12399;
	wire [4-1:0] node12400;
	wire [4-1:0] node12401;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12412;
	wire [4-1:0] node12414;
	wire [4-1:0] node12415;
	wire [4-1:0] node12419;
	wire [4-1:0] node12420;
	wire [4-1:0] node12421;
	wire [4-1:0] node12424;
	wire [4-1:0] node12426;
	wire [4-1:0] node12427;
	wire [4-1:0] node12431;
	wire [4-1:0] node12432;
	wire [4-1:0] node12433;
	wire [4-1:0] node12438;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12446;
	wire [4-1:0] node12449;
	wire [4-1:0] node12450;
	wire [4-1:0] node12453;
	wire [4-1:0] node12455;
	wire [4-1:0] node12458;
	wire [4-1:0] node12459;
	wire [4-1:0] node12460;
	wire [4-1:0] node12462;
	wire [4-1:0] node12465;
	wire [4-1:0] node12468;
	wire [4-1:0] node12469;
	wire [4-1:0] node12472;
	wire [4-1:0] node12474;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12480;
	wire [4-1:0] node12483;
	wire [4-1:0] node12484;
	wire [4-1:0] node12486;
	wire [4-1:0] node12490;
	wire [4-1:0] node12491;
	wire [4-1:0] node12492;
	wire [4-1:0] node12493;
	wire [4-1:0] node12495;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12504;
	wire [4-1:0] node12507;
	wire [4-1:0] node12510;
	wire [4-1:0] node12511;
	wire [4-1:0] node12512;
	wire [4-1:0] node12516;
	wire [4-1:0] node12517;
	wire [4-1:0] node12518;
	wire [4-1:0] node12522;
	wire [4-1:0] node12524;
	wire [4-1:0] node12527;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12531;
	wire [4-1:0] node12532;
	wire [4-1:0] node12534;
	wire [4-1:0] node12535;
	wire [4-1:0] node12538;
	wire [4-1:0] node12541;
	wire [4-1:0] node12542;
	wire [4-1:0] node12544;
	wire [4-1:0] node12546;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12554;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12557;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12564;
	wire [4-1:0] node12568;
	wire [4-1:0] node12569;
	wire [4-1:0] node12570;
	wire [4-1:0] node12571;
	wire [4-1:0] node12575;
	wire [4-1:0] node12578;
	wire [4-1:0] node12579;
	wire [4-1:0] node12583;
	wire [4-1:0] node12584;
	wire [4-1:0] node12585;
	wire [4-1:0] node12587;
	wire [4-1:0] node12589;
	wire [4-1:0] node12592;
	wire [4-1:0] node12593;
	wire [4-1:0] node12595;
	wire [4-1:0] node12596;
	wire [4-1:0] node12600;
	wire [4-1:0] node12601;
	wire [4-1:0] node12602;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12611;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12615;
	wire [4-1:0] node12618;
	wire [4-1:0] node12620;
	wire [4-1:0] node12623;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12628;
	wire [4-1:0] node12629;
	wire [4-1:0] node12634;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12637;
	wire [4-1:0] node12639;
	wire [4-1:0] node12641;
	wire [4-1:0] node12644;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12647;
	wire [4-1:0] node12651;
	wire [4-1:0] node12654;
	wire [4-1:0] node12655;
	wire [4-1:0] node12657;
	wire [4-1:0] node12660;
	wire [4-1:0] node12663;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12667;
	wire [4-1:0] node12670;
	wire [4-1:0] node12671;
	wire [4-1:0] node12674;
	wire [4-1:0] node12675;
	wire [4-1:0] node12679;
	wire [4-1:0] node12681;
	wire [4-1:0] node12684;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12692;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12699;
	wire [4-1:0] node12702;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12710;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12714;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12722;
	wire [4-1:0] node12724;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12730;
	wire [4-1:0] node12731;
	wire [4-1:0] node12732;
	wire [4-1:0] node12733;
	wire [4-1:0] node12736;
	wire [4-1:0] node12737;
	wire [4-1:0] node12741;
	wire [4-1:0] node12744;
	wire [4-1:0] node12745;
	wire [4-1:0] node12747;
	wire [4-1:0] node12750;
	wire [4-1:0] node12752;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12758;
	wire [4-1:0] node12759;
	wire [4-1:0] node12763;
	wire [4-1:0] node12764;
	wire [4-1:0] node12765;
	wire [4-1:0] node12768;
	wire [4-1:0] node12771;
	wire [4-1:0] node12773;
	wire [4-1:0] node12776;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12779;
	wire [4-1:0] node12781;
	wire [4-1:0] node12784;
	wire [4-1:0] node12787;
	wire [4-1:0] node12789;
	wire [4-1:0] node12790;
	wire [4-1:0] node12792;
	wire [4-1:0] node12795;
	wire [4-1:0] node12797;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12805;
	wire [4-1:0] node12807;
	wire [4-1:0] node12810;
	wire [4-1:0] node12812;
	wire [4-1:0] node12813;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12819;
	wire [4-1:0] node12820;
	wire [4-1:0] node12821;
	wire [4-1:0] node12823;
	wire [4-1:0] node12826;
	wire [4-1:0] node12827;
	wire [4-1:0] node12828;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12836;
	wire [4-1:0] node12839;
	wire [4-1:0] node12842;
	wire [4-1:0] node12843;
	wire [4-1:0] node12848;
	wire [4-1:0] node12849;
	wire [4-1:0] node12850;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12857;
	wire [4-1:0] node12858;
	wire [4-1:0] node12859;
	wire [4-1:0] node12863;
	wire [4-1:0] node12866;
	wire [4-1:0] node12867;
	wire [4-1:0] node12869;
	wire [4-1:0] node12871;
	wire [4-1:0] node12875;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12881;
	wire [4-1:0] node12882;
	wire [4-1:0] node12883;
	wire [4-1:0] node12886;
	wire [4-1:0] node12890;
	wire [4-1:0] node12892;
	wire [4-1:0] node12893;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12900;
	wire [4-1:0] node12901;
	wire [4-1:0] node12906;
	wire [4-1:0] node12908;
	wire [4-1:0] node12909;
	wire [4-1:0] node12910;
	wire [4-1:0] node12911;
	wire [4-1:0] node12912;
	wire [4-1:0] node12914;
	wire [4-1:0] node12916;
	wire [4-1:0] node12918;
	wire [4-1:0] node12919;
	wire [4-1:0] node12924;
	wire [4-1:0] node12926;
	wire [4-1:0] node12927;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12931;
	wire [4-1:0] node12932;
	wire [4-1:0] node12936;
	wire [4-1:0] node12938;
	wire [4-1:0] node12939;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12951;
	wire [4-1:0] node12952;
	wire [4-1:0] node12955;
	wire [4-1:0] node12956;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12962;
	wire [4-1:0] node12967;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12970;
	wire [4-1:0] node12971;
	wire [4-1:0] node12972;
	wire [4-1:0] node12974;
	wire [4-1:0] node12976;
	wire [4-1:0] node12980;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12985;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12993;
	wire [4-1:0] node12994;
	wire [4-1:0] node12995;
	wire [4-1:0] node12999;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13004;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13014;
	wire [4-1:0] node13018;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13026;
	wire [4-1:0] node13031;
	wire [4-1:0] node13033;
	wire [4-1:0] node13035;
	wire [4-1:0] node13036;
	wire [4-1:0] node13040;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13043;
	wire [4-1:0] node13047;
	wire [4-1:0] node13048;
	wire [4-1:0] node13049;
	wire [4-1:0] node13053;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13060;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13067;
	wire [4-1:0] node13068;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13072;
	wire [4-1:0] node13077;
	wire [4-1:0] node13080;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13084;
	wire [4-1:0] node13087;
	wire [4-1:0] node13088;
	wire [4-1:0] node13092;
	wire [4-1:0] node13094;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13103;
	wire [4-1:0] node13107;
	wire [4-1:0] node13108;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13118;
	wire [4-1:0] node13121;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13124;
	wire [4-1:0] node13125;
	wire [4-1:0] node13129;
	wire [4-1:0] node13131;
	wire [4-1:0] node13136;
	wire [4-1:0] node13138;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13149;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13157;
	wire [4-1:0] node13160;
	wire [4-1:0] node13161;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13168;
	wire [4-1:0] node13171;
	wire [4-1:0] node13172;
	wire [4-1:0] node13174;
	wire [4-1:0] node13175;
	wire [4-1:0] node13176;
	wire [4-1:0] node13180;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;

	assign outp = (inp[8]) ? node6754 : node1;
		assign node1 = (inp[9]) ? node3497 : node2;
			assign node2 = (inp[6]) ? node782 : node3;
				assign node3 = (inp[15]) ? node465 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[2]) ? node277 : node6;
							assign node6 = (inp[1]) ? node160 : node7;
								assign node7 = (inp[14]) ? node77 : node8;
									assign node8 = (inp[13]) ? node48 : node9;
										assign node9 = (inp[10]) ? node37 : node10;
											assign node10 = (inp[12]) ? node26 : node11;
												assign node11 = (inp[5]) ? node19 : node12;
													assign node12 = (inp[4]) ? node16 : node13;
														assign node13 = (inp[3]) ? 4'b0000 : 4'b1111;
														assign node16 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node19 = (inp[11]) ? 4'b0100 : node20;
														assign node20 = (inp[4]) ? node22 : 4'b0000;
															assign node22 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node26 = (inp[3]) ? node32 : node27;
													assign node27 = (inp[5]) ? node29 : 4'b1111;
														assign node29 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node32 = (inp[11]) ? 4'b1000 : node33;
														assign node33 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node37 = (inp[3]) ? node43 : node38;
												assign node38 = (inp[7]) ? node40 : 4'b0000;
													assign node40 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node43 = (inp[4]) ? 4'b0100 : node44;
													assign node44 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node48 = (inp[12]) ? node62 : node49;
											assign node49 = (inp[3]) ? node57 : node50;
												assign node50 = (inp[7]) ? node52 : 4'b1000;
													assign node52 = (inp[5]) ? node54 : 4'b1111;
														assign node54 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node57 = (inp[7]) ? node59 : 4'b1100;
													assign node59 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node62 = (inp[10]) ? node72 : node63;
												assign node63 = (inp[3]) ? node67 : node64;
													assign node64 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node67 = (inp[7]) ? node69 : 4'b0100;
														assign node69 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node72 = (inp[3]) ? node74 : 4'b1000;
													assign node74 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node77 = (inp[11]) ? node117 : node78;
										assign node78 = (inp[13]) ? node102 : node79;
											assign node79 = (inp[12]) ? node93 : node80;
												assign node80 = (inp[10]) ? node90 : node81;
													assign node81 = (inp[3]) ? 4'b1001 : node82;
														assign node82 = (inp[4]) ? node84 : 4'b1111;
															assign node84 = (inp[7]) ? node86 : 4'b1001;
																assign node86 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node90 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node93 = (inp[3]) ? 4'b1001 : node94;
													assign node94 = (inp[4]) ? node98 : node95;
														assign node95 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node98 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node102 = (inp[3]) ? node112 : node103;
												assign node103 = (inp[10]) ? node109 : node104;
													assign node104 = (inp[7]) ? node106 : 4'b0001;
														assign node106 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node109 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node112 = (inp[12]) ? 4'b0101 : node113;
													assign node113 = (inp[10]) ? 4'b1101 : 4'b0001;
										assign node117 = (inp[3]) ? node139 : node118;
											assign node118 = (inp[4]) ? node130 : node119;
												assign node119 = (inp[7]) ? node127 : node120;
													assign node120 = (inp[10]) ? 4'b0000 : node121;
														assign node121 = (inp[13]) ? 4'b0000 : node122;
															assign node122 = (inp[5]) ? 4'b1100 : 4'b1111;
													assign node127 = (inp[12]) ? 4'b1100 : 4'b1111;
												assign node130 = (inp[13]) ? node136 : node131;
													assign node131 = (inp[7]) ? 4'b0000 : node132;
														assign node132 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node136 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node139 = (inp[7]) ? node149 : node140;
												assign node140 = (inp[12]) ? node142 : 4'b1100;
													assign node142 = (inp[10]) ? node146 : node143;
														assign node143 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node146 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node149 = (inp[4]) ? node155 : node150;
													assign node150 = (inp[10]) ? node152 : 4'b0000;
														assign node152 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node155 = (inp[13]) ? 4'b1100 : node156;
														assign node156 = (inp[12]) ? 4'b1000 : 4'b0100;
								assign node160 = (inp[13]) ? node230 : node161;
									assign node161 = (inp[11]) ? node205 : node162;
										assign node162 = (inp[14]) ? node184 : node163;
											assign node163 = (inp[10]) ? node175 : node164;
												assign node164 = (inp[12]) ? node168 : node165;
													assign node165 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node168 = (inp[5]) ? 4'b1101 : node169;
														assign node169 = (inp[3]) ? 4'b1001 : node170;
															assign node170 = (inp[4]) ? 4'b1001 : 4'b1111;
												assign node175 = (inp[3]) ? node179 : node176;
													assign node176 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node179 = (inp[7]) ? node181 : 4'b0101;
														assign node181 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node184 = (inp[12]) ? node190 : node185;
												assign node185 = (inp[3]) ? node187 : 4'b0000;
													assign node187 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node190 = (inp[10]) ? node200 : node191;
													assign node191 = (inp[5]) ? node195 : node192;
														assign node192 = (inp[4]) ? 4'b1000 : 4'b1111;
														assign node195 = (inp[4]) ? 4'b1100 : node196;
															assign node196 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node200 = (inp[4]) ? node202 : 4'b0000;
														assign node202 = (inp[3]) ? 4'b0100 : 4'b0000;
										assign node205 = (inp[3]) ? node215 : node206;
											assign node206 = (inp[10]) ? 4'b0001 : node207;
												assign node207 = (inp[4]) ? node211 : node208;
													assign node208 = (inp[5]) ? 4'b0101 : 4'b1111;
													assign node211 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node215 = (inp[12]) ? node221 : node216;
												assign node216 = (inp[7]) ? node218 : 4'b0101;
													assign node218 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node221 = (inp[10]) ? node227 : node222;
													assign node222 = (inp[7]) ? 4'b1001 : node223;
														assign node223 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node227 = (inp[5]) ? 4'b0001 : 4'b0101;
									assign node230 = (inp[3]) ? node244 : node231;
										assign node231 = (inp[10]) ? node235 : node232;
											assign node232 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node235 = (inp[7]) ? node239 : node236;
												assign node236 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node239 = (inp[4]) ? 4'b1001 : node240;
													assign node240 = (inp[14]) ? 4'b1111 : 4'b1101;
										assign node244 = (inp[14]) ? node260 : node245;
											assign node245 = (inp[7]) ? node251 : node246;
												assign node246 = (inp[4]) ? 4'b1101 : node247;
													assign node247 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node251 = (inp[4]) ? node257 : node252;
													assign node252 = (inp[11]) ? node254 : 4'b1001;
														assign node254 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node257 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node260 = (inp[11]) ? node272 : node261;
												assign node261 = (inp[10]) ? 4'b1100 : node262;
													assign node262 = (inp[12]) ? node266 : node263;
														assign node263 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node266 = (inp[7]) ? node268 : 4'b0100;
															assign node268 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node272 = (inp[4]) ? 4'b1101 : node273;
													assign node273 = (inp[7]) ? 4'b1001 : 4'b1101;
							assign node277 = (inp[5]) ? node279 : 4'b1111;
								assign node279 = (inp[3]) ? node347 : node280;
									assign node280 = (inp[4]) ? node312 : node281;
										assign node281 = (inp[7]) ? 4'b1111 : node282;
											assign node282 = (inp[12]) ? node298 : node283;
												assign node283 = (inp[13]) ? node289 : node284;
													assign node284 = (inp[10]) ? node286 : 4'b0000;
														assign node286 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node289 = (inp[1]) ? node293 : node290;
														assign node290 = (inp[10]) ? 4'b1000 : 4'b0001;
														assign node293 = (inp[11]) ? 4'b1001 : node294;
															assign node294 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node298 = (inp[13]) ? node304 : node299;
													assign node299 = (inp[10]) ? node301 : 4'b1111;
														assign node301 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node304 = (inp[10]) ? 4'b1001 : node305;
														assign node305 = (inp[11]) ? node307 : 4'b0001;
															assign node307 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node312 = (inp[1]) ? node326 : node313;
											assign node313 = (inp[14]) ? node319 : node314;
												assign node314 = (inp[12]) ? 4'b0000 : node315;
													assign node315 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node319 = (inp[11]) ? 4'b1000 : node320;
													assign node320 = (inp[13]) ? 4'b0001 : node321;
														assign node321 = (inp[12]) ? 4'b1111 : 4'b1001;
											assign node326 = (inp[13]) ? node336 : node327;
												assign node327 = (inp[10]) ? node331 : node328;
													assign node328 = (inp[12]) ? 4'b1111 : 4'b0001;
													assign node331 = (inp[11]) ? 4'b0001 : node332;
														assign node332 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node336 = (inp[12]) ? node342 : node337;
													assign node337 = (inp[14]) ? node339 : 4'b1001;
														assign node339 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node342 = (inp[10]) ? 4'b1001 : node343;
														assign node343 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node347 = (inp[7]) ? node399 : node348;
										assign node348 = (inp[1]) ? node376 : node349;
											assign node349 = (inp[14]) ? node363 : node350;
												assign node350 = (inp[10]) ? node360 : node351;
													assign node351 = (inp[13]) ? node357 : node352;
														assign node352 = (inp[12]) ? node354 : 4'b0100;
															assign node354 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node357 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node360 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node363 = (inp[11]) ? node371 : node364;
													assign node364 = (inp[12]) ? 4'b1101 : node365;
														assign node365 = (inp[13]) ? node367 : 4'b0101;
															assign node367 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node371 = (inp[13]) ? node373 : 4'b0100;
														assign node373 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node376 = (inp[14]) ? node384 : node377;
												assign node377 = (inp[12]) ? node381 : node378;
													assign node378 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node381 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node384 = (inp[11]) ? node394 : node385;
													assign node385 = (inp[10]) ? 4'b0100 : node386;
														assign node386 = (inp[12]) ? node390 : node387;
															assign node387 = (inp[4]) ? 4'b1100 : 4'b0100;
															assign node390 = (inp[4]) ? 4'b0100 : 4'b1000;
													assign node394 = (inp[10]) ? 4'b0101 : node395;
														assign node395 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node399 = (inp[4]) ? node439 : node400;
											assign node400 = (inp[1]) ? node420 : node401;
												assign node401 = (inp[14]) ? node413 : node402;
													assign node402 = (inp[11]) ? node408 : node403;
														assign node403 = (inp[12]) ? 4'b0000 : node404;
															assign node404 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node408 = (inp[13]) ? 4'b1000 : node409;
															assign node409 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node413 = (inp[11]) ? 4'b1000 : node414;
														assign node414 = (inp[13]) ? node416 : 4'b0001;
															assign node416 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node420 = (inp[11]) ? node430 : node421;
													assign node421 = (inp[14]) ? node423 : 4'b0001;
														assign node423 = (inp[12]) ? node425 : 4'b0000;
															assign node425 = (inp[13]) ? node427 : 4'b1000;
																assign node427 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node430 = (inp[13]) ? node434 : node431;
														assign node431 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node434 = (inp[12]) ? node436 : 4'b1001;
															assign node436 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node439 = (inp[1]) ? node451 : node440;
												assign node440 = (inp[14]) ? node442 : 4'b0100;
													assign node442 = (inp[11]) ? node444 : 4'b1001;
														assign node444 = (inp[12]) ? node446 : 4'b1100;
															assign node446 = (inp[13]) ? 4'b0100 : node447;
																assign node447 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node451 = (inp[12]) ? node459 : node452;
													assign node452 = (inp[11]) ? node456 : node453;
														assign node453 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node456 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node459 = (inp[13]) ? node461 : 4'b1001;
														assign node461 = (inp[10]) ? 4'b1101 : 4'b0101;
					assign node465 = (inp[0]) ? 4'b1001 : node466;
						assign node466 = (inp[5]) ? node534 : node467;
							assign node467 = (inp[2]) ? 4'b1011 : node468;
								assign node468 = (inp[3]) ? node470 : 4'b1011;
									assign node470 = (inp[7]) ? node510 : node471;
										assign node471 = (inp[13]) ? node491 : node472;
											assign node472 = (inp[10]) ? node484 : node473;
												assign node473 = (inp[12]) ? node477 : node474;
													assign node474 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node477 = (inp[4]) ? node479 : 4'b1011;
														assign node479 = (inp[11]) ? node481 : 4'b1000;
															assign node481 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node484 = (inp[1]) ? node488 : node485;
													assign node485 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node488 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node491 = (inp[10]) ? node501 : node492;
												assign node492 = (inp[12]) ? node494 : 4'b1000;
													assign node494 = (inp[1]) ? 4'b0001 : node495;
														assign node495 = (inp[4]) ? 4'b0000 : node496;
															assign node496 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node501 = (inp[1]) ? node507 : node502;
													assign node502 = (inp[14]) ? node504 : 4'b1000;
														assign node504 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node507 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node510 = (inp[4]) ? node512 : 4'b1011;
											assign node512 = (inp[1]) ? node524 : node513;
												assign node513 = (inp[13]) ? node521 : node514;
													assign node514 = (inp[12]) ? node518 : node515;
														assign node515 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node518 = (inp[11]) ? 4'b0000 : 4'b1011;
													assign node521 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node524 = (inp[13]) ? node528 : node525;
													assign node525 = (inp[12]) ? 4'b1011 : 4'b0001;
													assign node528 = (inp[14]) ? node530 : 4'b1001;
														assign node530 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node534 = (inp[2]) ? node714 : node535;
								assign node535 = (inp[1]) ? node625 : node536;
									assign node536 = (inp[11]) ? node590 : node537;
										assign node537 = (inp[14]) ? node555 : node538;
											assign node538 = (inp[3]) ? node544 : node539;
												assign node539 = (inp[10]) ? 4'b1100 : node540;
													assign node540 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node544 = (inp[4]) ? node552 : node545;
													assign node545 = (inp[12]) ? node549 : node546;
														assign node546 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node549 = (inp[7]) ? 4'b0100 : 4'b1100;
													assign node552 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node555 = (inp[13]) ? node571 : node556;
												assign node556 = (inp[3]) ? node562 : node557;
													assign node557 = (inp[12]) ? 4'b1001 : node558;
														assign node558 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node562 = (inp[4]) ? node568 : node563;
														assign node563 = (inp[10]) ? node565 : 4'b1101;
															assign node565 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node568 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node571 = (inp[10]) ? node581 : node572;
													assign node572 = (inp[4]) ? 4'b0001 : node573;
														assign node573 = (inp[12]) ? 4'b0101 : node574;
															assign node574 = (inp[7]) ? 4'b0001 : node575;
																assign node575 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node581 = (inp[12]) ? 4'b0001 : node582;
														assign node582 = (inp[4]) ? 4'b1001 : node583;
															assign node583 = (inp[7]) ? 4'b1101 : node584;
																assign node584 = (inp[3]) ? 4'b1001 : 4'b1101;
										assign node590 = (inp[13]) ? node604 : node591;
											assign node591 = (inp[12]) ? node599 : node592;
												assign node592 = (inp[3]) ? 4'b0000 : node593;
													assign node593 = (inp[14]) ? 4'b0100 : node594;
														assign node594 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node599 = (inp[10]) ? node601 : 4'b1000;
													assign node601 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node604 = (inp[12]) ? node614 : node605;
												assign node605 = (inp[3]) ? node609 : node606;
													assign node606 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node609 = (inp[4]) ? 4'b1000 : node610;
														assign node610 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node614 = (inp[10]) ? node620 : node615;
													assign node615 = (inp[7]) ? 4'b0100 : node616;
														assign node616 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node620 = (inp[7]) ? node622 : 4'b1000;
														assign node622 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node625 = (inp[11]) ? node675 : node626;
										assign node626 = (inp[14]) ? node650 : node627;
											assign node627 = (inp[13]) ? node639 : node628;
												assign node628 = (inp[7]) ? node634 : node629;
													assign node629 = (inp[12]) ? node631 : 4'b0001;
														assign node631 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node634 = (inp[12]) ? node636 : 4'b0101;
														assign node636 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node639 = (inp[3]) ? node647 : node640;
													assign node640 = (inp[4]) ? 4'b1101 : node641;
														assign node641 = (inp[7]) ? node643 : 4'b0101;
															assign node643 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node647 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node650 = (inp[10]) ? node666 : node651;
												assign node651 = (inp[13]) ? node661 : node652;
													assign node652 = (inp[12]) ? node654 : 4'b0100;
														assign node654 = (inp[3]) ? node658 : node655;
															assign node655 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node658 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node661 = (inp[4]) ? node663 : 4'b1100;
														assign node663 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node666 = (inp[13]) ? node668 : 4'b0000;
													assign node668 = (inp[3]) ? 4'b1000 : node669;
														assign node669 = (inp[7]) ? node671 : 4'b1100;
															assign node671 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node675 = (inp[13]) ? node699 : node676;
											assign node676 = (inp[12]) ? node688 : node677;
												assign node677 = (inp[3]) ? node683 : node678;
													assign node678 = (inp[7]) ? node680 : 4'b0101;
														assign node680 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node683 = (inp[7]) ? node685 : 4'b0001;
														assign node685 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node688 = (inp[10]) ? node692 : node689;
													assign node689 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node692 = (inp[4]) ? 4'b0101 : node693;
														assign node693 = (inp[7]) ? node695 : 4'b0101;
															assign node695 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node699 = (inp[3]) ? node709 : node700;
												assign node700 = (inp[7]) ? node702 : 4'b1101;
													assign node702 = (inp[4]) ? node706 : node703;
														assign node703 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node706 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node709 = (inp[4]) ? 4'b1001 : node710;
													assign node710 = (inp[7]) ? 4'b1101 : 4'b1001;
								assign node714 = (inp[3]) ? node716 : 4'b1011;
									assign node716 = (inp[7]) ? node752 : node717;
										assign node717 = (inp[1]) ? node735 : node718;
											assign node718 = (inp[13]) ? node724 : node719;
												assign node719 = (inp[14]) ? node721 : 4'b0000;
													assign node721 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node724 = (inp[14]) ? node730 : node725;
													assign node725 = (inp[12]) ? node727 : 4'b1000;
														assign node727 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node730 = (inp[11]) ? node732 : 4'b0001;
														assign node732 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node735 = (inp[13]) ? node745 : node736;
												assign node736 = (inp[14]) ? node742 : node737;
													assign node737 = (inp[12]) ? node739 : 4'b0001;
														assign node739 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node742 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node745 = (inp[11]) ? node749 : node746;
													assign node746 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node749 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node752 = (inp[4]) ? node754 : 4'b1011;
											assign node754 = (inp[13]) ? node768 : node755;
												assign node755 = (inp[12]) ? node761 : node756;
													assign node756 = (inp[1]) ? node758 : 4'b0000;
														assign node758 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node761 = (inp[10]) ? node763 : 4'b1011;
														assign node763 = (inp[14]) ? 4'b0000 : node764;
															assign node764 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node768 = (inp[14]) ? node772 : node769;
													assign node769 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node772 = (inp[11]) ? node778 : node773;
														assign node773 = (inp[1]) ? node775 : 4'b0001;
															assign node775 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node778 = (inp[1]) ? 4'b1001 : 4'b1000;
				assign node782 = (inp[5]) ? node1956 : node783;
					assign node783 = (inp[0]) ? node1667 : node784;
						assign node784 = (inp[11]) ? node1256 : node785;
							assign node785 = (inp[10]) ? node1019 : node786;
								assign node786 = (inp[1]) ? node896 : node787;
									assign node787 = (inp[14]) ? node845 : node788;
										assign node788 = (inp[12]) ? node816 : node789;
											assign node789 = (inp[15]) ? node803 : node790;
												assign node790 = (inp[4]) ? node792 : 4'b0000;
													assign node792 = (inp[13]) ? node798 : node793;
														assign node793 = (inp[3]) ? 4'b0001 : node794;
															assign node794 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node798 = (inp[3]) ? 4'b0100 : node799;
															assign node799 = (inp[2]) ? 4'b1000 : 4'b0100;
												assign node803 = (inp[13]) ? node805 : 4'b0100;
													assign node805 = (inp[4]) ? node811 : node806;
														assign node806 = (inp[7]) ? node808 : 4'b1100;
															assign node808 = (inp[2]) ? 4'b1100 : 4'b0100;
														assign node811 = (inp[3]) ? 4'b0000 : node812;
															assign node812 = (inp[7]) ? 4'b0000 : 4'b1100;
											assign node816 = (inp[13]) ? node828 : node817;
												assign node817 = (inp[15]) ? node819 : 4'b1000;
													assign node819 = (inp[3]) ? node825 : node820;
														assign node820 = (inp[4]) ? node822 : 4'b1000;
															assign node822 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node825 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node828 = (inp[2]) ? node838 : node829;
													assign node829 = (inp[4]) ? node833 : node830;
														assign node830 = (inp[3]) ? 4'b1100 : 4'b0100;
														assign node833 = (inp[15]) ? 4'b1100 : node834;
															assign node834 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node838 = (inp[3]) ? node842 : node839;
														assign node839 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node842 = (inp[15]) ? 4'b0000 : 4'b1000;
										assign node845 = (inp[13]) ? node871 : node846;
											assign node846 = (inp[3]) ? node852 : node847;
												assign node847 = (inp[15]) ? 4'b1001 : node848;
													assign node848 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node852 = (inp[2]) ? node860 : node853;
													assign node853 = (inp[12]) ? 4'b1100 : node854;
														assign node854 = (inp[7]) ? 4'b0100 : node855;
															assign node855 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node860 = (inp[12]) ? node868 : node861;
														assign node861 = (inp[7]) ? 4'b1101 : node862;
															assign node862 = (inp[4]) ? node864 : 4'b1101;
																assign node864 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node868 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node871 = (inp[3]) ? node883 : node872;
												assign node872 = (inp[2]) ? 4'b0101 : node873;
													assign node873 = (inp[12]) ? node879 : node874;
														assign node874 = (inp[15]) ? node876 : 4'b0000;
															assign node876 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node879 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node883 = (inp[2]) ? node893 : node884;
													assign node884 = (inp[15]) ? node890 : node885;
														assign node885 = (inp[12]) ? node887 : 4'b1100;
															assign node887 = (inp[4]) ? 4'b0100 : 4'b1100;
														assign node890 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node893 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node896 = (inp[14]) ? node958 : node897;
										assign node897 = (inp[2]) ? node927 : node898;
											assign node898 = (inp[3]) ? node912 : node899;
												assign node899 = (inp[4]) ? node903 : node900;
													assign node900 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node903 = (inp[12]) ? 4'b0000 : node904;
														assign node904 = (inp[7]) ? node906 : 4'b0100;
															assign node906 = (inp[15]) ? node908 : 4'b0000;
																assign node908 = (inp[13]) ? 4'b0000 : 4'b0101;
												assign node912 = (inp[15]) ? node920 : node913;
													assign node913 = (inp[7]) ? 4'b0100 : node914;
														assign node914 = (inp[13]) ? 4'b1100 : node915;
															assign node915 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node920 = (inp[7]) ? node922 : 4'b0100;
														assign node922 = (inp[12]) ? 4'b0000 : node923;
															assign node923 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node927 = (inp[3]) ? node941 : node928;
												assign node928 = (inp[13]) ? node936 : node929;
													assign node929 = (inp[12]) ? 4'b1001 : node930;
														assign node930 = (inp[15]) ? node932 : 4'b0001;
															assign node932 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node936 = (inp[12]) ? 4'b0001 : node937;
														assign node937 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node941 = (inp[15]) ? node947 : node942;
													assign node942 = (inp[7]) ? node944 : 4'b0100;
														assign node944 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node947 = (inp[4]) ? 4'b0001 : node948;
														assign node948 = (inp[7]) ? node952 : node949;
															assign node949 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node952 = (inp[13]) ? node954 : 4'b0101;
																assign node954 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node958 = (inp[2]) ? node992 : node959;
											assign node959 = (inp[13]) ? node985 : node960;
												assign node960 = (inp[3]) ? node968 : node961;
													assign node961 = (inp[12]) ? 4'b0000 : node962;
														assign node962 = (inp[4]) ? node964 : 4'b0000;
															assign node964 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node968 = (inp[15]) ? node972 : node969;
														assign node969 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node972 = (inp[12]) ? node980 : node973;
															assign node973 = (inp[4]) ? node977 : node974;
																assign node974 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node977 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node980 = (inp[7]) ? node982 : 4'b0000;
																assign node982 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node985 = (inp[12]) ? node987 : 4'b1001;
													assign node987 = (inp[15]) ? node989 : 4'b0000;
														assign node989 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node992 = (inp[4]) ? node1016 : node993;
												assign node993 = (inp[15]) ? node1005 : node994;
													assign node994 = (inp[3]) ? node1000 : node995;
														assign node995 = (inp[12]) ? 4'b1100 : node996;
															assign node996 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node1000 = (inp[13]) ? 4'b0000 : node1001;
															assign node1001 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1005 = (inp[13]) ? node1007 : 4'b0100;
														assign node1007 = (inp[12]) ? 4'b0100 : node1008;
															assign node1008 = (inp[3]) ? node1012 : node1009;
																assign node1009 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node1012 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node1016 = (inp[7]) ? 4'b1100 : 4'b0100;
								assign node1019 = (inp[12]) ? node1133 : node1020;
									assign node1020 = (inp[13]) ? node1082 : node1021;
										assign node1021 = (inp[3]) ? node1053 : node1022;
											assign node1022 = (inp[2]) ? node1038 : node1023;
												assign node1023 = (inp[7]) ? node1033 : node1024;
													assign node1024 = (inp[1]) ? 4'b1000 : node1025;
														assign node1025 = (inp[14]) ? 4'b1000 : node1026;
															assign node1026 = (inp[4]) ? node1028 : 4'b0100;
																assign node1028 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node1033 = (inp[1]) ? node1035 : 4'b0101;
														assign node1035 = (inp[15]) ? 4'b0100 : 4'b1000;
												assign node1038 = (inp[14]) ? node1046 : node1039;
													assign node1039 = (inp[1]) ? 4'b0001 : node1040;
														assign node1040 = (inp[4]) ? node1042 : 4'b0000;
															assign node1042 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1046 = (inp[1]) ? 4'b0000 : node1047;
														assign node1047 = (inp[15]) ? 4'b0101 : node1048;
															assign node1048 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node1053 = (inp[15]) ? node1067 : node1054;
												assign node1054 = (inp[4]) ? node1058 : node1055;
													assign node1055 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node1058 = (inp[7]) ? node1064 : node1059;
														assign node1059 = (inp[2]) ? 4'b1100 : node1060;
															assign node1060 = (inp[1]) ? 4'b0100 : 4'b1001;
														assign node1064 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node1067 = (inp[14]) ? node1069 : 4'b1000;
													assign node1069 = (inp[4]) ? node1077 : node1070;
														assign node1070 = (inp[2]) ? node1074 : node1071;
															assign node1071 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node1074 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node1077 = (inp[1]) ? 4'b0001 : node1078;
															assign node1078 = (inp[7]) ? 4'b0001 : 4'b1000;
										assign node1082 = (inp[3]) ? node1104 : node1083;
											assign node1083 = (inp[15]) ? node1093 : node1084;
												assign node1084 = (inp[4]) ? node1088 : node1085;
													assign node1085 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node1088 = (inp[2]) ? node1090 : 4'b1100;
														assign node1090 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node1093 = (inp[7]) ? node1099 : node1094;
													assign node1094 = (inp[2]) ? 4'b1100 : node1095;
														assign node1095 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node1099 = (inp[1]) ? node1101 : 4'b1000;
														assign node1101 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node1104 = (inp[2]) ? node1120 : node1105;
												assign node1105 = (inp[15]) ? 4'b1100 : node1106;
													assign node1106 = (inp[1]) ? node1114 : node1107;
														assign node1107 = (inp[7]) ? node1111 : node1108;
															assign node1108 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node1111 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1114 = (inp[4]) ? 4'b1101 : node1115;
															assign node1115 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node1120 = (inp[15]) ? node1124 : node1121;
													assign node1121 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node1124 = (inp[4]) ? 4'b1000 : node1125;
														assign node1125 = (inp[7]) ? node1127 : 4'b1001;
															assign node1127 = (inp[1]) ? 4'b1101 : node1128;
																assign node1128 = (inp[14]) ? 4'b1101 : 4'b1100;
									assign node1133 = (inp[1]) ? node1211 : node1134;
										assign node1134 = (inp[2]) ? node1168 : node1135;
											assign node1135 = (inp[14]) ? node1155 : node1136;
												assign node1136 = (inp[4]) ? node1144 : node1137;
													assign node1137 = (inp[15]) ? 4'b0100 : node1138;
														assign node1138 = (inp[7]) ? node1140 : 4'b0000;
															assign node1140 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node1144 = (inp[3]) ? node1148 : node1145;
														assign node1145 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1148 = (inp[15]) ? node1152 : node1149;
															assign node1149 = (inp[13]) ? 4'b0101 : 4'b1001;
															assign node1152 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node1155 = (inp[15]) ? 4'b0000 : node1156;
													assign node1156 = (inp[4]) ? node1162 : node1157;
														assign node1157 = (inp[13]) ? 4'b0000 : node1158;
															assign node1158 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node1162 = (inp[13]) ? 4'b0100 : node1163;
															assign node1163 = (inp[3]) ? 4'b1000 : 4'b0000;
											assign node1168 = (inp[14]) ? node1192 : node1169;
												assign node1169 = (inp[13]) ? node1181 : node1170;
													assign node1170 = (inp[15]) ? node1176 : node1171;
														assign node1171 = (inp[7]) ? 4'b0000 : node1172;
															assign node1172 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1176 = (inp[3]) ? node1178 : 4'b0100;
															assign node1178 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1181 = (inp[3]) ? 4'b0000 : node1182;
														assign node1182 = (inp[7]) ? node1186 : node1183;
															assign node1183 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node1186 = (inp[4]) ? 4'b1100 : node1187;
																assign node1187 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node1192 = (inp[13]) ? node1200 : node1193;
													assign node1193 = (inp[7]) ? node1197 : node1194;
														assign node1194 = (inp[3]) ? 4'b0000 : 4'b1001;
														assign node1197 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node1200 = (inp[3]) ? node1204 : node1201;
														assign node1201 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node1204 = (inp[4]) ? node1208 : node1205;
															assign node1205 = (inp[15]) ? 4'b0101 : 4'b0000;
															assign node1208 = (inp[15]) ? 4'b0000 : 4'b0100;
										assign node1211 = (inp[13]) ? node1237 : node1212;
											assign node1212 = (inp[7]) ? node1226 : node1213;
												assign node1213 = (inp[15]) ? node1215 : 4'b1100;
													assign node1215 = (inp[2]) ? node1223 : node1216;
														assign node1216 = (inp[4]) ? 4'b1000 : node1217;
															assign node1217 = (inp[3]) ? 4'b1100 : node1218;
																assign node1218 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1223 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node1226 = (inp[2]) ? node1230 : node1227;
													assign node1227 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1230 = (inp[4]) ? node1234 : node1231;
														assign node1231 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node1234 = (inp[15]) ? 4'b0000 : 4'b1000;
											assign node1237 = (inp[4]) ? node1245 : node1238;
												assign node1238 = (inp[7]) ? 4'b1000 : node1239;
													assign node1239 = (inp[2]) ? 4'b1000 : node1240;
														assign node1240 = (inp[3]) ? 4'b0001 : 4'b1000;
												assign node1245 = (inp[15]) ? node1253 : node1246;
													assign node1246 = (inp[14]) ? node1248 : 4'b1100;
														assign node1248 = (inp[3]) ? 4'b1100 : node1249;
															assign node1249 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node1253 = (inp[3]) ? 4'b0001 : 4'b1000;
							assign node1256 = (inp[1]) ? node1490 : node1257;
								assign node1257 = (inp[3]) ? node1361 : node1258;
									assign node1258 = (inp[13]) ? node1318 : node1259;
										assign node1259 = (inp[2]) ? node1301 : node1260;
											assign node1260 = (inp[7]) ? node1282 : node1261;
												assign node1261 = (inp[14]) ? node1271 : node1262;
													assign node1262 = (inp[15]) ? node1268 : node1263;
														assign node1263 = (inp[10]) ? node1265 : 4'b0001;
															assign node1265 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1268 = (inp[4]) ? 4'b0001 : 4'b0100;
													assign node1271 = (inp[10]) ? node1275 : node1272;
														assign node1272 = (inp[12]) ? 4'b1100 : 4'b0101;
														assign node1275 = (inp[15]) ? node1279 : node1276;
															assign node1276 = (inp[12]) ? 4'b0101 : 4'b1001;
															assign node1279 = (inp[4]) ? 4'b0001 : 4'b0100;
												assign node1282 = (inp[12]) ? node1294 : node1283;
													assign node1283 = (inp[10]) ? node1289 : node1284;
														assign node1284 = (inp[4]) ? node1286 : 4'b0100;
															assign node1286 = (inp[14]) ? 4'b0001 : 4'b0100;
														assign node1289 = (inp[14]) ? 4'b0100 : node1290;
															assign node1290 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node1294 = (inp[10]) ? 4'b0100 : node1295;
														assign node1295 = (inp[4]) ? 4'b1001 : node1296;
															assign node1296 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node1301 = (inp[15]) ? node1309 : node1302;
												assign node1302 = (inp[7]) ? node1306 : node1303;
													assign node1303 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1306 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node1309 = (inp[4]) ? 4'b0100 : node1310;
													assign node1310 = (inp[10]) ? 4'b0100 : node1311;
														assign node1311 = (inp[14]) ? 4'b1000 : node1312;
															assign node1312 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node1318 = (inp[2]) ? node1342 : node1319;
											assign node1319 = (inp[15]) ? node1327 : node1320;
												assign node1320 = (inp[4]) ? node1322 : 4'b1001;
													assign node1322 = (inp[12]) ? 4'b1001 : node1323;
														assign node1323 = (inp[7]) ? 4'b0101 : 4'b1101;
												assign node1327 = (inp[4]) ? node1335 : node1328;
													assign node1328 = (inp[7]) ? node1330 : 4'b0100;
														assign node1330 = (inp[12]) ? node1332 : 4'b1000;
															assign node1332 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1335 = (inp[7]) ? node1339 : node1336;
														assign node1336 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node1339 = (inp[12]) ? 4'b0100 : 4'b0001;
											assign node1342 = (inp[15]) ? node1354 : node1343;
												assign node1343 = (inp[12]) ? node1349 : node1344;
													assign node1344 = (inp[4]) ? 4'b1000 : node1345;
														assign node1345 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node1349 = (inp[10]) ? 4'b1000 : node1350;
														assign node1350 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node1354 = (inp[10]) ? node1358 : node1355;
													assign node1355 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1358 = (inp[7]) ? 4'b1000 : 4'b1100;
									assign node1361 = (inp[13]) ? node1429 : node1362;
										assign node1362 = (inp[2]) ? node1400 : node1363;
											assign node1363 = (inp[4]) ? node1383 : node1364;
												assign node1364 = (inp[7]) ? node1374 : node1365;
													assign node1365 = (inp[15]) ? node1367 : 4'b0001;
														assign node1367 = (inp[12]) ? node1371 : node1368;
															assign node1368 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node1371 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node1374 = (inp[15]) ? node1380 : node1375;
														assign node1375 = (inp[14]) ? node1377 : 4'b1101;
															assign node1377 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node1380 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node1383 = (inp[15]) ? node1391 : node1384;
													assign node1384 = (inp[12]) ? node1388 : node1385;
														assign node1385 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1388 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1391 = (inp[7]) ? 4'b1101 : node1392;
														assign node1392 = (inp[12]) ? node1396 : node1393;
															assign node1393 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node1396 = (inp[10]) ? 4'b0001 : 4'b1101;
											assign node1400 = (inp[4]) ? node1414 : node1401;
												assign node1401 = (inp[15]) ? node1407 : node1402;
													assign node1402 = (inp[14]) ? 4'b0000 : node1403;
														assign node1403 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node1407 = (inp[7]) ? node1409 : 4'b0000;
														assign node1409 = (inp[12]) ? node1411 : 4'b0100;
															assign node1411 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node1414 = (inp[15]) ? node1420 : node1415;
													assign node1415 = (inp[12]) ? 4'b1001 : node1416;
														assign node1416 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node1420 = (inp[7]) ? node1426 : node1421;
														assign node1421 = (inp[10]) ? node1423 : 4'b1000;
															assign node1423 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1426 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node1429 = (inp[14]) ? node1449 : node1430;
											assign node1430 = (inp[12]) ? node1440 : node1431;
												assign node1431 = (inp[10]) ? node1433 : 4'b0001;
													assign node1433 = (inp[2]) ? node1435 : 4'b1000;
														assign node1435 = (inp[4]) ? node1437 : 4'b1001;
															assign node1437 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node1440 = (inp[2]) ? node1442 : 4'b0000;
													assign node1442 = (inp[7]) ? 4'b0000 : node1443;
														assign node1443 = (inp[4]) ? node1445 : 4'b1000;
															assign node1445 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node1449 = (inp[2]) ? node1471 : node1450;
												assign node1450 = (inp[4]) ? node1464 : node1451;
													assign node1451 = (inp[15]) ? node1461 : node1452;
														assign node1452 = (inp[10]) ? node1458 : node1453;
															assign node1453 = (inp[7]) ? 4'b1101 : node1454;
																assign node1454 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node1458 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node1461 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node1464 = (inp[15]) ? node1468 : node1465;
														assign node1465 = (inp[7]) ? 4'b1000 : 4'b0100;
														assign node1468 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node1471 = (inp[4]) ? node1475 : node1472;
													assign node1472 = (inp[10]) ? 4'b1001 : 4'b1100;
													assign node1475 = (inp[15]) ? node1487 : node1476;
														assign node1476 = (inp[7]) ? node1482 : node1477;
															assign node1477 = (inp[10]) ? node1479 : 4'b1101;
																assign node1479 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node1482 = (inp[12]) ? 4'b1001 : node1483;
																assign node1483 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node1487 = (inp[7]) ? 4'b0001 : 4'b1001;
								assign node1490 = (inp[10]) ? node1592 : node1491;
									assign node1491 = (inp[2]) ? node1539 : node1492;
										assign node1492 = (inp[7]) ? node1514 : node1493;
											assign node1493 = (inp[13]) ? node1503 : node1494;
												assign node1494 = (inp[12]) ? 4'b0001 : node1495;
													assign node1495 = (inp[3]) ? node1499 : node1496;
														assign node1496 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node1499 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node1503 = (inp[14]) ? node1509 : node1504;
													assign node1504 = (inp[12]) ? node1506 : 4'b0101;
														assign node1506 = (inp[15]) ? 4'b0101 : 4'b0001;
													assign node1509 = (inp[4]) ? node1511 : 4'b0001;
														assign node1511 = (inp[15]) ? 4'b0001 : 4'b1101;
											assign node1514 = (inp[4]) ? node1522 : node1515;
												assign node1515 = (inp[3]) ? node1519 : node1516;
													assign node1516 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node1519 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node1522 = (inp[3]) ? node1528 : node1523;
													assign node1523 = (inp[12]) ? node1525 : 4'b0001;
														assign node1525 = (inp[15]) ? 4'b1001 : 4'b0001;
													assign node1528 = (inp[15]) ? node1536 : node1529;
														assign node1529 = (inp[13]) ? node1533 : node1530;
															assign node1530 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node1533 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node1536 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node1539 = (inp[15]) ? node1563 : node1540;
											assign node1540 = (inp[12]) ? node1552 : node1541;
												assign node1541 = (inp[3]) ? node1547 : node1542;
													assign node1542 = (inp[13]) ? 4'b1001 : node1543;
														assign node1543 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1547 = (inp[4]) ? node1549 : 4'b0001;
														assign node1549 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node1552 = (inp[13]) ? node1556 : node1553;
													assign node1553 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node1556 = (inp[3]) ? node1560 : node1557;
														assign node1557 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node1560 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node1563 = (inp[12]) ? node1579 : node1564;
												assign node1564 = (inp[13]) ? node1568 : node1565;
													assign node1565 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node1568 = (inp[4]) ? node1576 : node1569;
														assign node1569 = (inp[3]) ? node1573 : node1570;
															assign node1570 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node1573 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1576 = (inp[3]) ? 4'b0001 : 4'b1101;
												assign node1579 = (inp[13]) ? node1583 : node1580;
													assign node1580 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node1583 = (inp[4]) ? 4'b0001 : node1584;
														assign node1584 = (inp[7]) ? node1588 : node1585;
															assign node1585 = (inp[3]) ? 4'b0001 : 4'b0101;
															assign node1588 = (inp[3]) ? 4'b0101 : 4'b0001;
									assign node1592 = (inp[13]) ? node1638 : node1593;
										assign node1593 = (inp[2]) ? node1621 : node1594;
											assign node1594 = (inp[15]) ? node1608 : node1595;
												assign node1595 = (inp[7]) ? node1601 : node1596;
													assign node1596 = (inp[4]) ? node1598 : 4'b1001;
														assign node1598 = (inp[3]) ? 4'b0101 : 4'b1101;
													assign node1601 = (inp[4]) ? node1605 : node1602;
														assign node1602 = (inp[3]) ? 4'b1101 : 4'b0101;
														assign node1605 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node1608 = (inp[3]) ? node1614 : node1609;
													assign node1609 = (inp[14]) ? node1611 : 4'b0101;
														assign node1611 = (inp[12]) ? 4'b0101 : 4'b1001;
													assign node1614 = (inp[4]) ? node1618 : node1615;
														assign node1615 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node1618 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node1621 = (inp[15]) ? node1625 : node1622;
												assign node1622 = (inp[3]) ? 4'b1001 : 4'b0001;
												assign node1625 = (inp[3]) ? node1631 : node1626;
													assign node1626 = (inp[4]) ? 4'b0101 : node1627;
														assign node1627 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1631 = (inp[7]) ? node1635 : node1632;
														assign node1632 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1635 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node1638 = (inp[7]) ? node1652 : node1639;
											assign node1639 = (inp[15]) ? node1645 : node1640;
												assign node1640 = (inp[3]) ? node1642 : 4'b1001;
													assign node1642 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node1645 = (inp[4]) ? node1647 : 4'b1101;
													assign node1647 = (inp[3]) ? 4'b1001 : node1648;
														assign node1648 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node1652 = (inp[15]) ? node1660 : node1653;
												assign node1653 = (inp[4]) ? node1655 : 4'b1001;
													assign node1655 = (inp[2]) ? node1657 : 4'b1101;
														assign node1657 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node1660 = (inp[4]) ? node1664 : node1661;
													assign node1661 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node1664 = (inp[3]) ? 4'b1001 : 4'b1101;
						assign node1667 = (inp[15]) ? node1869 : node1668;
							assign node1668 = (inp[2]) ? 4'b1101 : node1669;
								assign node1669 = (inp[1]) ? node1765 : node1670;
									assign node1670 = (inp[14]) ? node1712 : node1671;
										assign node1671 = (inp[13]) ? node1687 : node1672;
											assign node1672 = (inp[3]) ? node1678 : node1673;
												assign node1673 = (inp[7]) ? node1675 : 4'b0000;
													assign node1675 = (inp[4]) ? 4'b0000 : 4'b1101;
												assign node1678 = (inp[10]) ? 4'b0100 : node1679;
													assign node1679 = (inp[12]) ? node1683 : node1680;
														assign node1680 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1683 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node1687 = (inp[3]) ? node1695 : node1688;
												assign node1688 = (inp[7]) ? node1690 : 4'b1000;
													assign node1690 = (inp[4]) ? node1692 : 4'b1101;
														assign node1692 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node1695 = (inp[4]) ? node1707 : node1696;
													assign node1696 = (inp[7]) ? node1702 : node1697;
														assign node1697 = (inp[10]) ? 4'b1100 : node1698;
															assign node1698 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node1702 = (inp[10]) ? 4'b1000 : node1703;
															assign node1703 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node1707 = (inp[12]) ? node1709 : 4'b1100;
														assign node1709 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node1712 = (inp[11]) ? node1740 : node1713;
											assign node1713 = (inp[13]) ? node1735 : node1714;
												assign node1714 = (inp[10]) ? node1726 : node1715;
													assign node1715 = (inp[3]) ? node1721 : node1716;
														assign node1716 = (inp[7]) ? 4'b1101 : node1717;
															assign node1717 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node1721 = (inp[4]) ? node1723 : 4'b1001;
															assign node1723 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node1726 = (inp[12]) ? node1732 : node1727;
														assign node1727 = (inp[3]) ? node1729 : 4'b0001;
															assign node1729 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node1732 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node1735 = (inp[3]) ? node1737 : 4'b0001;
													assign node1737 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node1740 = (inp[4]) ? node1750 : node1741;
												assign node1741 = (inp[3]) ? node1747 : node1742;
													assign node1742 = (inp[7]) ? 4'b1101 : node1743;
														assign node1743 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1747 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node1750 = (inp[3]) ? node1754 : node1751;
													assign node1751 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node1754 = (inp[7]) ? node1760 : node1755;
														assign node1755 = (inp[12]) ? node1757 : 4'b1100;
															assign node1757 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node1760 = (inp[10]) ? node1762 : 4'b0100;
															assign node1762 = (inp[13]) ? 4'b1100 : 4'b0100;
									assign node1765 = (inp[14]) ? node1815 : node1766;
										assign node1766 = (inp[13]) ? node1790 : node1767;
											assign node1767 = (inp[12]) ? node1779 : node1768;
												assign node1768 = (inp[3]) ? node1774 : node1769;
													assign node1769 = (inp[4]) ? 4'b0001 : node1770;
														assign node1770 = (inp[11]) ? 4'b0001 : 4'b1101;
													assign node1774 = (inp[7]) ? node1776 : 4'b0101;
														assign node1776 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1779 = (inp[10]) ? node1787 : node1780;
													assign node1780 = (inp[3]) ? node1782 : 4'b1101;
														assign node1782 = (inp[4]) ? node1784 : 4'b1001;
															assign node1784 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node1787 = (inp[3]) ? 4'b0101 : 4'b1101;
											assign node1790 = (inp[12]) ? node1802 : node1791;
												assign node1791 = (inp[4]) ? node1799 : node1792;
													assign node1792 = (inp[11]) ? node1794 : 4'b1101;
														assign node1794 = (inp[3]) ? 4'b1001 : node1795;
															assign node1795 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node1799 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node1802 = (inp[10]) ? node1806 : node1803;
													assign node1803 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node1806 = (inp[7]) ? node1808 : 4'b1101;
														assign node1808 = (inp[3]) ? node1812 : node1809;
															assign node1809 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node1812 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node1815 = (inp[11]) ? node1843 : node1816;
											assign node1816 = (inp[13]) ? node1830 : node1817;
												assign node1817 = (inp[10]) ? node1823 : node1818;
													assign node1818 = (inp[12]) ? node1820 : 4'b0000;
														assign node1820 = (inp[3]) ? 4'b1000 : 4'b1101;
													assign node1823 = (inp[3]) ? node1825 : 4'b0000;
														assign node1825 = (inp[7]) ? node1827 : 4'b0100;
															assign node1827 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node1830 = (inp[3]) ? node1838 : node1831;
													assign node1831 = (inp[4]) ? node1835 : node1832;
														assign node1832 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node1835 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node1838 = (inp[7]) ? 4'b1000 : node1839;
														assign node1839 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node1843 = (inp[7]) ? node1855 : node1844;
												assign node1844 = (inp[3]) ? node1850 : node1845;
													assign node1845 = (inp[4]) ? node1847 : 4'b0001;
														assign node1847 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1850 = (inp[4]) ? 4'b0101 : node1851;
														assign node1851 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node1855 = (inp[3]) ? node1863 : node1856;
													assign node1856 = (inp[4]) ? node1858 : 4'b1101;
														assign node1858 = (inp[10]) ? 4'b0001 : node1859;
															assign node1859 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node1863 = (inp[4]) ? 4'b1101 : node1864;
														assign node1864 = (inp[12]) ? 4'b1001 : 4'b0001;
							assign node1869 = (inp[2]) ? 4'b1001 : node1870;
								assign node1870 = (inp[3]) ? node1872 : 4'b1001;
									assign node1872 = (inp[4]) ? node1910 : node1873;
										assign node1873 = (inp[7]) ? 4'b1001 : node1874;
											assign node1874 = (inp[10]) ? node1890 : node1875;
												assign node1875 = (inp[13]) ? node1879 : node1876;
													assign node1876 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node1879 = (inp[12]) ? node1887 : node1880;
														assign node1880 = (inp[1]) ? node1884 : node1881;
															assign node1881 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node1884 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1887 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node1890 = (inp[13]) ? node1900 : node1891;
													assign node1891 = (inp[11]) ? 4'b0000 : node1892;
														assign node1892 = (inp[1]) ? 4'b0000 : node1893;
															assign node1893 = (inp[12]) ? 4'b1001 : node1894;
																assign node1894 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node1900 = (inp[14]) ? node1902 : 4'b1000;
														assign node1902 = (inp[11]) ? node1906 : node1903;
															assign node1903 = (inp[12]) ? 4'b0001 : 4'b1000;
															assign node1906 = (inp[1]) ? 4'b1001 : 4'b1000;
										assign node1910 = (inp[1]) ? node1932 : node1911;
											assign node1911 = (inp[11]) ? node1921 : node1912;
												assign node1912 = (inp[14]) ? node1918 : node1913;
													assign node1913 = (inp[10]) ? 4'b0000 : node1914;
														assign node1914 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node1918 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node1921 = (inp[13]) ? node1927 : node1922;
													assign node1922 = (inp[12]) ? node1924 : 4'b0000;
														assign node1924 = (inp[14]) ? 4'b0000 : 4'b1001;
													assign node1927 = (inp[12]) ? node1929 : 4'b1000;
														assign node1929 = (inp[14]) ? 4'b0000 : 4'b1000;
											assign node1932 = (inp[14]) ? node1942 : node1933;
												assign node1933 = (inp[13]) ? node1939 : node1934;
													assign node1934 = (inp[10]) ? 4'b0001 : node1935;
														assign node1935 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node1939 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node1942 = (inp[11]) ? node1950 : node1943;
													assign node1943 = (inp[13]) ? 4'b1000 : node1944;
														assign node1944 = (inp[10]) ? 4'b0000 : node1945;
															assign node1945 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1950 = (inp[12]) ? 4'b0001 : node1951;
														assign node1951 = (inp[13]) ? 4'b1001 : 4'b0001;
					assign node1956 = (inp[3]) ? node2764 : node1957;
						assign node1957 = (inp[1]) ? node2421 : node1958;
							assign node1958 = (inp[2]) ? node2236 : node1959;
								assign node1959 = (inp[13]) ? node2109 : node1960;
									assign node1960 = (inp[12]) ? node2022 : node1961;
										assign node1961 = (inp[0]) ? node1991 : node1962;
											assign node1962 = (inp[11]) ? node1976 : node1963;
												assign node1963 = (inp[7]) ? node1971 : node1964;
													assign node1964 = (inp[15]) ? 4'b0101 : node1965;
														assign node1965 = (inp[14]) ? node1967 : 4'b0000;
															assign node1967 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node1971 = (inp[14]) ? 4'b0001 : node1972;
														assign node1972 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node1976 = (inp[4]) ? node1984 : node1977;
													assign node1977 = (inp[10]) ? 4'b0100 : node1978;
														assign node1978 = (inp[15]) ? node1980 : 4'b0100;
															assign node1980 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1984 = (inp[15]) ? node1986 : 4'b0001;
														assign node1986 = (inp[7]) ? 4'b0101 : node1987;
															assign node1987 = (inp[10]) ? 4'b1000 : 4'b0101;
											assign node1991 = (inp[11]) ? node2009 : node1992;
												assign node1992 = (inp[15]) ? node2002 : node1993;
													assign node1993 = (inp[10]) ? node1997 : node1994;
														assign node1994 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1997 = (inp[7]) ? 4'b1000 : node1998;
															assign node1998 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2002 = (inp[7]) ? node2006 : node2003;
														assign node2003 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node2006 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node2009 = (inp[15]) ? node2015 : node2010;
													assign node2010 = (inp[7]) ? 4'b0001 : node2011;
														assign node2011 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node2015 = (inp[7]) ? node2019 : node2016;
														assign node2016 = (inp[4]) ? 4'b1001 : 4'b0100;
														assign node2019 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node2022 = (inp[10]) ? node2070 : node2023;
											assign node2023 = (inp[0]) ? node2043 : node2024;
												assign node2024 = (inp[11]) ? node2032 : node2025;
													assign node2025 = (inp[15]) ? node2029 : node2026;
														assign node2026 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node2029 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2032 = (inp[14]) ? 4'b0001 : node2033;
														assign node2033 = (inp[7]) ? node2037 : node2034;
															assign node2034 = (inp[15]) ? 4'b0100 : 4'b0001;
															assign node2037 = (inp[4]) ? node2039 : 4'b0000;
																assign node2039 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node2043 = (inp[7]) ? node2057 : node2044;
													assign node2044 = (inp[15]) ? node2050 : node2045;
														assign node2045 = (inp[4]) ? node2047 : 4'b1100;
															assign node2047 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node2050 = (inp[4]) ? node2052 : 4'b1000;
															assign node2052 = (inp[14]) ? node2054 : 4'b1100;
																assign node2054 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node2057 = (inp[4]) ? node2065 : node2058;
														assign node2058 = (inp[15]) ? node2060 : 4'b1100;
															assign node2060 = (inp[11]) ? 4'b1000 : node2061;
																assign node2061 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node2065 = (inp[15]) ? node2067 : 4'b1001;
															assign node2067 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node2070 = (inp[14]) ? node2086 : node2071;
												assign node2071 = (inp[11]) ? node2075 : node2072;
													assign node2072 = (inp[0]) ? 4'b0000 : 4'b1001;
													assign node2075 = (inp[7]) ? node2081 : node2076;
														assign node2076 = (inp[4]) ? node2078 : 4'b0001;
															assign node2078 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node2081 = (inp[4]) ? node2083 : 4'b0000;
															assign node2083 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node2086 = (inp[7]) ? node2098 : node2087;
													assign node2087 = (inp[0]) ? node2093 : node2088;
														assign node2088 = (inp[4]) ? node2090 : 4'b1100;
															assign node2090 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node2093 = (inp[15]) ? 4'b0100 : node2094;
															assign node2094 = (inp[4]) ? 4'b0100 : 4'b0001;
													assign node2098 = (inp[4]) ? node2104 : node2099;
														assign node2099 = (inp[11]) ? 4'b0001 : node2100;
															assign node2100 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node2104 = (inp[15]) ? 4'b0101 : node2105;
															assign node2105 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node2109 = (inp[11]) ? node2173 : node2110;
										assign node2110 = (inp[0]) ? node2134 : node2111;
											assign node2111 = (inp[4]) ? node2125 : node2112;
												assign node2112 = (inp[7]) ? node2116 : node2113;
													assign node2113 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node2116 = (inp[12]) ? node2122 : node2117;
														assign node2117 = (inp[10]) ? 4'b0001 : node2118;
															assign node2118 = (inp[15]) ? 4'b1100 : 4'b0001;
														assign node2122 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node2125 = (inp[7]) ? node2131 : node2126;
													assign node2126 = (inp[15]) ? node2128 : 4'b0000;
														assign node2128 = (inp[10]) ? 4'b1000 : 4'b0001;
													assign node2131 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node2134 = (inp[14]) ? node2162 : node2135;
												assign node2135 = (inp[10]) ? node2157 : node2136;
													assign node2136 = (inp[15]) ? node2150 : node2137;
														assign node2137 = (inp[7]) ? node2143 : node2138;
															assign node2138 = (inp[4]) ? 4'b1001 : node2139;
																assign node2139 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node2143 = (inp[12]) ? node2147 : node2144;
																assign node2144 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node2147 = (inp[4]) ? 4'b1000 : 4'b0100;
														assign node2150 = (inp[12]) ? node2152 : 4'b1100;
															assign node2152 = (inp[7]) ? node2154 : 4'b0100;
																assign node2154 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2157 = (inp[15]) ? 4'b1000 : node2158;
														assign node2158 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node2162 = (inp[4]) ? node2168 : node2163;
													assign node2163 = (inp[12]) ? node2165 : 4'b0000;
														assign node2165 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2168 = (inp[10]) ? 4'b0000 : node2169;
														assign node2169 = (inp[15]) ? 4'b0000 : 4'b0100;
										assign node2173 = (inp[0]) ? node2201 : node2174;
											assign node2174 = (inp[4]) ? node2182 : node2175;
												assign node2175 = (inp[15]) ? 4'b0001 : node2176;
													assign node2176 = (inp[10]) ? 4'b0000 : node2177;
														assign node2177 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node2182 = (inp[12]) ? node2192 : node2183;
													assign node2183 = (inp[14]) ? 4'b0000 : node2184;
														assign node2184 = (inp[7]) ? node2186 : 4'b1001;
															assign node2186 = (inp[15]) ? node2188 : 4'b0000;
																assign node2188 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2192 = (inp[10]) ? node2196 : node2193;
														assign node2193 = (inp[15]) ? 4'b1000 : 4'b0001;
														assign node2196 = (inp[15]) ? 4'b1001 : node2197;
															assign node2197 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node2201 = (inp[10]) ? node2211 : node2202;
												assign node2202 = (inp[4]) ? node2208 : node2203;
													assign node2203 = (inp[15]) ? node2205 : 4'b0001;
														assign node2205 = (inp[14]) ? 4'b1100 : 4'b0000;
													assign node2208 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node2211 = (inp[12]) ? node2229 : node2212;
													assign node2212 = (inp[14]) ? node2220 : node2213;
														assign node2213 = (inp[4]) ? node2217 : node2214;
															assign node2214 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node2217 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node2220 = (inp[7]) ? node2222 : 4'b1001;
															assign node2222 = (inp[15]) ? node2226 : node2223;
																assign node2223 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node2226 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node2229 = (inp[15]) ? node2231 : 4'b0001;
														assign node2231 = (inp[4]) ? 4'b0001 : node2232;
															assign node2232 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node2236 = (inp[0]) ? node2376 : node2237;
									assign node2237 = (inp[4]) ? node2317 : node2238;
										assign node2238 = (inp[11]) ? node2282 : node2239;
											assign node2239 = (inp[13]) ? node2261 : node2240;
												assign node2240 = (inp[7]) ? node2254 : node2241;
													assign node2241 = (inp[15]) ? node2245 : node2242;
														assign node2242 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node2245 = (inp[14]) ? 4'b0100 : node2246;
															assign node2246 = (inp[12]) ? node2250 : node2247;
																assign node2247 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node2250 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node2254 = (inp[15]) ? node2256 : 4'b1100;
														assign node2256 = (inp[12]) ? 4'b1000 : node2257;
															assign node2257 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2261 = (inp[14]) ? node2267 : node2262;
													assign node2262 = (inp[15]) ? 4'b0100 : node2263;
														assign node2263 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2267 = (inp[10]) ? node2273 : node2268;
														assign node2268 = (inp[15]) ? node2270 : 4'b0000;
															assign node2270 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node2273 = (inp[12]) ? node2279 : node2274;
															assign node2274 = (inp[15]) ? 4'b0000 : node2275;
																assign node2275 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node2279 = (inp[15]) ? 4'b0100 : 4'b0000;
											assign node2282 = (inp[15]) ? node2298 : node2283;
												assign node2283 = (inp[13]) ? node2293 : node2284;
													assign node2284 = (inp[12]) ? node2286 : 4'b0000;
														assign node2286 = (inp[7]) ? node2290 : node2287;
															assign node2287 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node2290 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node2293 = (inp[14]) ? 4'b1000 : node2294;
														assign node2294 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node2298 = (inp[7]) ? node2308 : node2299;
													assign node2299 = (inp[13]) ? node2303 : node2300;
														assign node2300 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2303 = (inp[10]) ? node2305 : 4'b1101;
															assign node2305 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2308 = (inp[13]) ? node2314 : node2309;
														assign node2309 = (inp[12]) ? 4'b0001 : node2310;
															assign node2310 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node2314 = (inp[14]) ? 4'b0101 : 4'b1101;
										assign node2317 = (inp[11]) ? node2357 : node2318;
											assign node2318 = (inp[12]) ? node2334 : node2319;
												assign node2319 = (inp[15]) ? node2327 : node2320;
													assign node2320 = (inp[14]) ? node2322 : 4'b0001;
														assign node2322 = (inp[10]) ? 4'b0001 : node2323;
															assign node2323 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node2327 = (inp[14]) ? node2329 : 4'b1001;
														assign node2329 = (inp[7]) ? 4'b1000 : node2330;
															assign node2330 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2334 = (inp[15]) ? node2346 : node2335;
													assign node2335 = (inp[10]) ? node2337 : 4'b1001;
														assign node2337 = (inp[7]) ? node2343 : node2338;
															assign node2338 = (inp[14]) ? 4'b1001 : node2339;
																assign node2339 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node2343 = (inp[13]) ? 4'b1001 : 4'b1100;
													assign node2346 = (inp[13]) ? node2354 : node2347;
														assign node2347 = (inp[7]) ? node2349 : 4'b1001;
															assign node2349 = (inp[10]) ? node2351 : 4'b1100;
																assign node2351 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node2354 = (inp[7]) ? 4'b0001 : 4'b0100;
											assign node2357 = (inp[15]) ? node2367 : node2358;
												assign node2358 = (inp[10]) ? node2364 : node2359;
													assign node2359 = (inp[13]) ? node2361 : 4'b0100;
														assign node2361 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node2364 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node2367 = (inp[13]) ? node2371 : node2368;
													assign node2368 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node2371 = (inp[12]) ? 4'b0001 : node2372;
														assign node2372 = (inp[10]) ? 4'b0001 : 4'b1000;
									assign node2376 = (inp[15]) ? 4'b1001 : node2377;
										assign node2377 = (inp[11]) ? node2405 : node2378;
											assign node2378 = (inp[14]) ? node2388 : node2379;
												assign node2379 = (inp[4]) ? node2385 : node2380;
													assign node2380 = (inp[7]) ? 4'b1101 : node2381;
														assign node2381 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node2385 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node2388 = (inp[13]) ? node2394 : node2389;
													assign node2389 = (inp[12]) ? 4'b1101 : node2390;
														assign node2390 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node2394 = (inp[4]) ? node2400 : node2395;
														assign node2395 = (inp[7]) ? 4'b1101 : node2396;
															assign node2396 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2400 = (inp[12]) ? 4'b0001 : node2401;
															assign node2401 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node2405 = (inp[7]) ? node2415 : node2406;
												assign node2406 = (inp[13]) ? node2410 : node2407;
													assign node2407 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2410 = (inp[12]) ? node2412 : 4'b1000;
														assign node2412 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node2415 = (inp[4]) ? node2417 : 4'b1101;
													assign node2417 = (inp[12]) ? 4'b0000 : 4'b1000;
							assign node2421 = (inp[11]) ? node2603 : node2422;
								assign node2422 = (inp[2]) ? node2508 : node2423;
									assign node2423 = (inp[13]) ? node2467 : node2424;
										assign node2424 = (inp[0]) ? node2446 : node2425;
											assign node2425 = (inp[15]) ? node2437 : node2426;
												assign node2426 = (inp[12]) ? 4'b0001 : node2427;
													assign node2427 = (inp[7]) ? 4'b1100 : node2428;
														assign node2428 = (inp[4]) ? node2430 : 4'b1001;
															assign node2430 = (inp[14]) ? 4'b1000 : node2431;
																assign node2431 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node2437 = (inp[4]) ? node2441 : node2438;
													assign node2438 = (inp[7]) ? 4'b1001 : 4'b0101;
													assign node2441 = (inp[14]) ? node2443 : 4'b0001;
														assign node2443 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node2446 = (inp[14]) ? node2456 : node2447;
												assign node2447 = (inp[7]) ? node2449 : 4'b0000;
													assign node2449 = (inp[12]) ? node2451 : 4'b0101;
														assign node2451 = (inp[10]) ? node2453 : 4'b1001;
															assign node2453 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node2456 = (inp[15]) ? node2462 : node2457;
													assign node2457 = (inp[10]) ? 4'b0001 : node2458;
														assign node2458 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2462 = (inp[10]) ? node2464 : 4'b0000;
														assign node2464 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node2467 = (inp[10]) ? node2497 : node2468;
											assign node2468 = (inp[0]) ? node2482 : node2469;
												assign node2469 = (inp[15]) ? node2477 : node2470;
													assign node2470 = (inp[4]) ? node2474 : node2471;
														assign node2471 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node2474 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2477 = (inp[7]) ? node2479 : 4'b0001;
														assign node2479 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node2482 = (inp[15]) ? node2492 : node2483;
													assign node2483 = (inp[7]) ? node2489 : node2484;
														assign node2484 = (inp[12]) ? node2486 : 4'b0000;
															assign node2486 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node2489 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2492 = (inp[7]) ? 4'b0000 : node2493;
														assign node2493 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node2497 = (inp[0]) ? node2503 : node2498;
												assign node2498 = (inp[4]) ? node2500 : 4'b0101;
													assign node2500 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2503 = (inp[15]) ? 4'b1000 : node2504;
													assign node2504 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node2508 = (inp[0]) ? node2572 : node2509;
										assign node2509 = (inp[4]) ? node2535 : node2510;
											assign node2510 = (inp[14]) ? node2520 : node2511;
												assign node2511 = (inp[13]) ? 4'b0100 : node2512;
													assign node2512 = (inp[7]) ? node2514 : 4'b0000;
														assign node2514 = (inp[15]) ? 4'b0000 : node2515;
															assign node2515 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node2520 = (inp[13]) ? node2524 : node2521;
													assign node2521 = (inp[15]) ? 4'b0100 : 4'b0001;
													assign node2524 = (inp[15]) ? node2530 : node2525;
														assign node2525 = (inp[10]) ? node2527 : 4'b1001;
															assign node2527 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node2530 = (inp[10]) ? node2532 : 4'b0100;
															assign node2532 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2535 = (inp[12]) ? node2555 : node2536;
												assign node2536 = (inp[15]) ? node2546 : node2537;
													assign node2537 = (inp[13]) ? node2539 : 4'b1001;
														assign node2539 = (inp[10]) ? 4'b1000 : node2540;
															assign node2540 = (inp[7]) ? 4'b1001 : node2541;
																assign node2541 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2546 = (inp[13]) ? 4'b1001 : node2547;
														assign node2547 = (inp[14]) ? node2549 : 4'b0000;
															assign node2549 = (inp[7]) ? 4'b0001 : node2550;
																assign node2550 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node2555 = (inp[15]) ? node2561 : node2556;
													assign node2556 = (inp[14]) ? node2558 : 4'b0001;
														assign node2558 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node2561 = (inp[14]) ? node2563 : 4'b0001;
														assign node2563 = (inp[10]) ? node2569 : node2564;
															assign node2564 = (inp[13]) ? node2566 : 4'b0001;
																assign node2566 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node2569 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node2572 = (inp[15]) ? 4'b1001 : node2573;
											assign node2573 = (inp[14]) ? node2587 : node2574;
												assign node2574 = (inp[13]) ? node2580 : node2575;
													assign node2575 = (inp[10]) ? 4'b0001 : node2576;
														assign node2576 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node2580 = (inp[4]) ? node2584 : node2581;
														assign node2581 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node2584 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node2587 = (inp[4]) ? node2593 : node2588;
													assign node2588 = (inp[7]) ? 4'b1101 : node2589;
														assign node2589 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node2593 = (inp[13]) ? node2597 : node2594;
														assign node2594 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node2597 = (inp[12]) ? node2599 : 4'b1000;
															assign node2599 = (inp[10]) ? 4'b1000 : 4'b0000;
								assign node2603 = (inp[10]) ? node2697 : node2604;
									assign node2604 = (inp[4]) ? node2656 : node2605;
										assign node2605 = (inp[0]) ? node2631 : node2606;
											assign node2606 = (inp[2]) ? node2616 : node2607;
												assign node2607 = (inp[7]) ? 4'b0101 : node2608;
													assign node2608 = (inp[13]) ? node2612 : node2609;
														assign node2609 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2612 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node2616 = (inp[15]) ? node2626 : node2617;
													assign node2617 = (inp[13]) ? node2621 : node2618;
														assign node2618 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node2621 = (inp[7]) ? node2623 : 4'b0101;
															assign node2623 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2626 = (inp[7]) ? 4'b0001 : node2627;
														assign node2627 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node2631 = (inp[2]) ? node2647 : node2632;
												assign node2632 = (inp[7]) ? node2640 : node2633;
													assign node2633 = (inp[15]) ? node2635 : 4'b0001;
														assign node2635 = (inp[12]) ? node2637 : 4'b0101;
															assign node2637 = (inp[13]) ? 4'b0101 : 4'b1001;
													assign node2640 = (inp[15]) ? node2644 : node2641;
														assign node2641 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node2644 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2647 = (inp[15]) ? 4'b1001 : node2648;
													assign node2648 = (inp[7]) ? 4'b1101 : node2649;
														assign node2649 = (inp[13]) ? 4'b0001 : node2650;
															assign node2650 = (inp[12]) ? 4'b1101 : 4'b0001;
										assign node2656 = (inp[2]) ? node2680 : node2657;
											assign node2657 = (inp[7]) ? node2661 : node2658;
												assign node2658 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node2661 = (inp[14]) ? node2667 : node2662;
													assign node2662 = (inp[13]) ? node2664 : 4'b1001;
														assign node2664 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2667 = (inp[0]) ? node2675 : node2668;
														assign node2668 = (inp[13]) ? 4'b0001 : node2669;
															assign node2669 = (inp[15]) ? 4'b1001 : node2670;
																assign node2670 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2675 = (inp[12]) ? node2677 : 4'b0101;
															assign node2677 = (inp[15]) ? 4'b1001 : 4'b0001;
											assign node2680 = (inp[7]) ? node2688 : node2681;
												assign node2681 = (inp[15]) ? 4'b1001 : node2682;
													assign node2682 = (inp[12]) ? node2684 : 4'b1001;
														assign node2684 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node2688 = (inp[13]) ? node2692 : node2689;
													assign node2689 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node2692 = (inp[15]) ? node2694 : 4'b1001;
														assign node2694 = (inp[12]) ? 4'b1001 : 4'b0101;
									assign node2697 = (inp[13]) ? node2743 : node2698;
										assign node2698 = (inp[15]) ? node2724 : node2699;
											assign node2699 = (inp[0]) ? node2715 : node2700;
												assign node2700 = (inp[7]) ? node2706 : node2701;
													assign node2701 = (inp[4]) ? 4'b1001 : node2702;
														assign node2702 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node2706 = (inp[14]) ? node2708 : 4'b1001;
														assign node2708 = (inp[2]) ? node2712 : node2709;
															assign node2709 = (inp[4]) ? 4'b0101 : 4'b1001;
															assign node2712 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node2715 = (inp[7]) ? node2721 : node2716;
													assign node2716 = (inp[2]) ? 4'b0001 : node2717;
														assign node2717 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node2721 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node2724 = (inp[0]) ? node2736 : node2725;
												assign node2725 = (inp[7]) ? node2733 : node2726;
													assign node2726 = (inp[2]) ? node2730 : node2727;
														assign node2727 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2730 = (inp[4]) ? 4'b0101 : 4'b1101;
													assign node2733 = (inp[4]) ? 4'b0001 : 4'b1001;
												assign node2736 = (inp[2]) ? 4'b1001 : node2737;
													assign node2737 = (inp[12]) ? 4'b0101 : node2738;
														assign node2738 = (inp[4]) ? 4'b1001 : 4'b0001;
										assign node2743 = (inp[4]) ? 4'b1001 : node2744;
											assign node2744 = (inp[7]) ? node2750 : node2745;
												assign node2745 = (inp[0]) ? node2747 : 4'b1001;
													assign node2747 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node2750 = (inp[15]) ? node2758 : node2751;
													assign node2751 = (inp[0]) ? node2755 : node2752;
														assign node2752 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node2755 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node2758 = (inp[0]) ? 4'b1001 : node2759;
														assign node2759 = (inp[2]) ? 4'b1101 : 4'b1001;
						assign node2764 = (inp[4]) ? node3186 : node2765;
							assign node2765 = (inp[11]) ? node2979 : node2766;
								assign node2766 = (inp[2]) ? node2886 : node2767;
									assign node2767 = (inp[12]) ? node2827 : node2768;
										assign node2768 = (inp[13]) ? node2790 : node2769;
											assign node2769 = (inp[15]) ? node2781 : node2770;
												assign node2770 = (inp[1]) ? node2776 : node2771;
													assign node2771 = (inp[7]) ? 4'b0001 : node2772;
														assign node2772 = (inp[0]) ? 4'b0001 : 4'b1000;
													assign node2776 = (inp[10]) ? 4'b1001 : node2777;
														assign node2777 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node2781 = (inp[7]) ? node2785 : node2782;
													assign node2782 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2785 = (inp[1]) ? 4'b0000 : node2786;
														assign node2786 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node2790 = (inp[7]) ? node2806 : node2791;
												assign node2791 = (inp[10]) ? node2801 : node2792;
													assign node2792 = (inp[1]) ? node2798 : node2793;
														assign node2793 = (inp[0]) ? node2795 : 4'b1001;
															assign node2795 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node2798 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node2801 = (inp[0]) ? 4'b1000 : node2802;
														assign node2802 = (inp[14]) ? 4'b1000 : 4'b0001;
												assign node2806 = (inp[10]) ? node2820 : node2807;
													assign node2807 = (inp[15]) ? node2811 : node2808;
														assign node2808 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node2811 = (inp[0]) ? node2815 : node2812;
															assign node2812 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node2815 = (inp[14]) ? node2817 : 4'b1001;
																assign node2817 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node2820 = (inp[15]) ? node2822 : 4'b1001;
														assign node2822 = (inp[0]) ? node2824 : 4'b0001;
															assign node2824 = (inp[14]) ? 4'b0001 : 4'b1001;
										assign node2827 = (inp[7]) ? node2861 : node2828;
											assign node2828 = (inp[1]) ? node2850 : node2829;
												assign node2829 = (inp[0]) ? node2843 : node2830;
													assign node2830 = (inp[15]) ? node2836 : node2831;
														assign node2831 = (inp[14]) ? node2833 : 4'b0000;
															assign node2833 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2836 = (inp[13]) ? node2840 : node2837;
															assign node2837 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node2840 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node2843 = (inp[10]) ? 4'b1001 : node2844;
														assign node2844 = (inp[14]) ? 4'b1000 : node2845;
															assign node2845 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node2850 = (inp[15]) ? node2858 : node2851;
													assign node2851 = (inp[13]) ? node2853 : 4'b0001;
														assign node2853 = (inp[14]) ? 4'b0001 : node2854;
															assign node2854 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2858 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node2861 = (inp[14]) ? node2877 : node2862;
												assign node2862 = (inp[15]) ? node2864 : 4'b1001;
													assign node2864 = (inp[0]) ? node2874 : node2865;
														assign node2865 = (inp[10]) ? node2871 : node2866;
															assign node2866 = (inp[13]) ? node2868 : 4'b0000;
																assign node2868 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node2871 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node2874 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node2877 = (inp[13]) ? 4'b0000 : node2878;
													assign node2878 = (inp[15]) ? node2880 : 4'b1000;
														assign node2880 = (inp[10]) ? node2882 : 4'b0000;
															assign node2882 = (inp[1]) ? 4'b1000 : 4'b0000;
									assign node2886 = (inp[7]) ? node2942 : node2887;
										assign node2887 = (inp[10]) ? node2911 : node2888;
											assign node2888 = (inp[0]) ? node2906 : node2889;
												assign node2889 = (inp[1]) ? node2899 : node2890;
													assign node2890 = (inp[14]) ? node2892 : 4'b0000;
														assign node2892 = (inp[12]) ? node2894 : 4'b0000;
															assign node2894 = (inp[15]) ? node2896 : 4'b0000;
																assign node2896 = (inp[13]) ? 4'b0000 : 4'b1001;
													assign node2899 = (inp[13]) ? 4'b0001 : node2900;
														assign node2900 = (inp[12]) ? 4'b1000 : node2901;
															assign node2901 = (inp[15]) ? 4'b1000 : 4'b0000;
												assign node2906 = (inp[14]) ? 4'b0000 : node2907;
													assign node2907 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node2911 = (inp[12]) ? node2929 : node2912;
												assign node2912 = (inp[13]) ? node2924 : node2913;
													assign node2913 = (inp[0]) ? node2917 : node2914;
														assign node2914 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node2917 = (inp[15]) ? node2919 : 4'b1000;
															assign node2919 = (inp[14]) ? 4'b0001 : node2920;
																assign node2920 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node2924 = (inp[15]) ? node2926 : 4'b1001;
														assign node2926 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node2929 = (inp[13]) ? node2937 : node2930;
													assign node2930 = (inp[15]) ? 4'b0000 : node2931;
														assign node2931 = (inp[14]) ? 4'b1000 : node2932;
															assign node2932 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node2937 = (inp[15]) ? node2939 : 4'b0000;
														assign node2939 = (inp[14]) ? 4'b1000 : 4'b0001;
										assign node2942 = (inp[15]) ? node2968 : node2943;
											assign node2943 = (inp[14]) ? node2955 : node2944;
												assign node2944 = (inp[1]) ? node2948 : node2945;
													assign node2945 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node2948 = (inp[13]) ? node2952 : node2949;
														assign node2949 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2952 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node2955 = (inp[1]) ? node2965 : node2956;
													assign node2956 = (inp[12]) ? node2958 : 4'b1000;
														assign node2958 = (inp[13]) ? node2960 : 4'b1001;
															assign node2960 = (inp[0]) ? 4'b0001 : node2961;
																assign node2961 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node2965 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node2968 = (inp[0]) ? 4'b1001 : node2969;
												assign node2969 = (inp[13]) ? node2975 : node2970;
													assign node2970 = (inp[10]) ? 4'b0000 : node2971;
														assign node2971 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node2975 = (inp[12]) ? 4'b1000 : 4'b0000;
								assign node2979 = (inp[1]) ? node3105 : node2980;
									assign node2980 = (inp[2]) ? node3036 : node2981;
										assign node2981 = (inp[14]) ? node3019 : node2982;
											assign node2982 = (inp[10]) ? node3002 : node2983;
												assign node2983 = (inp[15]) ? node2989 : node2984;
													assign node2984 = (inp[0]) ? node2986 : 4'b1000;
														assign node2986 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2989 = (inp[0]) ? node2997 : node2990;
														assign node2990 = (inp[12]) ? node2992 : 4'b1000;
															assign node2992 = (inp[7]) ? node2994 : 4'b1000;
																assign node2994 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node2997 = (inp[12]) ? node2999 : 4'b0001;
															assign node2999 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node3002 = (inp[13]) ? node3012 : node3003;
													assign node3003 = (inp[15]) ? node3007 : node3004;
														assign node3004 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node3007 = (inp[0]) ? node3009 : 4'b1001;
															assign node3009 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node3012 = (inp[12]) ? 4'b0000 : node3013;
														assign node3013 = (inp[7]) ? 4'b0001 : node3014;
															assign node3014 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node3019 = (inp[0]) ? 4'b0001 : node3020;
												assign node3020 = (inp[12]) ? node3026 : node3021;
													assign node3021 = (inp[15]) ? 4'b1000 : node3022;
														assign node3022 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node3026 = (inp[7]) ? node3030 : node3027;
														assign node3027 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node3030 = (inp[13]) ? 4'b0000 : node3031;
															assign node3031 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node3036 = (inp[12]) ? node3076 : node3037;
											assign node3037 = (inp[13]) ? node3051 : node3038;
												assign node3038 = (inp[7]) ? node3042 : node3039;
													assign node3039 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node3042 = (inp[15]) ? node3048 : node3043;
														assign node3043 = (inp[10]) ? node3045 : 4'b1000;
															assign node3045 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3048 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node3051 = (inp[14]) ? node3057 : node3052;
													assign node3052 = (inp[0]) ? node3054 : 4'b1001;
														assign node3054 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3057 = (inp[0]) ? node3069 : node3058;
														assign node3058 = (inp[7]) ? node3062 : node3059;
															assign node3059 = (inp[15]) ? 4'b0000 : 4'b1001;
															assign node3062 = (inp[15]) ? node3066 : node3063;
																assign node3063 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node3066 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node3069 = (inp[15]) ? node3073 : node3070;
															assign node3070 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node3073 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node3076 = (inp[15]) ? node3094 : node3077;
												assign node3077 = (inp[0]) ? node3083 : node3078;
													assign node3078 = (inp[14]) ? 4'b1001 : node3079;
														assign node3079 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node3083 = (inp[14]) ? 4'b0000 : node3084;
														assign node3084 = (inp[10]) ? node3086 : 4'b0000;
															assign node3086 = (inp[7]) ? node3090 : node3087;
																assign node3087 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node3090 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node3094 = (inp[14]) ? node3102 : node3095;
													assign node3095 = (inp[0]) ? 4'b1001 : node3096;
														assign node3096 = (inp[10]) ? node3098 : 4'b0001;
															assign node3098 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node3102 = (inp[7]) ? 4'b1000 : 4'b0000;
									assign node3105 = (inp[13]) ? node3163 : node3106;
										assign node3106 = (inp[10]) ? node3130 : node3107;
											assign node3107 = (inp[15]) ? node3115 : node3108;
												assign node3108 = (inp[2]) ? 4'b0001 : node3109;
													assign node3109 = (inp[0]) ? node3111 : 4'b1001;
														assign node3111 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3115 = (inp[14]) ? node3123 : node3116;
													assign node3116 = (inp[2]) ? node3120 : node3117;
														assign node3117 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3120 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node3123 = (inp[12]) ? 4'b0001 : node3124;
														assign node3124 = (inp[0]) ? 4'b1001 : node3125;
															assign node3125 = (inp[2]) ? 4'b0001 : 4'b1001;
											assign node3130 = (inp[7]) ? node3142 : node3131;
												assign node3131 = (inp[0]) ? 4'b0001 : node3132;
													assign node3132 = (inp[14]) ? 4'b0001 : node3133;
														assign node3133 = (inp[15]) ? node3137 : node3134;
															assign node3134 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node3137 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node3142 = (inp[0]) ? node3148 : node3143;
													assign node3143 = (inp[12]) ? 4'b0001 : node3144;
														assign node3144 = (inp[15]) ? 4'b1001 : 4'b0001;
													assign node3148 = (inp[14]) ? node3154 : node3149;
														assign node3149 = (inp[2]) ? node3151 : 4'b1001;
															assign node3151 = (inp[15]) ? 4'b1001 : 4'b0001;
														assign node3154 = (inp[12]) ? node3158 : node3155;
															assign node3155 = (inp[15]) ? 4'b0001 : 4'b1001;
															assign node3158 = (inp[2]) ? node3160 : 4'b0001;
																assign node3160 = (inp[15]) ? 4'b1001 : 4'b0001;
										assign node3163 = (inp[10]) ? 4'b1001 : node3164;
											assign node3164 = (inp[0]) ? node3172 : node3165;
												assign node3165 = (inp[14]) ? node3167 : 4'b0001;
													assign node3167 = (inp[7]) ? 4'b0001 : node3168;
														assign node3168 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node3172 = (inp[15]) ? node3178 : node3173;
													assign node3173 = (inp[7]) ? node3175 : 4'b0001;
														assign node3175 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node3178 = (inp[14]) ? node3180 : 4'b1001;
														assign node3180 = (inp[2]) ? node3182 : 4'b1001;
															assign node3182 = (inp[7]) ? 4'b1001 : 4'b0001;
							assign node3186 = (inp[13]) ? node3392 : node3187;
								assign node3187 = (inp[1]) ? node3291 : node3188;
									assign node3188 = (inp[10]) ? node3228 : node3189;
										assign node3189 = (inp[0]) ? node3207 : node3190;
											assign node3190 = (inp[15]) ? node3200 : node3191;
												assign node3191 = (inp[11]) ? node3195 : node3192;
													assign node3192 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node3195 = (inp[14]) ? 4'b0001 : node3196;
														assign node3196 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node3200 = (inp[2]) ? node3202 : 4'b1000;
													assign node3202 = (inp[12]) ? 4'b0000 : node3203;
														assign node3203 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node3207 = (inp[14]) ? node3213 : node3208;
												assign node3208 = (inp[7]) ? node3210 : 4'b0000;
													assign node3210 = (inp[15]) ? 4'b0000 : 4'b1000;
												assign node3213 = (inp[12]) ? node3219 : node3214;
													assign node3214 = (inp[7]) ? 4'b0001 : node3215;
														assign node3215 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node3219 = (inp[2]) ? node3221 : 4'b0000;
														assign node3221 = (inp[11]) ? node3225 : node3222;
															assign node3222 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node3225 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node3228 = (inp[15]) ? node3264 : node3229;
											assign node3229 = (inp[2]) ? node3251 : node3230;
												assign node3230 = (inp[7]) ? node3240 : node3231;
													assign node3231 = (inp[14]) ? node3235 : node3232;
														assign node3232 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node3235 = (inp[0]) ? node3237 : 4'b0000;
															assign node3237 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3240 = (inp[14]) ? node3246 : node3241;
														assign node3241 = (inp[0]) ? 4'b0000 : node3242;
															assign node3242 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3246 = (inp[11]) ? node3248 : 4'b0001;
															assign node3248 = (inp[12]) ? 4'b0001 : 4'b1000;
												assign node3251 = (inp[11]) ? node3259 : node3252;
													assign node3252 = (inp[0]) ? 4'b0001 : node3253;
														assign node3253 = (inp[12]) ? node3255 : 4'b1001;
															assign node3255 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node3259 = (inp[14]) ? node3261 : 4'b1000;
														assign node3261 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node3264 = (inp[0]) ? node3278 : node3265;
												assign node3265 = (inp[2]) ? node3271 : node3266;
													assign node3266 = (inp[12]) ? node3268 : 4'b0001;
														assign node3268 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node3271 = (inp[7]) ? node3273 : 4'b0000;
														assign node3273 = (inp[12]) ? node3275 : 4'b0001;
															assign node3275 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node3278 = (inp[7]) ? node3280 : 4'b1000;
													assign node3280 = (inp[2]) ? 4'b0000 : node3281;
														assign node3281 = (inp[14]) ? node3287 : node3282;
															assign node3282 = (inp[11]) ? node3284 : 4'b1000;
																assign node3284 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node3287 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node3291 = (inp[11]) ? node3355 : node3292;
										assign node3292 = (inp[10]) ? node3322 : node3293;
											assign node3293 = (inp[0]) ? node3309 : node3294;
												assign node3294 = (inp[15]) ? node3300 : node3295;
													assign node3295 = (inp[7]) ? 4'b0000 : node3296;
														assign node3296 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node3300 = (inp[14]) ? 4'b1001 : node3301;
														assign node3301 = (inp[7]) ? node3303 : 4'b0001;
															assign node3303 = (inp[12]) ? 4'b1000 : node3304;
																assign node3304 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node3309 = (inp[12]) ? node3313 : node3310;
													assign node3310 = (inp[15]) ? 4'b0000 : 4'b1001;
													assign node3313 = (inp[7]) ? node3315 : 4'b0000;
														assign node3315 = (inp[15]) ? 4'b1001 : node3316;
															assign node3316 = (inp[2]) ? node3318 : 4'b0001;
																assign node3318 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node3322 = (inp[15]) ? node3338 : node3323;
												assign node3323 = (inp[14]) ? node3333 : node3324;
													assign node3324 = (inp[7]) ? node3330 : node3325;
														assign node3325 = (inp[12]) ? 4'b0001 : node3326;
															assign node3326 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node3330 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node3333 = (inp[7]) ? 4'b0000 : node3334;
														assign node3334 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3338 = (inp[12]) ? node3348 : node3339;
													assign node3339 = (inp[14]) ? node3341 : 4'b0001;
														assign node3341 = (inp[7]) ? node3343 : 4'b0001;
															assign node3343 = (inp[0]) ? 4'b0001 : node3344;
																assign node3344 = (inp[2]) ? 4'b0001 : 4'b1000;
													assign node3348 = (inp[14]) ? node3352 : node3349;
														assign node3349 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node3352 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node3355 = (inp[10]) ? 4'b0001 : node3356;
											assign node3356 = (inp[2]) ? node3376 : node3357;
												assign node3357 = (inp[12]) ? node3363 : node3358;
													assign node3358 = (inp[7]) ? 4'b0001 : node3359;
														assign node3359 = (inp[15]) ? 4'b1001 : 4'b0001;
													assign node3363 = (inp[15]) ? node3369 : node3364;
														assign node3364 = (inp[14]) ? node3366 : 4'b1001;
															assign node3366 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node3369 = (inp[14]) ? 4'b1001 : node3370;
															assign node3370 = (inp[7]) ? node3372 : 4'b0001;
																assign node3372 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node3376 = (inp[15]) ? 4'b0001 : node3377;
													assign node3377 = (inp[0]) ? node3383 : node3378;
														assign node3378 = (inp[7]) ? 4'b0001 : node3379;
															assign node3379 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3383 = (inp[14]) ? node3387 : node3384;
															assign node3384 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node3387 = (inp[12]) ? 4'b0001 : 4'b1001;
								assign node3392 = (inp[10]) ? node3472 : node3393;
									assign node3393 = (inp[11]) ? node3443 : node3394;
										assign node3394 = (inp[0]) ? node3416 : node3395;
											assign node3395 = (inp[15]) ? node3409 : node3396;
												assign node3396 = (inp[1]) ? 4'b0000 : node3397;
													assign node3397 = (inp[7]) ? node3405 : node3398;
														assign node3398 = (inp[14]) ? 4'b0000 : node3399;
															assign node3399 = (inp[12]) ? node3401 : 4'b0001;
																assign node3401 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node3405 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node3409 = (inp[1]) ? node3411 : 4'b0000;
													assign node3411 = (inp[14]) ? 4'b0001 : node3412;
														assign node3412 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node3416 = (inp[15]) ? node3432 : node3417;
												assign node3417 = (inp[7]) ? node3419 : 4'b0001;
													assign node3419 = (inp[14]) ? node3427 : node3420;
														assign node3420 = (inp[1]) ? node3424 : node3421;
															assign node3421 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node3424 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node3427 = (inp[1]) ? node3429 : 4'b0000;
															assign node3429 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node3432 = (inp[1]) ? 4'b0000 : node3433;
													assign node3433 = (inp[14]) ? node3437 : node3434;
														assign node3434 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node3437 = (inp[7]) ? node3439 : 4'b0001;
															assign node3439 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node3443 = (inp[1]) ? 4'b0001 : node3444;
											assign node3444 = (inp[14]) ? node3460 : node3445;
												assign node3445 = (inp[7]) ? node3453 : node3446;
													assign node3446 = (inp[2]) ? node3448 : 4'b0001;
														assign node3448 = (inp[0]) ? node3450 : 4'b0000;
															assign node3450 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node3453 = (inp[2]) ? node3455 : 4'b0000;
														assign node3455 = (inp[15]) ? 4'b0001 : node3456;
															assign node3456 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node3460 = (inp[7]) ? 4'b0000 : node3461;
													assign node3461 = (inp[2]) ? node3463 : 4'b0001;
														assign node3463 = (inp[0]) ? node3465 : 4'b0000;
															assign node3465 = (inp[15]) ? node3467 : 4'b0000;
																assign node3467 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node3472 = (inp[11]) ? 4'b0000 : node3473;
										assign node3473 = (inp[1]) ? 4'b0000 : node3474;
											assign node3474 = (inp[0]) ? node3486 : node3475;
												assign node3475 = (inp[7]) ? node3481 : node3476;
													assign node3476 = (inp[2]) ? node3478 : 4'b0001;
														assign node3478 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node3481 = (inp[2]) ? 4'b0000 : node3482;
														assign node3482 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node3486 = (inp[14]) ? node3488 : 4'b0000;
													assign node3488 = (inp[12]) ? node3490 : 4'b0000;
														assign node3490 = (inp[15]) ? node3492 : 4'b0000;
															assign node3492 = (inp[7]) ? 4'b0001 : 4'b0000;
			assign node3497 = (inp[15]) ? node5271 : node3498;
				assign node3498 = (inp[6]) ? node3982 : node3499;
					assign node3499 = (inp[0]) ? 4'b0101 : node3500;
						assign node3500 = (inp[2]) ? node3820 : node3501;
							assign node3501 = (inp[1]) ? node3651 : node3502;
								assign node3502 = (inp[3]) ? node3582 : node3503;
									assign node3503 = (inp[5]) ? node3537 : node3504;
										assign node3504 = (inp[13]) ? node3516 : node3505;
											assign node3505 = (inp[4]) ? node3507 : 4'b0111;
												assign node3507 = (inp[7]) ? 4'b0111 : node3508;
													assign node3508 = (inp[11]) ? node3510 : 4'b0000;
														assign node3510 = (inp[14]) ? node3512 : 4'b1000;
															assign node3512 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3516 = (inp[12]) ? node3522 : node3517;
												assign node3517 = (inp[14]) ? node3519 : 4'b0000;
													assign node3519 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node3522 = (inp[7]) ? node3530 : node3523;
													assign node3523 = (inp[4]) ? node3527 : node3524;
														assign node3524 = (inp[10]) ? 4'b0000 : 4'b0111;
														assign node3527 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node3530 = (inp[10]) ? node3532 : 4'b0111;
														assign node3532 = (inp[4]) ? node3534 : 4'b0111;
															assign node3534 = (inp[14]) ? 4'b0111 : 4'b0000;
										assign node3537 = (inp[4]) ? node3565 : node3538;
											assign node3538 = (inp[11]) ? node3554 : node3539;
												assign node3539 = (inp[14]) ? node3543 : node3540;
													assign node3540 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node3543 = (inp[7]) ? node3545 : 4'b1101;
														assign node3545 = (inp[10]) ? node3547 : 4'b0101;
															assign node3547 = (inp[12]) ? node3551 : node3548;
																assign node3548 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node3551 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node3554 = (inp[13]) ? node3560 : node3555;
													assign node3555 = (inp[10]) ? 4'b1100 : node3556;
														assign node3556 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node3560 = (inp[12]) ? 4'b1100 : node3561;
														assign node3561 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node3565 = (inp[7]) ? node3571 : node3566;
												assign node3566 = (inp[11]) ? 4'b1000 : node3567;
													assign node3567 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node3571 = (inp[13]) ? node3579 : node3572;
													assign node3572 = (inp[10]) ? 4'b1100 : node3573;
														assign node3573 = (inp[11]) ? node3575 : 4'b0101;
															assign node3575 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node3579 = (inp[10]) ? 4'b0000 : 4'b1101;
									assign node3582 = (inp[11]) ? node3624 : node3583;
										assign node3583 = (inp[14]) ? node3599 : node3584;
											assign node3584 = (inp[13]) ? node3592 : node3585;
												assign node3585 = (inp[12]) ? node3587 : 4'b1000;
													assign node3587 = (inp[7]) ? node3589 : 4'b1100;
														assign node3589 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node3592 = (inp[10]) ? node3596 : node3593;
													assign node3593 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node3596 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node3599 = (inp[13]) ? node3613 : node3600;
												assign node3600 = (inp[7]) ? node3608 : node3601;
													assign node3601 = (inp[4]) ? node3603 : 4'b0001;
														assign node3603 = (inp[5]) ? 4'b0101 : node3604;
															assign node3604 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node3608 = (inp[12]) ? 4'b0001 : node3609;
														assign node3609 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3613 = (inp[10]) ? node3619 : node3614;
													assign node3614 = (inp[4]) ? node3616 : 4'b1001;
														assign node3616 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3619 = (inp[12]) ? 4'b1001 : node3620;
														assign node3620 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node3624 = (inp[13]) ? node3638 : node3625;
											assign node3625 = (inp[10]) ? node3633 : node3626;
												assign node3626 = (inp[12]) ? node3628 : 4'b1000;
													assign node3628 = (inp[7]) ? 4'b0000 : node3629;
														assign node3629 = (inp[14]) ? 4'b0000 : 4'b0100;
												assign node3633 = (inp[7]) ? 4'b1000 : node3634;
													assign node3634 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node3638 = (inp[4]) ? node3644 : node3639;
												assign node3639 = (inp[12]) ? 4'b1000 : node3640;
													assign node3640 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node3644 = (inp[10]) ? 4'b0100 : node3645;
													assign node3645 = (inp[12]) ? node3647 : 4'b0100;
														assign node3647 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node3651 = (inp[11]) ? node3751 : node3652;
									assign node3652 = (inp[14]) ? node3704 : node3653;
										assign node3653 = (inp[7]) ? node3679 : node3654;
											assign node3654 = (inp[3]) ? node3666 : node3655;
												assign node3655 = (inp[13]) ? node3663 : node3656;
													assign node3656 = (inp[4]) ? node3658 : 4'b1101;
														assign node3658 = (inp[5]) ? node3660 : 4'b1001;
															assign node3660 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3663 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node3666 = (inp[4]) ? node3672 : node3667;
													assign node3667 = (inp[10]) ? 4'b1001 : node3668;
														assign node3668 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3672 = (inp[5]) ? 4'b1101 : node3673;
														assign node3673 = (inp[10]) ? 4'b0101 : node3674;
															assign node3674 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node3679 = (inp[3]) ? node3691 : node3680;
												assign node3680 = (inp[5]) ? node3686 : node3681;
													assign node3681 = (inp[13]) ? node3683 : 4'b0111;
														assign node3683 = (inp[4]) ? 4'b0001 : 4'b0111;
													assign node3686 = (inp[13]) ? 4'b1101 : node3687;
														assign node3687 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node3691 = (inp[5]) ? node3697 : node3692;
													assign node3692 = (inp[12]) ? node3694 : 4'b1001;
														assign node3694 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3697 = (inp[10]) ? node3701 : node3698;
														assign node3698 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node3701 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node3704 = (inp[13]) ? node3730 : node3705;
											assign node3705 = (inp[10]) ? node3719 : node3706;
												assign node3706 = (inp[7]) ? node3714 : node3707;
													assign node3707 = (inp[12]) ? node3709 : 4'b1000;
														assign node3709 = (inp[3]) ? node3711 : 4'b0000;
															assign node3711 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node3714 = (inp[5]) ? node3716 : 4'b0111;
														assign node3716 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node3719 = (inp[4]) ? node3725 : node3720;
													assign node3720 = (inp[3]) ? 4'b1000 : node3721;
														assign node3721 = (inp[12]) ? 4'b0111 : 4'b1100;
													assign node3725 = (inp[3]) ? node3727 : 4'b1000;
														assign node3727 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node3730 = (inp[12]) ? node3738 : node3731;
												assign node3731 = (inp[3]) ? node3733 : 4'b0000;
													assign node3733 = (inp[7]) ? node3735 : 4'b0100;
														assign node3735 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node3738 = (inp[10]) ? node3744 : node3739;
													assign node3739 = (inp[3]) ? node3741 : 4'b1100;
														assign node3741 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node3744 = (inp[3]) ? 4'b0100 : node3745;
														assign node3745 = (inp[5]) ? node3747 : 4'b0111;
															assign node3747 = (inp[7]) ? 4'b0100 : 4'b0000;
									assign node3751 = (inp[13]) ? node3783 : node3752;
										assign node3752 = (inp[3]) ? node3770 : node3753;
											assign node3753 = (inp[7]) ? node3763 : node3754;
												assign node3754 = (inp[4]) ? node3758 : node3755;
													assign node3755 = (inp[5]) ? 4'b1101 : 4'b0111;
													assign node3758 = (inp[10]) ? 4'b1001 : node3759;
														assign node3759 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3763 = (inp[5]) ? node3765 : 4'b0111;
													assign node3765 = (inp[4]) ? node3767 : 4'b1101;
														assign node3767 = (inp[14]) ? 4'b0101 : 4'b1101;
											assign node3770 = (inp[4]) ? node3776 : node3771;
												assign node3771 = (inp[10]) ? 4'b1001 : node3772;
													assign node3772 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3776 = (inp[7]) ? 4'b1001 : node3777;
													assign node3777 = (inp[12]) ? node3779 : 4'b1101;
														assign node3779 = (inp[10]) ? 4'b1101 : 4'b0101;
										assign node3783 = (inp[12]) ? node3797 : node3784;
											assign node3784 = (inp[3]) ? node3792 : node3785;
												assign node3785 = (inp[4]) ? 4'b0001 : node3786;
													assign node3786 = (inp[7]) ? node3788 : 4'b0001;
														assign node3788 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node3792 = (inp[7]) ? node3794 : 4'b0101;
													assign node3794 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node3797 = (inp[10]) ? node3813 : node3798;
												assign node3798 = (inp[5]) ? node3804 : node3799;
													assign node3799 = (inp[3]) ? node3801 : 4'b0111;
														assign node3801 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3804 = (inp[4]) ? node3806 : 4'b1001;
														assign node3806 = (inp[7]) ? node3810 : node3807;
															assign node3807 = (inp[14]) ? 4'b1001 : 4'b1101;
															assign node3810 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node3813 = (inp[3]) ? node3815 : 4'b0001;
													assign node3815 = (inp[4]) ? 4'b0101 : node3816;
														assign node3816 = (inp[7]) ? 4'b0001 : 4'b0101;
							assign node3820 = (inp[5]) ? node3822 : 4'b0111;
								assign node3822 = (inp[3]) ? node3878 : node3823;
									assign node3823 = (inp[7]) ? node3861 : node3824;
										assign node3824 = (inp[4]) ? node3836 : node3825;
											assign node3825 = (inp[13]) ? node3827 : 4'b0111;
												assign node3827 = (inp[1]) ? node3833 : node3828;
													assign node3828 = (inp[14]) ? node3830 : 4'b0000;
														assign node3830 = (inp[10]) ? 4'b0000 : 4'b0111;
													assign node3833 = (inp[12]) ? 4'b0111 : 4'b0001;
											assign node3836 = (inp[1]) ? node3850 : node3837;
												assign node3837 = (inp[11]) ? node3841 : node3838;
													assign node3838 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node3841 = (inp[13]) ? node3847 : node3842;
														assign node3842 = (inp[12]) ? node3844 : 4'b1000;
															assign node3844 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3847 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node3850 = (inp[14]) ? node3856 : node3851;
													assign node3851 = (inp[13]) ? 4'b1001 : node3852;
														assign node3852 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3856 = (inp[13]) ? node3858 : 4'b1001;
														assign node3858 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node3861 = (inp[4]) ? node3863 : 4'b0111;
											assign node3863 = (inp[13]) ? node3865 : 4'b0111;
												assign node3865 = (inp[10]) ? node3873 : node3866;
													assign node3866 = (inp[12]) ? 4'b0111 : node3867;
														assign node3867 = (inp[11]) ? node3869 : 4'b0111;
															assign node3869 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node3873 = (inp[1]) ? 4'b0001 : node3874;
														assign node3874 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node3878 = (inp[4]) ? node3924 : node3879;
										assign node3879 = (inp[13]) ? node3895 : node3880;
											assign node3880 = (inp[10]) ? node3888 : node3881;
												assign node3881 = (inp[11]) ? node3885 : node3882;
													assign node3882 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node3885 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3888 = (inp[14]) ? node3890 : 4'b1000;
													assign node3890 = (inp[1]) ? node3892 : 4'b1001;
														assign node3892 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node3895 = (inp[12]) ? node3911 : node3896;
												assign node3896 = (inp[7]) ? node3900 : node3897;
													assign node3897 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node3900 = (inp[10]) ? node3906 : node3901;
														assign node3901 = (inp[1]) ? node3903 : 4'b0000;
															assign node3903 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3906 = (inp[1]) ? 4'b0001 : node3907;
															assign node3907 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node3911 = (inp[10]) ? node3919 : node3912;
													assign node3912 = (inp[11]) ? node3916 : node3913;
														assign node3913 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node3916 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node3919 = (inp[11]) ? node3921 : 4'b0100;
														assign node3921 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node3924 = (inp[7]) ? node3956 : node3925;
											assign node3925 = (inp[1]) ? node3943 : node3926;
												assign node3926 = (inp[11]) ? node3936 : node3927;
													assign node3927 = (inp[14]) ? node3931 : node3928;
														assign node3928 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node3931 = (inp[12]) ? node3933 : 4'b1101;
															assign node3933 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node3936 = (inp[14]) ? node3938 : 4'b1100;
														assign node3938 = (inp[13]) ? node3940 : 4'b0100;
															assign node3940 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node3943 = (inp[14]) ? node3951 : node3944;
													assign node3944 = (inp[10]) ? 4'b0101 : node3945;
														assign node3945 = (inp[12]) ? node3947 : 4'b1101;
															assign node3947 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node3951 = (inp[12]) ? node3953 : 4'b1100;
														assign node3953 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node3956 = (inp[13]) ? node3970 : node3957;
												assign node3957 = (inp[10]) ? node3967 : node3958;
													assign node3958 = (inp[12]) ? node3960 : 4'b1000;
														assign node3960 = (inp[1]) ? node3964 : node3961;
															assign node3961 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node3964 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node3967 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node3970 = (inp[12]) ? 4'b1001 : node3971;
													assign node3971 = (inp[10]) ? 4'b0100 : node3972;
														assign node3972 = (inp[14]) ? node3976 : node3973;
															assign node3973 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node3976 = (inp[1]) ? 4'b0100 : 4'b1001;
					assign node3982 = (inp[5]) ? node4560 : node3983;
						assign node3983 = (inp[0]) ? node4413 : node3984;
							assign node3984 = (inp[11]) ? node4206 : node3985;
								assign node3985 = (inp[3]) ? node4103 : node3986;
									assign node3986 = (inp[4]) ? node4050 : node3987;
										assign node3987 = (inp[10]) ? node4023 : node3988;
											assign node3988 = (inp[7]) ? node4006 : node3989;
												assign node3989 = (inp[2]) ? node3997 : node3990;
													assign node3990 = (inp[13]) ? node3994 : node3991;
														assign node3991 = (inp[12]) ? 4'b0101 : 4'b1100;
														assign node3994 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node3997 = (inp[13]) ? node3999 : 4'b1100;
														assign node3999 = (inp[12]) ? node4001 : 4'b1101;
															assign node4001 = (inp[14]) ? 4'b1100 : node4002;
																assign node4002 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node4006 = (inp[2]) ? node4014 : node4007;
													assign node4007 = (inp[13]) ? node4009 : 4'b0101;
														assign node4009 = (inp[14]) ? 4'b1101 : node4010;
															assign node4010 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node4014 = (inp[12]) ? node4018 : node4015;
														assign node4015 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node4018 = (inp[13]) ? 4'b1101 : node4019;
															assign node4019 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node4023 = (inp[7]) ? node4037 : node4024;
												assign node4024 = (inp[13]) ? node4032 : node4025;
													assign node4025 = (inp[2]) ? node4029 : node4026;
														assign node4026 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node4029 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node4032 = (inp[14]) ? 4'b0000 : node4033;
														assign node4033 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node4037 = (inp[2]) ? node4043 : node4038;
													assign node4038 = (inp[13]) ? node4040 : 4'b1101;
														assign node4040 = (inp[1]) ? 4'b0000 : 4'b1101;
													assign node4043 = (inp[14]) ? node4047 : node4044;
														assign node4044 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node4047 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node4050 = (inp[2]) ? node4070 : node4051;
											assign node4051 = (inp[12]) ? node4063 : node4052;
												assign node4052 = (inp[10]) ? node4058 : node4053;
													assign node4053 = (inp[13]) ? node4055 : 4'b1000;
														assign node4055 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node4058 = (inp[13]) ? 4'b0100 : node4059;
														assign node4059 = (inp[14]) ? 4'b0000 : 4'b0100;
												assign node4063 = (inp[10]) ? node4067 : node4064;
													assign node4064 = (inp[1]) ? 4'b1100 : 4'b0000;
													assign node4067 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node4070 = (inp[7]) ? node4084 : node4071;
												assign node4071 = (inp[13]) ? node4075 : node4072;
													assign node4072 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4075 = (inp[12]) ? node4081 : node4076;
														assign node4076 = (inp[10]) ? 4'b0000 : node4077;
															assign node4077 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4081 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node4084 = (inp[13]) ? node4096 : node4085;
													assign node4085 = (inp[10]) ? node4093 : node4086;
														assign node4086 = (inp[12]) ? node4088 : 4'b1100;
															assign node4088 = (inp[1]) ? 4'b0100 : node4089;
																assign node4089 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node4093 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node4096 = (inp[10]) ? 4'b0000 : node4097;
														assign node4097 = (inp[12]) ? node4099 : 4'b0001;
															assign node4099 = (inp[1]) ? 4'b1101 : 4'b1100;
									assign node4103 = (inp[7]) ? node4147 : node4104;
										assign node4104 = (inp[4]) ? node4126 : node4105;
											assign node4105 = (inp[10]) ? node4117 : node4106;
												assign node4106 = (inp[2]) ? node4114 : node4107;
													assign node4107 = (inp[13]) ? 4'b1000 : node4108;
														assign node4108 = (inp[12]) ? node4110 : 4'b1100;
															assign node4110 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node4114 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4117 = (inp[12]) ? node4123 : node4118;
													assign node4118 = (inp[2]) ? 4'b0000 : node4119;
														assign node4119 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4123 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node4126 = (inp[2]) ? node4138 : node4127;
												assign node4127 = (inp[13]) ? node4133 : node4128;
													assign node4128 = (inp[10]) ? 4'b0001 : node4129;
														assign node4129 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node4133 = (inp[14]) ? 4'b0101 : node4134;
														assign node4134 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node4138 = (inp[10]) ? node4144 : node4139;
													assign node4139 = (inp[13]) ? node4141 : 4'b1000;
														assign node4141 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node4144 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node4147 = (inp[2]) ? node4173 : node4148;
											assign node4148 = (inp[4]) ? node4158 : node4149;
												assign node4149 = (inp[10]) ? node4153 : node4150;
													assign node4150 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node4153 = (inp[1]) ? 4'b0000 : node4154;
														assign node4154 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node4158 = (inp[10]) ? node4170 : node4159;
													assign node4159 = (inp[1]) ? node4161 : 4'b1000;
														assign node4161 = (inp[14]) ? 4'b0001 : node4162;
															assign node4162 = (inp[12]) ? node4166 : node4163;
																assign node4163 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node4166 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node4170 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node4173 = (inp[4]) ? node4189 : node4174;
												assign node4174 = (inp[13]) ? node4180 : node4175;
													assign node4175 = (inp[14]) ? 4'b1000 : node4176;
														assign node4176 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node4180 = (inp[14]) ? node4186 : node4181;
														assign node4181 = (inp[10]) ? 4'b0000 : node4182;
															assign node4182 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4186 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node4189 = (inp[13]) ? node4201 : node4190;
													assign node4190 = (inp[10]) ? node4196 : node4191;
														assign node4191 = (inp[1]) ? 4'b1000 : node4192;
															assign node4192 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4196 = (inp[14]) ? node4198 : 4'b0000;
															assign node4198 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4201 = (inp[12]) ? node4203 : 4'b0100;
														assign node4203 = (inp[10]) ? 4'b1000 : 4'b0000;
								assign node4206 = (inp[1]) ? node4316 : node4207;
									assign node4207 = (inp[3]) ? node4263 : node4208;
										assign node4208 = (inp[2]) ? node4230 : node4209;
											assign node4209 = (inp[4]) ? node4219 : node4210;
												assign node4210 = (inp[12]) ? node4214 : node4211;
													assign node4211 = (inp[10]) ? 4'b0001 : 4'b1100;
													assign node4214 = (inp[10]) ? 4'b1100 : node4215;
														assign node4215 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node4219 = (inp[13]) ? node4225 : node4220;
													assign node4220 = (inp[14]) ? node4222 : 4'b1001;
														assign node4222 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node4225 = (inp[12]) ? 4'b1101 : node4226;
														assign node4226 = (inp[10]) ? 4'b0101 : 4'b1101;
											assign node4230 = (inp[4]) ? node4244 : node4231;
												assign node4231 = (inp[13]) ? node4237 : node4232;
													assign node4232 = (inp[7]) ? 4'b1100 : node4233;
														assign node4233 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node4237 = (inp[10]) ? node4241 : node4238;
														assign node4238 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node4241 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node4244 = (inp[7]) ? node4254 : node4245;
													assign node4245 = (inp[10]) ? node4251 : node4246;
														assign node4246 = (inp[12]) ? node4248 : 4'b1000;
															assign node4248 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node4251 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node4254 = (inp[13]) ? node4258 : node4255;
														assign node4255 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node4258 = (inp[12]) ? node4260 : 4'b0000;
															assign node4260 = (inp[10]) ? 4'b0000 : 4'b1100;
										assign node4263 = (inp[10]) ? node4291 : node4264;
											assign node4264 = (inp[12]) ? node4278 : node4265;
												assign node4265 = (inp[13]) ? node4271 : node4266;
													assign node4266 = (inp[7]) ? node4268 : 4'b1000;
														assign node4268 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node4271 = (inp[4]) ? node4275 : node4272;
														assign node4272 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node4275 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node4278 = (inp[7]) ? node4288 : node4279;
													assign node4279 = (inp[2]) ? node4283 : node4280;
														assign node4280 = (inp[4]) ? 4'b1000 : 4'b0001;
														assign node4283 = (inp[13]) ? node4285 : 4'b0001;
															assign node4285 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4288 = (inp[13]) ? 4'b1000 : 4'b0101;
											assign node4291 = (inp[12]) ? node4305 : node4292;
												assign node4292 = (inp[13]) ? node4300 : node4293;
													assign node4293 = (inp[7]) ? node4297 : node4294;
														assign node4294 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node4297 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node4300 = (inp[2]) ? 4'b0001 : node4301;
														assign node4301 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node4305 = (inp[2]) ? node4311 : node4306;
													assign node4306 = (inp[4]) ? 4'b0000 : node4307;
														assign node4307 = (inp[14]) ? 4'b1001 : 4'b1101;
													assign node4311 = (inp[4]) ? 4'b1001 : node4312;
														assign node4312 = (inp[14]) ? 4'b0000 : 4'b1000;
									assign node4316 = (inp[10]) ? node4364 : node4317;
										assign node4317 = (inp[3]) ? node4335 : node4318;
											assign node4318 = (inp[2]) ? node4328 : node4319;
												assign node4319 = (inp[4]) ? node4325 : node4320;
													assign node4320 = (inp[12]) ? 4'b1001 : node4321;
														assign node4321 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node4325 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node4328 = (inp[12]) ? node4332 : node4329;
													assign node4329 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node4332 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node4335 = (inp[7]) ? node4347 : node4336;
												assign node4336 = (inp[4]) ? node4342 : node4337;
													assign node4337 = (inp[12]) ? 4'b1001 : node4338;
														assign node4338 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node4342 = (inp[13]) ? 4'b1101 : node4343;
														assign node4343 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node4347 = (inp[14]) ? node4359 : node4348;
													assign node4348 = (inp[13]) ? node4350 : 4'b1001;
														assign node4350 = (inp[4]) ? node4354 : node4351;
															assign node4351 = (inp[2]) ? 4'b0001 : 4'b1101;
															assign node4354 = (inp[12]) ? node4356 : 4'b1001;
																assign node4356 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node4359 = (inp[13]) ? 4'b0001 : node4360;
														assign node4360 = (inp[4]) ? 4'b0001 : 4'b1001;
										assign node4364 = (inp[13]) ? node4400 : node4365;
											assign node4365 = (inp[14]) ? node4379 : node4366;
												assign node4366 = (inp[2]) ? node4372 : node4367;
													assign node4367 = (inp[3]) ? node4369 : 4'b0001;
														assign node4369 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node4372 = (inp[3]) ? node4376 : node4373;
														assign node4373 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node4376 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4379 = (inp[4]) ? node4385 : node4380;
													assign node4380 = (inp[3]) ? node4382 : 4'b1101;
														assign node4382 = (inp[2]) ? 4'b1001 : 4'b0101;
													assign node4385 = (inp[12]) ? node4395 : node4386;
														assign node4386 = (inp[7]) ? node4392 : node4387;
															assign node4387 = (inp[2]) ? node4389 : 4'b0101;
																assign node4389 = (inp[3]) ? 4'b0101 : 4'b1001;
															assign node4392 = (inp[3]) ? 4'b1001 : 4'b1101;
														assign node4395 = (inp[3]) ? 4'b1001 : node4396;
															assign node4396 = (inp[2]) ? 4'b1001 : 4'b0001;
											assign node4400 = (inp[4]) ? node4408 : node4401;
												assign node4401 = (inp[14]) ? 4'b0001 : node4402;
													assign node4402 = (inp[2]) ? node4404 : 4'b0001;
														assign node4404 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node4408 = (inp[2]) ? node4410 : 4'b0101;
													assign node4410 = (inp[3]) ? 4'b0101 : 4'b0001;
							assign node4413 = (inp[2]) ? 4'b0101 : node4414;
								assign node4414 = (inp[3]) ? node4466 : node4415;
									assign node4415 = (inp[4]) ? node4431 : node4416;
										assign node4416 = (inp[12]) ? 4'b0101 : node4417;
											assign node4417 = (inp[7]) ? 4'b0101 : node4418;
												assign node4418 = (inp[13]) ? node4420 : 4'b0101;
													assign node4420 = (inp[14]) ? node4424 : node4421;
														assign node4421 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node4424 = (inp[1]) ? 4'b0001 : node4425;
															assign node4425 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node4431 = (inp[7]) ? node4449 : node4432;
											assign node4432 = (inp[1]) ? node4444 : node4433;
												assign node4433 = (inp[14]) ? 4'b0000 : node4434;
													assign node4434 = (inp[10]) ? node4440 : node4435;
														assign node4435 = (inp[13]) ? node4437 : 4'b0000;
															assign node4437 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4440 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node4444 = (inp[13]) ? 4'b0001 : node4445;
													assign node4445 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node4449 = (inp[13]) ? node4451 : 4'b0101;
												assign node4451 = (inp[10]) ? node4459 : node4452;
													assign node4452 = (inp[14]) ? 4'b0101 : node4453;
														assign node4453 = (inp[1]) ? node4455 : 4'b0000;
															assign node4455 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node4459 = (inp[14]) ? node4461 : 4'b0000;
														assign node4461 = (inp[1]) ? 4'b0000 : node4462;
															assign node4462 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node4466 = (inp[7]) ? node4514 : node4467;
										assign node4467 = (inp[4]) ? node4481 : node4468;
											assign node4468 = (inp[1]) ? node4474 : node4469;
												assign node4469 = (inp[13]) ? 4'b0100 : node4470;
													assign node4470 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4474 = (inp[12]) ? node4476 : 4'b1001;
													assign node4476 = (inp[10]) ? 4'b0101 : node4477;
														assign node4477 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node4481 = (inp[11]) ? node4499 : node4482;
												assign node4482 = (inp[14]) ? node4488 : node4483;
													assign node4483 = (inp[1]) ? node4485 : 4'b0100;
														assign node4485 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node4488 = (inp[1]) ? node4492 : node4489;
														assign node4489 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node4492 = (inp[10]) ? 4'b0100 : node4493;
															assign node4493 = (inp[12]) ? node4495 : 4'b0100;
																assign node4495 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node4499 = (inp[1]) ? node4505 : node4500;
													assign node4500 = (inp[14]) ? 4'b1100 : node4501;
														assign node4501 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node4505 = (inp[13]) ? node4509 : node4506;
														assign node4506 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4509 = (inp[12]) ? node4511 : 4'b0101;
															assign node4511 = (inp[10]) ? 4'b0101 : 4'b1101;
										assign node4514 = (inp[1]) ? node4538 : node4515;
											assign node4515 = (inp[14]) ? node4525 : node4516;
												assign node4516 = (inp[13]) ? node4522 : node4517;
													assign node4517 = (inp[12]) ? node4519 : 4'b1000;
														assign node4519 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node4522 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node4525 = (inp[11]) ? node4531 : node4526;
													assign node4526 = (inp[12]) ? node4528 : 4'b1001;
														assign node4528 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node4531 = (inp[10]) ? 4'b1000 : node4532;
														assign node4532 = (inp[12]) ? node4534 : 4'b0100;
															assign node4534 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node4538 = (inp[13]) ? node4544 : node4539;
												assign node4539 = (inp[14]) ? node4541 : 4'b1001;
													assign node4541 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4544 = (inp[12]) ? node4552 : node4545;
													assign node4545 = (inp[4]) ? node4549 : node4546;
														assign node4546 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node4549 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4552 = (inp[10]) ? 4'b0101 : node4553;
														assign node4553 = (inp[11]) ? 4'b1001 : node4554;
															assign node4554 = (inp[14]) ? 4'b1000 : 4'b1001;
						assign node4560 = (inp[3]) ? node4936 : node4561;
							assign node4561 = (inp[4]) ? node4725 : node4562;
								assign node4562 = (inp[7]) ? node4642 : node4563;
									assign node4563 = (inp[2]) ? node4601 : node4564;
										assign node4564 = (inp[0]) ? node4586 : node4565;
											assign node4565 = (inp[1]) ? node4573 : node4566;
												assign node4566 = (inp[14]) ? 4'b1001 : node4567;
													assign node4567 = (inp[13]) ? node4569 : 4'b1100;
														assign node4569 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node4573 = (inp[11]) ? node4581 : node4574;
													assign node4574 = (inp[12]) ? node4576 : 4'b0001;
														assign node4576 = (inp[13]) ? node4578 : 4'b1001;
															assign node4578 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node4581 = (inp[13]) ? node4583 : 4'b0001;
														assign node4583 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node4586 = (inp[11]) ? node4594 : node4587;
												assign node4587 = (inp[10]) ? 4'b0000 : node4588;
													assign node4588 = (inp[13]) ? 4'b0000 : node4589;
														assign node4589 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node4594 = (inp[10]) ? node4596 : 4'b1001;
													assign node4596 = (inp[12]) ? node4598 : 4'b0001;
														assign node4598 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node4601 = (inp[0]) ? node4629 : node4602;
											assign node4602 = (inp[1]) ? node4616 : node4603;
												assign node4603 = (inp[12]) ? node4609 : node4604;
													assign node4604 = (inp[13]) ? node4606 : 4'b0000;
														assign node4606 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node4609 = (inp[13]) ? node4613 : node4610;
														assign node4610 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node4613 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node4616 = (inp[11]) ? node4626 : node4617;
													assign node4617 = (inp[14]) ? node4621 : node4618;
														assign node4618 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node4621 = (inp[10]) ? node4623 : 4'b1100;
															assign node4623 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node4626 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node4629 = (inp[13]) ? node4631 : 4'b0101;
												assign node4631 = (inp[10]) ? node4639 : node4632;
													assign node4632 = (inp[1]) ? node4634 : 4'b0101;
														assign node4634 = (inp[14]) ? node4636 : 4'b0101;
															assign node4636 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node4639 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node4642 = (inp[13]) ? node4684 : node4643;
										assign node4643 = (inp[2]) ? node4667 : node4644;
											assign node4644 = (inp[12]) ? node4654 : node4645;
												assign node4645 = (inp[11]) ? node4651 : node4646;
													assign node4646 = (inp[10]) ? 4'b1100 : node4647;
														assign node4647 = (inp[0]) ? 4'b0101 : 4'b1100;
													assign node4651 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node4654 = (inp[1]) ? node4662 : node4655;
													assign node4655 = (inp[0]) ? 4'b1100 : node4656;
														assign node4656 = (inp[10]) ? 4'b0100 : node4657;
															assign node4657 = (inp[11]) ? 4'b1100 : 4'b0101;
													assign node4662 = (inp[14]) ? 4'b0101 : node4663;
														assign node4663 = (inp[10]) ? 4'b1100 : 4'b0101;
											assign node4667 = (inp[11]) ? node4673 : node4668;
												assign node4668 = (inp[0]) ? 4'b0101 : node4669;
													assign node4669 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node4673 = (inp[0]) ? 4'b0101 : node4674;
													assign node4674 = (inp[12]) ? node4676 : 4'b0101;
														assign node4676 = (inp[1]) ? node4680 : node4677;
															assign node4677 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node4680 = (inp[10]) ? 4'b0101 : 4'b1101;
										assign node4684 = (inp[0]) ? node4702 : node4685;
											assign node4685 = (inp[2]) ? node4697 : node4686;
												assign node4686 = (inp[1]) ? node4692 : node4687;
													assign node4687 = (inp[11]) ? 4'b1001 : node4688;
														assign node4688 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4692 = (inp[12]) ? 4'b1001 : node4693;
														assign node4693 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node4697 = (inp[1]) ? 4'b0001 : node4698;
													assign node4698 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node4702 = (inp[2]) ? 4'b0101 : node4703;
												assign node4703 = (inp[12]) ? node4711 : node4704;
													assign node4704 = (inp[10]) ? node4708 : node4705;
														assign node4705 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node4708 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node4711 = (inp[10]) ? node4717 : node4712;
														assign node4712 = (inp[1]) ? 4'b1101 : node4713;
															assign node4713 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node4717 = (inp[1]) ? 4'b0001 : node4718;
															assign node4718 = (inp[14]) ? node4720 : 4'b0100;
																assign node4720 = (inp[11]) ? 4'b0100 : 4'b1101;
								assign node4725 = (inp[11]) ? node4863 : node4726;
									assign node4726 = (inp[2]) ? node4794 : node4727;
										assign node4727 = (inp[1]) ? node4763 : node4728;
											assign node4728 = (inp[13]) ? node4740 : node4729;
												assign node4729 = (inp[0]) ? node4733 : node4730;
													assign node4730 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node4733 = (inp[7]) ? 4'b1000 : node4734;
														assign node4734 = (inp[12]) ? node4736 : 4'b1000;
															assign node4736 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node4740 = (inp[12]) ? node4752 : node4741;
													assign node4741 = (inp[7]) ? node4747 : node4742;
														assign node4742 = (inp[10]) ? 4'b1001 : node4743;
															assign node4743 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4747 = (inp[14]) ? node4749 : 4'b0000;
															assign node4749 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node4752 = (inp[10]) ? node4760 : node4753;
														assign node4753 = (inp[0]) ? 4'b0100 : node4754;
															assign node4754 = (inp[14]) ? node4756 : 4'b0100;
																assign node4756 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node4760 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node4763 = (inp[10]) ? node4779 : node4764;
												assign node4764 = (inp[12]) ? node4770 : node4765;
													assign node4765 = (inp[13]) ? node4767 : 4'b0001;
														assign node4767 = (inp[0]) ? 4'b0001 : 4'b1000;
													assign node4770 = (inp[7]) ? 4'b0000 : node4771;
														assign node4771 = (inp[13]) ? 4'b0001 : node4772;
															assign node4772 = (inp[0]) ? 4'b1000 : node4773;
																assign node4773 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4779 = (inp[13]) ? node4787 : node4780;
													assign node4780 = (inp[7]) ? 4'b0000 : node4781;
														assign node4781 = (inp[12]) ? 4'b0100 : node4782;
															assign node4782 = (inp[0]) ? 4'b0100 : 4'b0000;
													assign node4787 = (inp[7]) ? node4791 : node4788;
														assign node4788 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4791 = (inp[14]) ? 4'b0100 : 4'b1000;
										assign node4794 = (inp[7]) ? node4836 : node4795;
											assign node4795 = (inp[0]) ? node4821 : node4796;
												assign node4796 = (inp[10]) ? node4812 : node4797;
													assign node4797 = (inp[14]) ? node4809 : node4798;
														assign node4798 = (inp[12]) ? node4806 : node4799;
															assign node4799 = (inp[1]) ? node4803 : node4800;
																assign node4800 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node4803 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4806 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node4809 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node4812 = (inp[1]) ? node4816 : node4813;
														assign node4813 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4816 = (inp[12]) ? node4818 : 4'b0001;
															assign node4818 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node4821 = (inp[1]) ? node4829 : node4822;
													assign node4822 = (inp[14]) ? node4824 : 4'b1000;
														assign node4824 = (inp[10]) ? node4826 : 4'b1001;
															assign node4826 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node4829 = (inp[14]) ? node4831 : 4'b0001;
														assign node4831 = (inp[13]) ? 4'b0000 : node4832;
															assign node4832 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node4836 = (inp[0]) ? node4856 : node4837;
												assign node4837 = (inp[10]) ? node4849 : node4838;
													assign node4838 = (inp[14]) ? node4844 : node4839;
														assign node4839 = (inp[13]) ? 4'b0001 : node4840;
															assign node4840 = (inp[1]) ? 4'b1000 : 4'b0001;
														assign node4844 = (inp[13]) ? node4846 : 4'b1001;
															assign node4846 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node4849 = (inp[12]) ? 4'b0101 : node4850;
														assign node4850 = (inp[1]) ? node4852 : 4'b0100;
															assign node4852 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node4856 = (inp[13]) ? node4858 : 4'b0101;
													assign node4858 = (inp[12]) ? node4860 : 4'b0000;
														assign node4860 = (inp[14]) ? 4'b0101 : 4'b0001;
									assign node4863 = (inp[1]) ? node4909 : node4864;
										assign node4864 = (inp[2]) ? node4892 : node4865;
											assign node4865 = (inp[0]) ? node4881 : node4866;
												assign node4866 = (inp[13]) ? node4872 : node4867;
													assign node4867 = (inp[12]) ? node4869 : 4'b0000;
														assign node4869 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node4872 = (inp[12]) ? node4876 : node4873;
														assign node4873 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node4876 = (inp[7]) ? 4'b0100 : node4877;
															assign node4877 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node4881 = (inp[7]) ? node4885 : node4882;
													assign node4882 = (inp[14]) ? 4'b0101 : 4'b1001;
													assign node4885 = (inp[12]) ? node4889 : node4886;
														assign node4886 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node4889 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node4892 = (inp[7]) ? node4900 : node4893;
												assign node4893 = (inp[0]) ? node4897 : node4894;
													assign node4894 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node4897 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node4900 = (inp[0]) ? node4904 : node4901;
													assign node4901 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node4904 = (inp[13]) ? node4906 : 4'b0101;
														assign node4906 = (inp[10]) ? 4'b0000 : 4'b0101;
										assign node4909 = (inp[10]) ? node4923 : node4910;
											assign node4910 = (inp[2]) ? node4912 : 4'b1001;
												assign node4912 = (inp[14]) ? node4918 : node4913;
													assign node4913 = (inp[0]) ? 4'b0101 : node4914;
														assign node4914 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4918 = (inp[7]) ? 4'b0001 : node4919;
														assign node4919 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node4923 = (inp[13]) ? 4'b0001 : node4924;
												assign node4924 = (inp[0]) ? node4926 : 4'b0001;
													assign node4926 = (inp[14]) ? node4932 : node4927;
														assign node4927 = (inp[2]) ? 4'b0101 : node4928;
															assign node4928 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4932 = (inp[2]) ? 4'b1001 : 4'b0101;
							assign node4936 = (inp[13]) ? node5132 : node4937;
								assign node4937 = (inp[1]) ? node5033 : node4938;
									assign node4938 = (inp[0]) ? node4980 : node4939;
										assign node4939 = (inp[10]) ? node4967 : node4940;
											assign node4940 = (inp[7]) ? node4952 : node4941;
												assign node4941 = (inp[2]) ? node4947 : node4942;
													assign node4942 = (inp[11]) ? node4944 : 4'b0001;
														assign node4944 = (inp[4]) ? 4'b1000 : 4'b0001;
													assign node4947 = (inp[4]) ? node4949 : 4'b1001;
														assign node4949 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node4952 = (inp[12]) ? node4960 : node4953;
													assign node4953 = (inp[4]) ? 4'b0001 : node4954;
														assign node4954 = (inp[14]) ? 4'b1000 : node4955;
															assign node4955 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node4960 = (inp[14]) ? node4964 : node4961;
														assign node4961 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node4964 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node4967 = (inp[4]) ? 4'b0001 : node4968;
												assign node4968 = (inp[2]) ? node4976 : node4969;
													assign node4969 = (inp[14]) ? 4'b0001 : node4970;
														assign node4970 = (inp[12]) ? node4972 : 4'b1000;
															assign node4972 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node4976 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node4980 = (inp[10]) ? node5010 : node4981;
											assign node4981 = (inp[12]) ? node4999 : node4982;
												assign node4982 = (inp[4]) ? node4990 : node4983;
													assign node4983 = (inp[11]) ? 4'b1000 : node4984;
														assign node4984 = (inp[14]) ? 4'b0001 : node4985;
															assign node4985 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node4990 = (inp[2]) ? node4994 : node4991;
														assign node4991 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node4994 = (inp[11]) ? node4996 : 4'b1000;
															assign node4996 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node4999 = (inp[4]) ? node5001 : 4'b1000;
													assign node5001 = (inp[14]) ? node5005 : node5002;
														assign node5002 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node5005 = (inp[2]) ? node5007 : 4'b1000;
															assign node5007 = (inp[11]) ? 4'b1000 : 4'b0000;
											assign node5010 = (inp[11]) ? node5026 : node5011;
												assign node5011 = (inp[12]) ? node5015 : node5012;
													assign node5012 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node5015 = (inp[14]) ? node5017 : 4'b0001;
														assign node5017 = (inp[4]) ? node5019 : 4'b0000;
															assign node5019 = (inp[2]) ? node5023 : node5020;
																assign node5020 = (inp[7]) ? 4'b1001 : 4'b0000;
																assign node5023 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node5026 = (inp[7]) ? 4'b1000 : node5027;
													assign node5027 = (inp[4]) ? node5029 : 4'b0001;
														assign node5029 = (inp[2]) ? 4'b0000 : 4'b1000;
									assign node5033 = (inp[11]) ? node5085 : node5034;
										assign node5034 = (inp[10]) ? node5064 : node5035;
											assign node5035 = (inp[2]) ? node5051 : node5036;
												assign node5036 = (inp[12]) ? node5048 : node5037;
													assign node5037 = (inp[14]) ? node5045 : node5038;
														assign node5038 = (inp[7]) ? node5040 : 4'b0000;
															assign node5040 = (inp[0]) ? node5042 : 4'b1001;
																assign node5042 = (inp[4]) ? 4'b1000 : 4'b0000;
														assign node5045 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node5048 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node5051 = (inp[4]) ? node5057 : node5052;
													assign node5052 = (inp[7]) ? 4'b0001 : node5053;
														assign node5053 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5057 = (inp[12]) ? node5061 : node5058;
														assign node5058 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node5061 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node5064 = (inp[12]) ? node5078 : node5065;
												assign node5065 = (inp[2]) ? node5073 : node5066;
													assign node5066 = (inp[4]) ? 4'b0000 : node5067;
														assign node5067 = (inp[14]) ? node5069 : 4'b0001;
															assign node5069 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node5073 = (inp[7]) ? 4'b0000 : node5074;
														assign node5074 = (inp[0]) ? 4'b0000 : 4'b1000;
												assign node5078 = (inp[4]) ? node5080 : 4'b1001;
													assign node5080 = (inp[7]) ? 4'b0001 : node5081;
														assign node5081 = (inp[0]) ? 4'b0001 : 4'b1000;
										assign node5085 = (inp[4]) ? node5111 : node5086;
											assign node5086 = (inp[2]) ? node5100 : node5087;
												assign node5087 = (inp[7]) ? node5089 : 4'b0001;
													assign node5089 = (inp[14]) ? node5093 : node5090;
														assign node5090 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node5093 = (inp[0]) ? node5095 : 4'b0001;
															assign node5095 = (inp[10]) ? 4'b0001 : node5096;
																assign node5096 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node5100 = (inp[12]) ? node5108 : node5101;
													assign node5101 = (inp[0]) ? 4'b1001 : node5102;
														assign node5102 = (inp[7]) ? node5104 : 4'b1001;
															assign node5104 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node5108 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node5111 = (inp[10]) ? 4'b0001 : node5112;
												assign node5112 = (inp[0]) ? node5118 : node5113;
													assign node5113 = (inp[2]) ? node5115 : 4'b0001;
														assign node5115 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node5118 = (inp[14]) ? node5126 : node5119;
														assign node5119 = (inp[7]) ? 4'b0001 : node5120;
															assign node5120 = (inp[12]) ? 4'b0001 : node5121;
																assign node5121 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node5126 = (inp[7]) ? node5128 : 4'b0001;
															assign node5128 = (inp[2]) ? 4'b1001 : 4'b0001;
								assign node5132 = (inp[4]) ? node5222 : node5133;
									assign node5133 = (inp[11]) ? node5179 : node5134;
										assign node5134 = (inp[0]) ? node5154 : node5135;
											assign node5135 = (inp[10]) ? node5143 : node5136;
												assign node5136 = (inp[12]) ? node5138 : 4'b0000;
													assign node5138 = (inp[14]) ? node5140 : 4'b0000;
														assign node5140 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node5143 = (inp[14]) ? node5151 : node5144;
													assign node5144 = (inp[1]) ? 4'b1001 : node5145;
														assign node5145 = (inp[12]) ? 4'b1001 : node5146;
															assign node5146 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node5151 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node5154 = (inp[2]) ? node5170 : node5155;
												assign node5155 = (inp[10]) ? node5165 : node5156;
													assign node5156 = (inp[14]) ? 4'b0001 : node5157;
														assign node5157 = (inp[1]) ? node5161 : node5158;
															assign node5158 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node5161 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node5165 = (inp[1]) ? node5167 : 4'b0000;
														assign node5167 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node5170 = (inp[12]) ? node5172 : 4'b0000;
													assign node5172 = (inp[7]) ? 4'b1000 : node5173;
														assign node5173 = (inp[10]) ? node5175 : 4'b0000;
															assign node5175 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node5179 = (inp[1]) ? node5209 : node5180;
											assign node5180 = (inp[0]) ? node5194 : node5181;
												assign node5181 = (inp[7]) ? node5189 : node5182;
													assign node5182 = (inp[12]) ? node5184 : 4'b0001;
														assign node5184 = (inp[10]) ? 4'b0000 : node5185;
															assign node5185 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node5189 = (inp[2]) ? node5191 : 4'b1001;
														assign node5191 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node5194 = (inp[12]) ? node5204 : node5195;
													assign node5195 = (inp[2]) ? node5201 : node5196;
														assign node5196 = (inp[10]) ? node5198 : 4'b1000;
															assign node5198 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node5201 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node5204 = (inp[2]) ? 4'b1001 : node5205;
														assign node5205 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node5209 = (inp[12]) ? 4'b0001 : node5210;
												assign node5210 = (inp[10]) ? 4'b0001 : node5211;
													assign node5211 = (inp[7]) ? node5215 : node5212;
														assign node5212 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node5215 = (inp[14]) ? 4'b0001 : node5216;
															assign node5216 = (inp[0]) ? 4'b0001 : 4'b1001;
									assign node5222 = (inp[10]) ? node5256 : node5223;
										assign node5223 = (inp[11]) ? node5245 : node5224;
											assign node5224 = (inp[0]) ? node5234 : node5225;
												assign node5225 = (inp[7]) ? 4'b0001 : node5226;
													assign node5226 = (inp[2]) ? node5228 : 4'b0000;
														assign node5228 = (inp[14]) ? 4'b0001 : node5229;
															assign node5229 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node5234 = (inp[12]) ? node5242 : node5235;
													assign node5235 = (inp[14]) ? 4'b0001 : node5236;
														assign node5236 = (inp[1]) ? node5238 : 4'b0000;
															assign node5238 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node5242 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node5245 = (inp[1]) ? 4'b0001 : node5246;
												assign node5246 = (inp[0]) ? node5248 : 4'b0001;
													assign node5248 = (inp[12]) ? node5252 : node5249;
														assign node5249 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node5252 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node5256 = (inp[11]) ? 4'b0000 : node5257;
											assign node5257 = (inp[1]) ? 4'b0000 : node5258;
												assign node5258 = (inp[2]) ? node5264 : node5259;
													assign node5259 = (inp[7]) ? node5261 : 4'b0001;
														assign node5261 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node5264 = (inp[12]) ? 4'b0000 : node5265;
														assign node5265 = (inp[0]) ? 4'b0000 : 4'b0001;
				assign node5271 = (inp[0]) ? node6433 : node5272;
					assign node5272 = (inp[6]) ? node5616 : node5273;
						assign node5273 = (inp[2]) ? node5549 : node5274;
							assign node5274 = (inp[5]) ? node5340 : node5275;
								assign node5275 = (inp[3]) ? node5277 : 4'b0011;
									assign node5277 = (inp[7]) ? node5321 : node5278;
										assign node5278 = (inp[4]) ? node5296 : node5279;
											assign node5279 = (inp[13]) ? node5281 : 4'b0011;
												assign node5281 = (inp[12]) ? node5291 : node5282;
													assign node5282 = (inp[14]) ? node5284 : 4'b0001;
														assign node5284 = (inp[10]) ? node5286 : 4'b0000;
															assign node5286 = (inp[11]) ? node5288 : 4'b0001;
																assign node5288 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node5291 = (inp[14]) ? 4'b0011 : node5292;
														assign node5292 = (inp[1]) ? 4'b0011 : 4'b0000;
											assign node5296 = (inp[1]) ? node5312 : node5297;
												assign node5297 = (inp[11]) ? node5307 : node5298;
													assign node5298 = (inp[14]) ? node5302 : node5299;
														assign node5299 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node5302 = (inp[13]) ? node5304 : 4'b0001;
															assign node5304 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5307 = (inp[14]) ? node5309 : 4'b1000;
														assign node5309 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node5312 = (inp[10]) ? node5318 : node5313;
													assign node5313 = (inp[14]) ? node5315 : 4'b1001;
														assign node5315 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node5318 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node5321 = (inp[13]) ? node5323 : 4'b0011;
											assign node5323 = (inp[4]) ? node5325 : 4'b0011;
												assign node5325 = (inp[11]) ? node5337 : node5326;
													assign node5326 = (inp[12]) ? node5332 : node5327;
														assign node5327 = (inp[14]) ? node5329 : 4'b0001;
															assign node5329 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node5332 = (inp[1]) ? node5334 : 4'b0011;
															assign node5334 = (inp[10]) ? 4'b0000 : 4'b0011;
													assign node5337 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node5340 = (inp[1]) ? node5450 : node5341;
									assign node5341 = (inp[14]) ? node5387 : node5342;
										assign node5342 = (inp[13]) ? node5370 : node5343;
											assign node5343 = (inp[12]) ? node5359 : node5344;
												assign node5344 = (inp[11]) ? node5354 : node5345;
													assign node5345 = (inp[3]) ? node5349 : node5346;
														assign node5346 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5349 = (inp[7]) ? 4'b1100 : node5350;
															assign node5350 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node5354 = (inp[7]) ? node5356 : 4'b1000;
														assign node5356 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node5359 = (inp[10]) ? node5363 : node5360;
													assign node5360 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node5363 = (inp[3]) ? node5365 : 4'b1000;
														assign node5365 = (inp[4]) ? node5367 : 4'b1100;
															assign node5367 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node5370 = (inp[10]) ? node5380 : node5371;
												assign node5371 = (inp[12]) ? node5377 : node5372;
													assign node5372 = (inp[3]) ? 4'b0000 : node5373;
														assign node5373 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node5377 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node5380 = (inp[3]) ? 4'b0000 : node5381;
													assign node5381 = (inp[7]) ? node5383 : 4'b0100;
														assign node5383 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node5387 = (inp[11]) ? node5421 : node5388;
											assign node5388 = (inp[13]) ? node5404 : node5389;
												assign node5389 = (inp[10]) ? node5395 : node5390;
													assign node5390 = (inp[3]) ? 4'b0101 : node5391;
														assign node5391 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node5395 = (inp[12]) ? node5397 : 4'b1001;
														assign node5397 = (inp[4]) ? node5399 : 4'b0001;
															assign node5399 = (inp[7]) ? 4'b0101 : node5400;
																assign node5400 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node5404 = (inp[10]) ? node5412 : node5405;
													assign node5405 = (inp[3]) ? node5407 : 4'b1001;
														assign node5407 = (inp[4]) ? node5409 : 4'b1101;
															assign node5409 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node5412 = (inp[12]) ? node5418 : node5413;
														assign node5413 = (inp[3]) ? 4'b0001 : node5414;
															assign node5414 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node5418 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node5421 = (inp[13]) ? node5431 : node5422;
												assign node5422 = (inp[10]) ? node5426 : node5423;
													assign node5423 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node5426 = (inp[3]) ? 4'b1100 : node5427;
														assign node5427 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node5431 = (inp[12]) ? node5439 : node5432;
													assign node5432 = (inp[10]) ? 4'b0100 : node5433;
														assign node5433 = (inp[3]) ? node5435 : 4'b0000;
															assign node5435 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node5439 = (inp[10]) ? 4'b0100 : node5440;
														assign node5440 = (inp[4]) ? node5444 : node5441;
															assign node5441 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node5444 = (inp[3]) ? node5446 : 4'b1100;
																assign node5446 = (inp[7]) ? 4'b1100 : 4'b1000;
									assign node5450 = (inp[11]) ? node5510 : node5451;
										assign node5451 = (inp[14]) ? node5469 : node5452;
											assign node5452 = (inp[3]) ? node5458 : node5453;
												assign node5453 = (inp[7]) ? 4'b1001 : node5454;
													assign node5454 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node5458 = (inp[13]) ? node5466 : node5459;
													assign node5459 = (inp[12]) ? node5463 : node5460;
														assign node5460 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node5463 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node5466 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node5469 = (inp[13]) ? node5493 : node5470;
												assign node5470 = (inp[10]) ? node5482 : node5471;
													assign node5471 = (inp[12]) ? node5473 : 4'b1100;
														assign node5473 = (inp[3]) ? node5477 : node5474;
															assign node5474 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node5477 = (inp[4]) ? node5479 : 4'b0100;
																assign node5479 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node5482 = (inp[7]) ? 4'b1100 : node5483;
														assign node5483 = (inp[12]) ? node5487 : node5484;
															assign node5484 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node5487 = (inp[3]) ? node5489 : 4'b1000;
																assign node5489 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node5493 = (inp[12]) ? node5501 : node5494;
													assign node5494 = (inp[7]) ? node5496 : 4'b0100;
														assign node5496 = (inp[4]) ? 4'b0000 : node5497;
															assign node5497 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node5501 = (inp[10]) ? 4'b0000 : node5502;
														assign node5502 = (inp[4]) ? node5504 : 4'b1000;
															assign node5504 = (inp[3]) ? 4'b1000 : node5505;
																assign node5505 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node5510 = (inp[13]) ? node5534 : node5511;
											assign node5511 = (inp[10]) ? node5525 : node5512;
												assign node5512 = (inp[12]) ? node5520 : node5513;
													assign node5513 = (inp[7]) ? 4'b1101 : node5514;
														assign node5514 = (inp[14]) ? node5516 : 4'b1001;
															assign node5516 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node5520 = (inp[7]) ? node5522 : 4'b0101;
														assign node5522 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node5525 = (inp[4]) ? node5529 : node5526;
													assign node5526 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node5529 = (inp[7]) ? 4'b1001 : node5530;
														assign node5530 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node5534 = (inp[4]) ? node5544 : node5535;
												assign node5535 = (inp[10]) ? 4'b0101 : node5536;
													assign node5536 = (inp[12]) ? node5540 : node5537;
														assign node5537 = (inp[14]) ? 4'b0001 : 4'b0101;
														assign node5540 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node5544 = (inp[12]) ? node5546 : 4'b0001;
													assign node5546 = (inp[10]) ? 4'b0001 : 4'b1001;
							assign node5549 = (inp[5]) ? node5551 : 4'b0011;
								assign node5551 = (inp[3]) ? node5553 : 4'b0011;
									assign node5553 = (inp[7]) ? node5599 : node5554;
										assign node5554 = (inp[4]) ? node5568 : node5555;
											assign node5555 = (inp[13]) ? node5557 : 4'b0011;
												assign node5557 = (inp[14]) ? node5561 : node5558;
													assign node5558 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node5561 = (inp[11]) ? node5565 : node5562;
														assign node5562 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node5565 = (inp[1]) ? 4'b0011 : 4'b0000;
											assign node5568 = (inp[13]) ? node5580 : node5569;
												assign node5569 = (inp[1]) ? node5575 : node5570;
													assign node5570 = (inp[10]) ? 4'b1000 : node5571;
														assign node5571 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node5575 = (inp[10]) ? 4'b1001 : node5576;
														assign node5576 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node5580 = (inp[12]) ? node5592 : node5581;
													assign node5581 = (inp[11]) ? 4'b0001 : node5582;
														assign node5582 = (inp[10]) ? node5584 : 4'b0000;
															assign node5584 = (inp[14]) ? node5588 : node5585;
																assign node5585 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node5588 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node5592 = (inp[10]) ? node5596 : node5593;
														assign node5593 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node5596 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node5599 = (inp[13]) ? node5601 : 4'b0011;
											assign node5601 = (inp[4]) ? node5603 : 4'b0011;
												assign node5603 = (inp[1]) ? node5609 : node5604;
													assign node5604 = (inp[10]) ? 4'b0000 : node5605;
														assign node5605 = (inp[12]) ? 4'b0011 : 4'b0000;
													assign node5609 = (inp[14]) ? node5611 : 4'b0001;
														assign node5611 = (inp[12]) ? 4'b0011 : node5612;
															assign node5612 = (inp[11]) ? 4'b0001 : 4'b0000;
						assign node5616 = (inp[5]) ? node6024 : node5617;
							assign node5617 = (inp[11]) ? node5827 : node5618;
								assign node5618 = (inp[3]) ? node5734 : node5619;
									assign node5619 = (inp[7]) ? node5683 : node5620;
										assign node5620 = (inp[2]) ? node5650 : node5621;
											assign node5621 = (inp[1]) ? node5635 : node5622;
												assign node5622 = (inp[13]) ? node5626 : node5623;
													assign node5623 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node5626 = (inp[4]) ? node5630 : node5627;
														assign node5627 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5630 = (inp[12]) ? 4'b0000 : node5631;
															assign node5631 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node5635 = (inp[14]) ? node5641 : node5636;
													assign node5636 = (inp[13]) ? 4'b0101 : node5637;
														assign node5637 = (inp[4]) ? 4'b0000 : 4'b1001;
													assign node5641 = (inp[4]) ? 4'b1100 : node5642;
														assign node5642 = (inp[13]) ? 4'b1000 : node5643;
															assign node5643 = (inp[12]) ? node5645 : 4'b1000;
																assign node5645 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node5650 = (inp[4]) ? node5662 : node5651;
												assign node5651 = (inp[10]) ? node5659 : node5652;
													assign node5652 = (inp[14]) ? node5656 : node5653;
														assign node5653 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node5656 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node5659 = (inp[13]) ? 4'b0100 : 4'b1001;
												assign node5662 = (inp[13]) ? node5672 : node5663;
													assign node5663 = (inp[10]) ? node5667 : node5664;
														assign node5664 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5667 = (inp[1]) ? node5669 : 4'b1100;
															assign node5669 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node5672 = (inp[14]) ? node5676 : node5673;
														assign node5673 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node5676 = (inp[1]) ? node5678 : 4'b1101;
															assign node5678 = (inp[10]) ? 4'b0100 : node5679;
																assign node5679 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node5683 = (inp[13]) ? node5709 : node5684;
											assign node5684 = (inp[12]) ? node5696 : node5685;
												assign node5685 = (inp[2]) ? node5691 : node5686;
													assign node5686 = (inp[1]) ? 4'b1000 : node5687;
														assign node5687 = (inp[10]) ? 4'b1000 : 4'b0001;
													assign node5691 = (inp[10]) ? 4'b1001 : node5692;
														assign node5692 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node5696 = (inp[2]) ? node5704 : node5697;
													assign node5697 = (inp[14]) ? 4'b0001 : node5698;
														assign node5698 = (inp[10]) ? node5700 : 4'b0001;
															assign node5700 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node5704 = (inp[10]) ? node5706 : 4'b0000;
														assign node5706 = (inp[4]) ? 4'b1000 : 4'b0001;
											assign node5709 = (inp[4]) ? node5721 : node5710;
												assign node5710 = (inp[12]) ? node5714 : node5711;
													assign node5711 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5714 = (inp[10]) ? node5716 : 4'b1001;
														assign node5716 = (inp[2]) ? node5718 : 4'b0000;
															assign node5718 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node5721 = (inp[14]) ? node5729 : node5722;
													assign node5722 = (inp[2]) ? 4'b0101 : node5723;
														assign node5723 = (inp[10]) ? node5725 : 4'b0101;
															assign node5725 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node5729 = (inp[10]) ? node5731 : 4'b1000;
														assign node5731 = (inp[12]) ? 4'b0100 : 4'b0000;
									assign node5734 = (inp[2]) ? node5768 : node5735;
										assign node5735 = (inp[10]) ? node5749 : node5736;
											assign node5736 = (inp[1]) ? node5738 : 4'b0000;
												assign node5738 = (inp[4]) ? node5742 : node5739;
													assign node5739 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node5742 = (inp[13]) ? node5744 : 4'b1100;
														assign node5744 = (inp[7]) ? 4'b1100 : node5745;
															assign node5745 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node5749 = (inp[1]) ? node5757 : node5750;
												assign node5750 = (inp[13]) ? 4'b1001 : node5751;
													assign node5751 = (inp[7]) ? 4'b1100 : node5752;
														assign node5752 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node5757 = (inp[7]) ? node5761 : node5758;
													assign node5758 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node5761 = (inp[14]) ? node5763 : 4'b0000;
														assign node5763 = (inp[4]) ? node5765 : 4'b0000;
															assign node5765 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node5768 = (inp[7]) ? node5798 : node5769;
											assign node5769 = (inp[4]) ? node5785 : node5770;
												assign node5770 = (inp[12]) ? node5774 : node5771;
													assign node5771 = (inp[13]) ? 4'b0000 : 4'b1101;
													assign node5774 = (inp[13]) ? 4'b1101 : node5775;
														assign node5775 = (inp[10]) ? node5781 : node5776;
															assign node5776 = (inp[1]) ? node5778 : 4'b0100;
																assign node5778 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node5781 = (inp[14]) ? 4'b0101 : 4'b1100;
												assign node5785 = (inp[1]) ? node5793 : node5786;
													assign node5786 = (inp[14]) ? node5788 : 4'b1000;
														assign node5788 = (inp[10]) ? 4'b0000 : node5789;
															assign node5789 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5793 = (inp[14]) ? 4'b0000 : node5794;
														assign node5794 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node5798 = (inp[4]) ? node5814 : node5799;
												assign node5799 = (inp[10]) ? node5805 : node5800;
													assign node5800 = (inp[14]) ? node5802 : 4'b0101;
														assign node5802 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node5805 = (inp[13]) ? node5809 : node5806;
														assign node5806 = (inp[12]) ? 4'b1101 : 4'b1100;
														assign node5809 = (inp[14]) ? node5811 : 4'b0101;
															assign node5811 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node5814 = (inp[12]) ? node5816 : 4'b1100;
													assign node5816 = (inp[10]) ? node5820 : node5817;
														assign node5817 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node5820 = (inp[13]) ? node5822 : 4'b1101;
															assign node5822 = (inp[14]) ? node5824 : 4'b0000;
																assign node5824 = (inp[1]) ? 4'b0000 : 4'b1101;
								assign node5827 = (inp[1]) ? node5939 : node5828;
									assign node5828 = (inp[3]) ? node5872 : node5829;
										assign node5829 = (inp[4]) ? node5845 : node5830;
											assign node5830 = (inp[13]) ? node5836 : node5831;
												assign node5831 = (inp[12]) ? node5833 : 4'b1000;
													assign node5833 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node5836 = (inp[10]) ? node5842 : node5837;
													assign node5837 = (inp[12]) ? 4'b1000 : node5838;
														assign node5838 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node5842 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node5845 = (inp[2]) ? node5861 : node5846;
												assign node5846 = (inp[13]) ? node5856 : node5847;
													assign node5847 = (inp[7]) ? node5853 : node5848;
														assign node5848 = (inp[10]) ? 4'b0001 : node5849;
															assign node5849 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node5853 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node5856 = (inp[7]) ? node5858 : 4'b1001;
														assign node5858 = (inp[14]) ? 4'b0100 : 4'b0001;
												assign node5861 = (inp[13]) ? node5867 : node5862;
													assign node5862 = (inp[14]) ? 4'b1000 : node5863;
														assign node5863 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node5867 = (inp[14]) ? 4'b0100 : node5868;
														assign node5868 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node5872 = (inp[2]) ? node5914 : node5873;
											assign node5873 = (inp[4]) ? node5897 : node5874;
												assign node5874 = (inp[7]) ? node5886 : node5875;
													assign node5875 = (inp[14]) ? node5883 : node5876;
														assign node5876 = (inp[10]) ? 4'b0101 : node5877;
															assign node5877 = (inp[13]) ? 4'b0101 : node5878;
																assign node5878 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5883 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node5886 = (inp[13]) ? 4'b1001 : node5887;
														assign node5887 = (inp[14]) ? node5891 : node5888;
															assign node5888 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5891 = (inp[10]) ? 4'b1001 : node5892;
																assign node5892 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node5897 = (inp[13]) ? node5903 : node5898;
													assign node5898 = (inp[12]) ? node5900 : 4'b1101;
														assign node5900 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node5903 = (inp[7]) ? node5907 : node5904;
														assign node5904 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5907 = (inp[14]) ? 4'b0000 : node5908;
															assign node5908 = (inp[10]) ? 4'b1101 : node5909;
																assign node5909 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node5914 = (inp[4]) ? node5924 : node5915;
												assign node5915 = (inp[13]) ? node5921 : node5916;
													assign node5916 = (inp[12]) ? node5918 : 4'b1100;
														assign node5918 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node5921 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node5924 = (inp[12]) ? node5928 : node5925;
													assign node5925 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node5928 = (inp[7]) ? node5936 : node5929;
														assign node5929 = (inp[13]) ? node5933 : node5930;
															assign node5930 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node5933 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node5936 = (inp[10]) ? 4'b0000 : 4'b1100;
									assign node5939 = (inp[10]) ? node5989 : node5940;
										assign node5940 = (inp[3]) ? node5966 : node5941;
											assign node5941 = (inp[7]) ? node5957 : node5942;
												assign node5942 = (inp[4]) ? node5950 : node5943;
													assign node5943 = (inp[13]) ? node5947 : node5944;
														assign node5944 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5947 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node5950 = (inp[13]) ? node5952 : 4'b0101;
														assign node5952 = (inp[2]) ? node5954 : 4'b1001;
															assign node5954 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node5957 = (inp[2]) ? node5959 : 4'b0001;
													assign node5959 = (inp[13]) ? node5963 : node5960;
														assign node5960 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5963 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node5966 = (inp[2]) ? node5974 : node5967;
												assign node5967 = (inp[4]) ? node5969 : 4'b1001;
													assign node5969 = (inp[7]) ? 4'b1101 : node5970;
														assign node5970 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node5974 = (inp[7]) ? node5982 : node5975;
													assign node5975 = (inp[14]) ? node5977 : 4'b0001;
														assign node5977 = (inp[4]) ? node5979 : 4'b1101;
															assign node5979 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5982 = (inp[4]) ? node5984 : 4'b0101;
														assign node5984 = (inp[12]) ? node5986 : 4'b1101;
															assign node5986 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node5989 = (inp[13]) ? node5999 : node5990;
											assign node5990 = (inp[3]) ? node5992 : 4'b1001;
												assign node5992 = (inp[12]) ? 4'b0101 : node5993;
													assign node5993 = (inp[7]) ? 4'b0001 : node5994;
														assign node5994 = (inp[4]) ? 4'b0001 : 4'b1101;
											assign node5999 = (inp[14]) ? node6007 : node6000;
												assign node6000 = (inp[7]) ? node6002 : 4'b0001;
													assign node6002 = (inp[2]) ? 4'b0101 : node6003;
														assign node6003 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node6007 = (inp[4]) ? node6019 : node6008;
													assign node6008 = (inp[2]) ? node6010 : 4'b0101;
														assign node6010 = (inp[12]) ? 4'b0001 : node6011;
															assign node6011 = (inp[7]) ? node6015 : node6012;
																assign node6012 = (inp[3]) ? 4'b0001 : 4'b0101;
																assign node6015 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node6019 = (inp[2]) ? node6021 : 4'b0001;
														assign node6021 = (inp[3]) ? 4'b0001 : 4'b0101;
							assign node6024 = (inp[3]) ? node6262 : node6025;
								assign node6025 = (inp[1]) ? node6155 : node6026;
									assign node6026 = (inp[4]) ? node6096 : node6027;
										assign node6027 = (inp[13]) ? node6059 : node6028;
											assign node6028 = (inp[10]) ? node6046 : node6029;
												assign node6029 = (inp[12]) ? node6039 : node6030;
													assign node6030 = (inp[14]) ? node6034 : node6031;
														assign node6031 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node6034 = (inp[11]) ? node6036 : 4'b1000;
															assign node6036 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node6039 = (inp[11]) ? node6043 : node6040;
														assign node6040 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6043 = (inp[2]) ? 4'b0001 : 4'b1000;
												assign node6046 = (inp[7]) ? node6052 : node6047;
													assign node6047 = (inp[12]) ? 4'b1000 : node6048;
														assign node6048 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node6052 = (inp[12]) ? 4'b0000 : node6053;
														assign node6053 = (inp[14]) ? node6055 : 4'b0001;
															assign node6055 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node6059 = (inp[12]) ? node6071 : node6060;
												assign node6060 = (inp[2]) ? node6062 : 4'b0100;
													assign node6062 = (inp[10]) ? node6066 : node6063;
														assign node6063 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node6066 = (inp[14]) ? 4'b0101 : node6067;
															assign node6067 = (inp[11]) ? 4'b0000 : 4'b0100;
												assign node6071 = (inp[10]) ? node6083 : node6072;
													assign node6072 = (inp[14]) ? node6080 : node6073;
														assign node6073 = (inp[7]) ? 4'b0100 : node6074;
															assign node6074 = (inp[2]) ? node6076 : 4'b1101;
																assign node6076 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node6080 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node6083 = (inp[14]) ? node6093 : node6084;
														assign node6084 = (inp[11]) ? node6086 : 4'b1000;
															assign node6086 = (inp[7]) ? node6090 : node6087;
																assign node6087 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node6090 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node6093 = (inp[11]) ? 4'b1001 : 4'b0001;
										assign node6096 = (inp[11]) ? node6130 : node6097;
											assign node6097 = (inp[14]) ? node6117 : node6098;
												assign node6098 = (inp[13]) ? node6112 : node6099;
													assign node6099 = (inp[12]) ? node6105 : node6100;
														assign node6100 = (inp[2]) ? node6102 : 4'b0000;
															assign node6102 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node6105 = (inp[2]) ? node6107 : 4'b0001;
															assign node6107 = (inp[10]) ? 4'b0001 : node6108;
																assign node6108 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node6112 = (inp[2]) ? 4'b1001 : node6113;
														assign node6113 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node6117 = (inp[10]) ? node6125 : node6118;
													assign node6118 = (inp[2]) ? 4'b0100 : node6119;
														assign node6119 = (inp[13]) ? 4'b0101 : node6120;
															assign node6120 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node6125 = (inp[7]) ? node6127 : 4'b0000;
														assign node6127 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node6130 = (inp[2]) ? node6144 : node6131;
												assign node6131 = (inp[13]) ? node6137 : node6132;
													assign node6132 = (inp[10]) ? node6134 : 4'b1001;
														assign node6134 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node6137 = (inp[7]) ? 4'b1000 : node6138;
														assign node6138 = (inp[10]) ? node6140 : 4'b1000;
															assign node6140 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node6144 = (inp[7]) ? 4'b0000 : node6145;
													assign node6145 = (inp[14]) ? node6149 : node6146;
														assign node6146 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node6149 = (inp[13]) ? 4'b0100 : node6150;
															assign node6150 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node6155 = (inp[11]) ? node6217 : node6156;
										assign node6156 = (inp[4]) ? node6180 : node6157;
											assign node6157 = (inp[2]) ? node6171 : node6158;
												assign node6158 = (inp[10]) ? node6164 : node6159;
													assign node6159 = (inp[14]) ? 4'b0101 : node6160;
														assign node6160 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node6164 = (inp[13]) ? node6166 : 4'b0001;
														assign node6166 = (inp[7]) ? 4'b1101 : node6167;
															assign node6167 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node6171 = (inp[10]) ? node6175 : node6172;
													assign node6172 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node6175 = (inp[13]) ? 4'b0100 : node6176;
														assign node6176 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node6180 = (inp[14]) ? node6200 : node6181;
												assign node6181 = (inp[2]) ? node6189 : node6182;
													assign node6182 = (inp[12]) ? 4'b1001 : node6183;
														assign node6183 = (inp[13]) ? 4'b0000 : node6184;
															assign node6184 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node6189 = (inp[10]) ? node6197 : node6190;
														assign node6190 = (inp[7]) ? node6194 : node6191;
															assign node6191 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node6194 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node6197 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node6200 = (inp[10]) ? node6210 : node6201;
													assign node6201 = (inp[13]) ? node6205 : node6202;
														assign node6202 = (inp[2]) ? 4'b1100 : 4'b0101;
														assign node6205 = (inp[12]) ? node6207 : 4'b0001;
															assign node6207 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node6210 = (inp[12]) ? node6212 : 4'b1001;
														assign node6212 = (inp[7]) ? node6214 : 4'b0000;
															assign node6214 = (inp[2]) ? 4'b0001 : 4'b1001;
										assign node6217 = (inp[13]) ? node6243 : node6218;
											assign node6218 = (inp[10]) ? node6232 : node6219;
												assign node6219 = (inp[12]) ? node6227 : node6220;
													assign node6220 = (inp[4]) ? node6222 : 4'b1001;
														assign node6222 = (inp[7]) ? 4'b0001 : node6223;
															assign node6223 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node6227 = (inp[2]) ? node6229 : 4'b0101;
														assign node6229 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node6232 = (inp[4]) ? node6238 : node6233;
													assign node6233 = (inp[7]) ? 4'b1001 : node6234;
														assign node6234 = (inp[2]) ? 4'b0101 : 4'b1101;
													assign node6238 = (inp[7]) ? node6240 : 4'b1001;
														assign node6240 = (inp[2]) ? 4'b1001 : 4'b0101;
											assign node6243 = (inp[10]) ? node6255 : node6244;
												assign node6244 = (inp[12]) ? node6252 : node6245;
													assign node6245 = (inp[14]) ? node6249 : node6246;
														assign node6246 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node6249 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node6252 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node6255 = (inp[4]) ? 4'b0001 : node6256;
													assign node6256 = (inp[2]) ? node6258 : 4'b0001;
														assign node6258 = (inp[7]) ? 4'b0101 : 4'b0001;
								assign node6262 = (inp[4]) ? node6358 : node6263;
									assign node6263 = (inp[11]) ? node6301 : node6264;
										assign node6264 = (inp[13]) ? node6284 : node6265;
											assign node6265 = (inp[12]) ? node6275 : node6266;
												assign node6266 = (inp[1]) ? node6268 : 4'b1001;
													assign node6268 = (inp[2]) ? node6272 : node6269;
														assign node6269 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6272 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node6275 = (inp[10]) ? node6279 : node6276;
													assign node6276 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node6279 = (inp[2]) ? node6281 : 4'b0001;
														assign node6281 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node6284 = (inp[14]) ? node6292 : node6285;
												assign node6285 = (inp[1]) ? node6287 : 4'b1000;
													assign node6287 = (inp[10]) ? node6289 : 4'b0000;
														assign node6289 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node6292 = (inp[12]) ? node6294 : 4'b1000;
													assign node6294 = (inp[10]) ? node6298 : node6295;
														assign node6295 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node6298 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node6301 = (inp[1]) ? node6331 : node6302;
											assign node6302 = (inp[12]) ? node6312 : node6303;
												assign node6303 = (inp[10]) ? node6307 : node6304;
													assign node6304 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node6307 = (inp[7]) ? 4'b0000 : node6308;
														assign node6308 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node6312 = (inp[14]) ? node6322 : node6313;
													assign node6313 = (inp[10]) ? node6315 : 4'b1000;
														assign node6315 = (inp[7]) ? 4'b0000 : node6316;
															assign node6316 = (inp[13]) ? 4'b0001 : node6317;
																assign node6317 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node6322 = (inp[2]) ? 4'b1001 : node6323;
														assign node6323 = (inp[13]) ? 4'b1000 : node6324;
															assign node6324 = (inp[7]) ? 4'b1000 : node6325;
																assign node6325 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node6331 = (inp[10]) ? node6353 : node6332;
												assign node6332 = (inp[13]) ? node6340 : node6333;
													assign node6333 = (inp[7]) ? node6335 : 4'b0001;
														assign node6335 = (inp[12]) ? node6337 : 4'b0001;
															assign node6337 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node6340 = (inp[14]) ? 4'b1001 : node6341;
														assign node6341 = (inp[7]) ? node6347 : node6342;
															assign node6342 = (inp[2]) ? node6344 : 4'b1001;
																assign node6344 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node6347 = (inp[12]) ? 4'b1001 : node6348;
																assign node6348 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node6353 = (inp[7]) ? node6355 : 4'b0001;
													assign node6355 = (inp[2]) ? 4'b1001 : 4'b0001;
									assign node6358 = (inp[10]) ? node6396 : node6359;
										assign node6359 = (inp[13]) ? node6379 : node6360;
											assign node6360 = (inp[14]) ? node6364 : node6361;
												assign node6361 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node6364 = (inp[7]) ? node6374 : node6365;
													assign node6365 = (inp[2]) ? node6367 : 4'b1001;
														assign node6367 = (inp[1]) ? 4'b0001 : node6368;
															assign node6368 = (inp[11]) ? node6370 : 4'b1001;
																assign node6370 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6374 = (inp[12]) ? 4'b1001 : node6375;
														assign node6375 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node6379 = (inp[11]) ? node6387 : node6380;
												assign node6380 = (inp[7]) ? node6384 : node6381;
													assign node6381 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node6384 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node6387 = (inp[1]) ? 4'b0001 : node6388;
													assign node6388 = (inp[2]) ? node6390 : 4'b0000;
														assign node6390 = (inp[14]) ? 4'b0001 : node6391;
															assign node6391 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node6396 = (inp[13]) ? node6426 : node6397;
											assign node6397 = (inp[2]) ? node6413 : node6398;
												assign node6398 = (inp[1]) ? node6408 : node6399;
													assign node6399 = (inp[7]) ? node6401 : 4'b0000;
														assign node6401 = (inp[11]) ? node6405 : node6402;
															assign node6402 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node6405 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6408 = (inp[11]) ? 4'b0001 : node6409;
														assign node6409 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node6413 = (inp[7]) ? node6415 : 4'b0001;
													assign node6415 = (inp[12]) ? node6421 : node6416;
														assign node6416 = (inp[1]) ? 4'b0001 : node6417;
															assign node6417 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node6421 = (inp[11]) ? node6423 : 4'b0000;
															assign node6423 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node6426 = (inp[11]) ? 4'b0000 : node6427;
												assign node6427 = (inp[7]) ? node6429 : 4'b0000;
													assign node6429 = (inp[14]) ? 4'b0001 : 4'b0000;
					assign node6433 = (inp[6]) ? node6435 : 4'b0001;
						assign node6435 = (inp[5]) ? node6489 : node6436;
							assign node6436 = (inp[3]) ? node6438 : 4'b0001;
								assign node6438 = (inp[2]) ? 4'b0001 : node6439;
									assign node6439 = (inp[4]) ? node6447 : node6440;
										assign node6440 = (inp[7]) ? 4'b0001 : node6441;
											assign node6441 = (inp[12]) ? 4'b0001 : node6442;
												assign node6442 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node6447 = (inp[7]) ? node6483 : node6448;
											assign node6448 = (inp[1]) ? node6466 : node6449;
												assign node6449 = (inp[13]) ? node6461 : node6450;
													assign node6450 = (inp[14]) ? node6452 : 4'b1000;
														assign node6452 = (inp[11]) ? node6456 : node6453;
															assign node6453 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node6456 = (inp[12]) ? node6458 : 4'b1000;
																assign node6458 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node6461 = (inp[10]) ? 4'b0000 : node6462;
														assign node6462 = (inp[11]) ? 4'b0000 : 4'b1001;
												assign node6466 = (inp[14]) ? node6476 : node6467;
													assign node6467 = (inp[10]) ? 4'b1001 : node6468;
														assign node6468 = (inp[12]) ? node6472 : node6469;
															assign node6469 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node6472 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node6476 = (inp[11]) ? node6480 : node6477;
														assign node6477 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node6480 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node6483 = (inp[1]) ? 4'b0001 : node6484;
												assign node6484 = (inp[13]) ? 4'b0000 : 4'b0001;
							assign node6489 = (inp[2]) ? node6687 : node6490;
								assign node6490 = (inp[1]) ? node6598 : node6491;
									assign node6491 = (inp[3]) ? node6545 : node6492;
										assign node6492 = (inp[13]) ? node6516 : node6493;
											assign node6493 = (inp[10]) ? node6501 : node6494;
												assign node6494 = (inp[12]) ? node6496 : 4'b1000;
													assign node6496 = (inp[14]) ? node6498 : 4'b0000;
														assign node6498 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node6501 = (inp[7]) ? node6511 : node6502;
													assign node6502 = (inp[12]) ? node6508 : node6503;
														assign node6503 = (inp[4]) ? node6505 : 4'b1000;
															assign node6505 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6508 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node6511 = (inp[11]) ? 4'b1000 : node6512;
														assign node6512 = (inp[12]) ? 4'b1000 : 4'b1001;
											assign node6516 = (inp[4]) ? node6524 : node6517;
												assign node6517 = (inp[14]) ? node6521 : node6518;
													assign node6518 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node6521 = (inp[11]) ? 4'b0100 : 4'b1001;
												assign node6524 = (inp[7]) ? node6538 : node6525;
													assign node6525 = (inp[11]) ? node6533 : node6526;
														assign node6526 = (inp[10]) ? node6530 : node6527;
															assign node6527 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node6530 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node6533 = (inp[14]) ? node6535 : 4'b1001;
															assign node6535 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6538 = (inp[11]) ? node6540 : 4'b0000;
														assign node6540 = (inp[10]) ? 4'b0100 : node6541;
															assign node6541 = (inp[12]) ? 4'b1000 : 4'b0100;
										assign node6545 = (inp[7]) ? node6575 : node6546;
											assign node6546 = (inp[12]) ? node6560 : node6547;
												assign node6547 = (inp[4]) ? node6557 : node6548;
													assign node6548 = (inp[14]) ? node6552 : node6549;
														assign node6549 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node6552 = (inp[10]) ? node6554 : 4'b0000;
															assign node6554 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node6557 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node6560 = (inp[13]) ? node6570 : node6561;
													assign node6561 = (inp[14]) ? node6563 : 4'b0001;
														assign node6563 = (inp[4]) ? node6565 : 4'b0000;
															assign node6565 = (inp[11]) ? 4'b0001 : node6566;
																assign node6566 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node6570 = (inp[11]) ? 4'b0000 : node6571;
														assign node6571 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node6575 = (inp[4]) ? node6587 : node6576;
												assign node6576 = (inp[14]) ? node6580 : node6577;
													assign node6577 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node6580 = (inp[11]) ? node6584 : node6581;
														assign node6581 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node6584 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node6587 = (inp[13]) ? 4'b0000 : node6588;
													assign node6588 = (inp[10]) ? 4'b0000 : node6589;
														assign node6589 = (inp[14]) ? 4'b1001 : node6590;
															assign node6590 = (inp[11]) ? 4'b0000 : node6591;
																assign node6591 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node6598 = (inp[11]) ? node6654 : node6599;
										assign node6599 = (inp[14]) ? node6637 : node6600;
											assign node6600 = (inp[3]) ? node6620 : node6601;
												assign node6601 = (inp[7]) ? node6615 : node6602;
													assign node6602 = (inp[10]) ? 4'b0101 : node6603;
														assign node6603 = (inp[4]) ? node6611 : node6604;
															assign node6604 = (inp[12]) ? node6608 : node6605;
																assign node6605 = (inp[13]) ? 4'b0101 : 4'b1001;
																assign node6608 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node6611 = (inp[12]) ? 4'b0101 : 4'b1000;
													assign node6615 = (inp[13]) ? node6617 : 4'b1001;
														assign node6617 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node6620 = (inp[10]) ? node6632 : node6621;
													assign node6621 = (inp[12]) ? node6627 : node6622;
														assign node6622 = (inp[7]) ? node6624 : 4'b0001;
															assign node6624 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node6627 = (inp[13]) ? 4'b0001 : node6628;
															assign node6628 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node6632 = (inp[12]) ? node6634 : 4'b1000;
														assign node6634 = (inp[4]) ? 4'b0001 : 4'b1000;
											assign node6637 = (inp[3]) ? node6643 : node6638;
												assign node6638 = (inp[12]) ? node6640 : 4'b1000;
													assign node6640 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node6643 = (inp[4]) ? node6649 : node6644;
													assign node6644 = (inp[12]) ? node6646 : 4'b1001;
														assign node6646 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node6649 = (inp[7]) ? 4'b0000 : node6650;
														assign node6650 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node6654 = (inp[13]) ? node6670 : node6655;
											assign node6655 = (inp[4]) ? node6657 : 4'b1001;
												assign node6657 = (inp[10]) ? 4'b0001 : node6658;
													assign node6658 = (inp[3]) ? node6664 : node6659;
														assign node6659 = (inp[12]) ? node6661 : 4'b1101;
															assign node6661 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node6664 = (inp[12]) ? node6666 : 4'b1001;
															assign node6666 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node6670 = (inp[12]) ? node6680 : node6671;
												assign node6671 = (inp[3]) ? node6677 : node6672;
													assign node6672 = (inp[10]) ? node6674 : 4'b0101;
														assign node6674 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node6677 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node6680 = (inp[3]) ? node6684 : node6681;
													assign node6681 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node6684 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node6687 = (inp[3]) ? node6689 : 4'b0001;
									assign node6689 = (inp[13]) ? node6713 : node6690;
										assign node6690 = (inp[4]) ? node6692 : 4'b0001;
											assign node6692 = (inp[7]) ? 4'b0001 : node6693;
												assign node6693 = (inp[12]) ? node6699 : node6694;
													assign node6694 = (inp[10]) ? 4'b0001 : node6695;
														assign node6695 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node6699 = (inp[10]) ? node6709 : node6700;
														assign node6700 = (inp[11]) ? node6706 : node6701;
															assign node6701 = (inp[1]) ? node6703 : 4'b0001;
																assign node6703 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6706 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node6709 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node6713 = (inp[10]) ? node6731 : node6714;
											assign node6714 = (inp[1]) ? 4'b0001 : node6715;
												assign node6715 = (inp[4]) ? node6721 : node6716;
													assign node6716 = (inp[12]) ? 4'b0001 : node6717;
														assign node6717 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6721 = (inp[7]) ? node6723 : 4'b0000;
														assign node6723 = (inp[12]) ? 4'b0001 : node6724;
															assign node6724 = (inp[14]) ? node6726 : 4'b0000;
																assign node6726 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node6731 = (inp[4]) ? node6745 : node6732;
												assign node6732 = (inp[7]) ? 4'b0001 : node6733;
													assign node6733 = (inp[14]) ? node6735 : 4'b0000;
														assign node6735 = (inp[12]) ? node6737 : 4'b0000;
															assign node6737 = (inp[11]) ? node6741 : node6738;
																assign node6738 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node6741 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node6745 = (inp[14]) ? node6747 : 4'b0000;
													assign node6747 = (inp[11]) ? 4'b0000 : node6748;
														assign node6748 = (inp[7]) ? node6750 : 4'b0000;
															assign node6750 = (inp[1]) ? 4'b0000 : 4'b0001;
		assign node6754 = (inp[9]) ? node10070 : node6755;
			assign node6755 = (inp[15]) ? node8531 : node6756;
				assign node6756 = (inp[6]) ? node7224 : node6757;
					assign node6757 = (inp[0]) ? 4'b1100 : node6758;
						assign node6758 = (inp[5]) ? node6926 : node6759;
							assign node6759 = (inp[2]) ? 4'b1110 : node6760;
								assign node6760 = (inp[3]) ? node6842 : node6761;
									assign node6761 = (inp[7]) ? node6813 : node6762;
										assign node6762 = (inp[1]) ? node6788 : node6763;
											assign node6763 = (inp[13]) ? node6775 : node6764;
												assign node6764 = (inp[4]) ? node6766 : 4'b1110;
													assign node6766 = (inp[14]) ? node6772 : node6767;
														assign node6767 = (inp[10]) ? node6769 : 4'b1001;
															assign node6769 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node6772 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6775 = (inp[12]) ? node6783 : node6776;
													assign node6776 = (inp[10]) ? node6778 : 4'b0001;
														assign node6778 = (inp[14]) ? node6780 : 4'b1001;
															assign node6780 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node6783 = (inp[14]) ? node6785 : 4'b0001;
														assign node6785 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node6788 = (inp[14]) ? node6800 : node6789;
												assign node6789 = (inp[13]) ? node6795 : node6790;
													assign node6790 = (inp[10]) ? 4'b0000 : node6791;
														assign node6791 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node6795 = (inp[10]) ? 4'b1000 : node6796;
														assign node6796 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6800 = (inp[11]) ? node6808 : node6801;
													assign node6801 = (inp[13]) ? node6805 : node6802;
														assign node6802 = (inp[4]) ? 4'b1001 : 4'b1110;
														assign node6805 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6808 = (inp[12]) ? node6810 : 4'b1000;
														assign node6810 = (inp[4]) ? 4'b1000 : 4'b0000;
										assign node6813 = (inp[4]) ? node6815 : 4'b1110;
											assign node6815 = (inp[13]) ? node6827 : node6816;
												assign node6816 = (inp[12]) ? node6822 : node6817;
													assign node6817 = (inp[14]) ? node6819 : 4'b0000;
														assign node6819 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node6822 = (inp[11]) ? node6824 : 4'b1110;
														assign node6824 = (inp[10]) ? 4'b0000 : 4'b1110;
												assign node6827 = (inp[1]) ? node6831 : node6828;
													assign node6828 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node6831 = (inp[11]) ? node6837 : node6832;
														assign node6832 = (inp[14]) ? node6834 : 4'b1000;
															assign node6834 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6837 = (inp[10]) ? 4'b1000 : node6838;
															assign node6838 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node6842 = (inp[1]) ? node6892 : node6843;
										assign node6843 = (inp[13]) ? node6869 : node6844;
											assign node6844 = (inp[14]) ? node6854 : node6845;
												assign node6845 = (inp[10]) ? node6847 : 4'b1001;
													assign node6847 = (inp[12]) ? node6851 : node6848;
														assign node6848 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node6851 = (inp[11]) ? 4'b1001 : 4'b1101;
												assign node6854 = (inp[11]) ? node6864 : node6855;
													assign node6855 = (inp[12]) ? node6859 : node6856;
														assign node6856 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node6859 = (inp[7]) ? 4'b1000 : node6860;
															assign node6860 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node6864 = (inp[12]) ? 4'b1001 : node6865;
														assign node6865 = (inp[10]) ? 4'b0101 : 4'b1001;
											assign node6869 = (inp[12]) ? node6881 : node6870;
												assign node6870 = (inp[10]) ? node6872 : 4'b0101;
													assign node6872 = (inp[4]) ? node6876 : node6873;
														assign node6873 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node6876 = (inp[14]) ? node6878 : 4'b1101;
															assign node6878 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node6881 = (inp[14]) ? node6887 : node6882;
													assign node6882 = (inp[4]) ? 4'b0101 : node6883;
														assign node6883 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node6887 = (inp[11]) ? 4'b0101 : node6888;
														assign node6888 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node6892 = (inp[14]) ? node6906 : node6893;
											assign node6893 = (inp[13]) ? node6901 : node6894;
												assign node6894 = (inp[4]) ? 4'b0100 : node6895;
													assign node6895 = (inp[12]) ? node6897 : 4'b0100;
														assign node6897 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node6901 = (inp[11]) ? node6903 : 4'b1100;
													assign node6903 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node6906 = (inp[11]) ? node6916 : node6907;
												assign node6907 = (inp[7]) ? node6911 : node6908;
													assign node6908 = (inp[4]) ? 4'b1101 : 4'b0101;
													assign node6911 = (inp[12]) ? node6913 : 4'b1001;
														assign node6913 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node6916 = (inp[13]) ? node6920 : node6917;
													assign node6917 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node6920 = (inp[4]) ? 4'b1100 : node6921;
														assign node6921 = (inp[7]) ? 4'b1000 : 4'b1100;
							assign node6926 = (inp[1]) ? node7084 : node6927;
								assign node6927 = (inp[13]) ? node7009 : node6928;
									assign node6928 = (inp[11]) ? node6970 : node6929;
										assign node6929 = (inp[14]) ? node6947 : node6930;
											assign node6930 = (inp[10]) ? node6936 : node6931;
												assign node6931 = (inp[3]) ? 4'b1001 : node6932;
													assign node6932 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node6936 = (inp[3]) ? node6938 : 4'b1110;
													assign node6938 = (inp[12]) ? node6944 : node6939;
														assign node6939 = (inp[4]) ? 4'b0101 : node6940;
															assign node6940 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node6944 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node6947 = (inp[12]) ? node6961 : node6948;
												assign node6948 = (inp[10]) ? node6956 : node6949;
													assign node6949 = (inp[3]) ? node6953 : node6950;
														assign node6950 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node6953 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node6956 = (inp[3]) ? 4'b0100 : node6957;
														assign node6957 = (inp[2]) ? 4'b1110 : 4'b0100;
												assign node6961 = (inp[7]) ? node6967 : node6962;
													assign node6962 = (inp[3]) ? node6964 : 4'b1000;
														assign node6964 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node6967 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node6970 = (inp[10]) ? node6986 : node6971;
											assign node6971 = (inp[3]) ? node6977 : node6972;
												assign node6972 = (inp[7]) ? node6974 : 4'b1001;
													assign node6974 = (inp[2]) ? 4'b1110 : 4'b1101;
												assign node6977 = (inp[14]) ? node6979 : 4'b1001;
													assign node6979 = (inp[2]) ? node6981 : 4'b1101;
														assign node6981 = (inp[4]) ? node6983 : 4'b1001;
															assign node6983 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node6986 = (inp[12]) ? node6990 : node6987;
												assign node6987 = (inp[14]) ? 4'b0001 : 4'b0101;
												assign node6990 = (inp[14]) ? node6998 : node6991;
													assign node6991 = (inp[4]) ? node6993 : 4'b1001;
														assign node6993 = (inp[2]) ? 4'b1001 : node6994;
															assign node6994 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node6998 = (inp[2]) ? 4'b1101 : node6999;
														assign node6999 = (inp[4]) ? node7001 : 4'b1101;
															assign node7001 = (inp[7]) ? node7005 : node7002;
																assign node7002 = (inp[3]) ? 4'b1101 : 4'b1001;
																assign node7005 = (inp[3]) ? 4'b1001 : 4'b1101;
									assign node7009 = (inp[14]) ? node7045 : node7010;
										assign node7010 = (inp[12]) ? node7034 : node7011;
											assign node7011 = (inp[10]) ? node7025 : node7012;
												assign node7012 = (inp[3]) ? node7020 : node7013;
													assign node7013 = (inp[2]) ? 4'b1110 : node7014;
														assign node7014 = (inp[4]) ? 4'b0001 : node7015;
															assign node7015 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node7020 = (inp[4]) ? 4'b0101 : node7021;
														assign node7021 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7025 = (inp[3]) ? node7029 : node7026;
													assign node7026 = (inp[11]) ? 4'b1001 : 4'b1110;
													assign node7029 = (inp[4]) ? 4'b1101 : node7030;
														assign node7030 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node7034 = (inp[7]) ? node7038 : node7035;
												assign node7035 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node7038 = (inp[4]) ? node7042 : node7039;
													assign node7039 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node7042 = (inp[3]) ? 4'b0101 : 4'b0001;
										assign node7045 = (inp[11]) ? node7067 : node7046;
											assign node7046 = (inp[3]) ? node7056 : node7047;
												assign node7047 = (inp[7]) ? node7051 : node7048;
													assign node7048 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node7051 = (inp[4]) ? 4'b0000 : node7052;
														assign node7052 = (inp[10]) ? 4'b1100 : 4'b1110;
												assign node7056 = (inp[4]) ? node7062 : node7057;
													assign node7057 = (inp[7]) ? node7059 : 4'b0100;
														assign node7059 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7062 = (inp[12]) ? 4'b0100 : node7063;
														assign node7063 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node7067 = (inp[10]) ? node7075 : node7068;
												assign node7068 = (inp[3]) ? 4'b0101 : node7069;
													assign node7069 = (inp[4]) ? 4'b0001 : node7070;
														assign node7070 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node7075 = (inp[12]) ? node7079 : node7076;
													assign node7076 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node7079 = (inp[7]) ? node7081 : 4'b0101;
														assign node7081 = (inp[2]) ? 4'b1110 : 4'b0101;
								assign node7084 = (inp[11]) ? node7168 : node7085;
									assign node7085 = (inp[14]) ? node7119 : node7086;
										assign node7086 = (inp[13]) ? node7094 : node7087;
											assign node7087 = (inp[7]) ? node7091 : node7088;
												assign node7088 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node7091 = (inp[2]) ? 4'b1110 : 4'b0100;
											assign node7094 = (inp[10]) ? node7104 : node7095;
												assign node7095 = (inp[12]) ? node7099 : node7096;
													assign node7096 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node7099 = (inp[3]) ? node7101 : 4'b0000;
														assign node7101 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7104 = (inp[12]) ? node7112 : node7105;
													assign node7105 = (inp[4]) ? 4'b1000 : node7106;
														assign node7106 = (inp[7]) ? node7108 : 4'b1000;
															assign node7108 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node7112 = (inp[3]) ? 4'b1100 : node7113;
														assign node7113 = (inp[4]) ? 4'b1000 : node7114;
															assign node7114 = (inp[7]) ? 4'b1100 : 4'b1000;
										assign node7119 = (inp[13]) ? node7143 : node7120;
											assign node7120 = (inp[12]) ? node7132 : node7121;
												assign node7121 = (inp[10]) ? node7127 : node7122;
													assign node7122 = (inp[3]) ? 4'b1001 : node7123;
														assign node7123 = (inp[2]) ? 4'b1110 : 4'b1101;
													assign node7127 = (inp[3]) ? 4'b0101 : node7128;
														assign node7128 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node7132 = (inp[4]) ? node7134 : 4'b1001;
													assign node7134 = (inp[3]) ? node7140 : node7135;
														assign node7135 = (inp[7]) ? node7137 : 4'b1001;
															assign node7137 = (inp[2]) ? 4'b1110 : 4'b1101;
														assign node7140 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node7143 = (inp[12]) ? node7157 : node7144;
												assign node7144 = (inp[10]) ? node7148 : node7145;
													assign node7145 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node7148 = (inp[3]) ? node7152 : node7149;
														assign node7149 = (inp[7]) ? 4'b1110 : 4'b1001;
														assign node7152 = (inp[7]) ? node7154 : 4'b1101;
															assign node7154 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node7157 = (inp[3]) ? node7163 : node7158;
													assign node7158 = (inp[10]) ? 4'b0001 : node7159;
														assign node7159 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node7163 = (inp[7]) ? node7165 : 4'b0101;
														assign node7165 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node7168 = (inp[13]) ? node7192 : node7169;
										assign node7169 = (inp[3]) ? node7179 : node7170;
											assign node7170 = (inp[4]) ? 4'b0000 : node7171;
												assign node7171 = (inp[14]) ? node7173 : 4'b1110;
													assign node7173 = (inp[7]) ? node7175 : 4'b0000;
														assign node7175 = (inp[2]) ? 4'b1110 : 4'b0100;
											assign node7179 = (inp[10]) ? node7187 : node7180;
												assign node7180 = (inp[12]) ? 4'b1000 : node7181;
													assign node7181 = (inp[4]) ? 4'b0100 : node7182;
														assign node7182 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7187 = (inp[4]) ? 4'b0100 : node7188;
													assign node7188 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node7192 = (inp[12]) ? node7206 : node7193;
											assign node7193 = (inp[3]) ? node7201 : node7194;
												assign node7194 = (inp[4]) ? 4'b1000 : node7195;
													assign node7195 = (inp[7]) ? node7197 : 4'b1000;
														assign node7197 = (inp[2]) ? 4'b1110 : 4'b1100;
												assign node7201 = (inp[7]) ? node7203 : 4'b1100;
													assign node7203 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node7206 = (inp[10]) ? node7218 : node7207;
												assign node7207 = (inp[3]) ? node7213 : node7208;
													assign node7208 = (inp[7]) ? node7210 : 4'b0000;
														assign node7210 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node7213 = (inp[7]) ? node7215 : 4'b0100;
														assign node7215 = (inp[14]) ? 4'b0100 : 4'b0000;
												assign node7218 = (inp[3]) ? node7220 : 4'b1000;
													assign node7220 = (inp[2]) ? 4'b1100 : 4'b1000;
					assign node7224 = (inp[5]) ? node7816 : node7225;
						assign node7225 = (inp[0]) ? node7635 : node7226;
							assign node7226 = (inp[11]) ? node7438 : node7227;
								assign node7227 = (inp[3]) ? node7351 : node7228;
									assign node7228 = (inp[7]) ? node7282 : node7229;
										assign node7229 = (inp[2]) ? node7255 : node7230;
											assign node7230 = (inp[4]) ? node7244 : node7231;
												assign node7231 = (inp[10]) ? node7239 : node7232;
													assign node7232 = (inp[1]) ? node7236 : node7233;
														assign node7233 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node7236 = (inp[14]) ? 4'b1101 : 4'b0001;
													assign node7239 = (inp[12]) ? 4'b0001 : node7240;
														assign node7240 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node7244 = (inp[10]) ? node7250 : node7245;
													assign node7245 = (inp[13]) ? 4'b1101 : node7246;
														assign node7246 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node7250 = (inp[13]) ? 4'b0101 : node7251;
														assign node7251 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node7255 = (inp[1]) ? node7267 : node7256;
												assign node7256 = (inp[14]) ? node7264 : node7257;
													assign node7257 = (inp[12]) ? node7261 : node7258;
														assign node7258 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7261 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node7264 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node7267 = (inp[14]) ? 4'b0001 : node7268;
													assign node7268 = (inp[13]) ? node7276 : node7269;
														assign node7269 = (inp[12]) ? node7271 : 4'b0000;
															assign node7271 = (inp[10]) ? 4'b0000 : node7272;
																assign node7272 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node7276 = (inp[12]) ? node7278 : 4'b1000;
															assign node7278 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node7282 = (inp[4]) ? node7322 : node7283;
											assign node7283 = (inp[13]) ? node7303 : node7284;
												assign node7284 = (inp[12]) ? node7294 : node7285;
													assign node7285 = (inp[1]) ? node7291 : node7286;
														assign node7286 = (inp[10]) ? 4'b0101 : node7287;
															assign node7287 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node7291 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node7294 = (inp[2]) ? 4'b1101 : node7295;
														assign node7295 = (inp[14]) ? node7299 : node7296;
															assign node7296 = (inp[1]) ? 4'b0100 : 4'b1101;
															assign node7299 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node7303 = (inp[10]) ? node7313 : node7304;
													assign node7304 = (inp[12]) ? node7308 : node7305;
														assign node7305 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node7308 = (inp[14]) ? node7310 : 4'b0100;
															assign node7310 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node7313 = (inp[12]) ? node7317 : node7314;
														assign node7314 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node7317 = (inp[2]) ? node7319 : 4'b0001;
															assign node7319 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node7322 = (inp[10]) ? node7342 : node7323;
												assign node7323 = (inp[13]) ? node7333 : node7324;
													assign node7324 = (inp[2]) ? node7326 : 4'b1001;
														assign node7326 = (inp[12]) ? node7328 : 4'b1101;
															assign node7328 = (inp[1]) ? node7330 : 4'b1100;
																assign node7330 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node7333 = (inp[2]) ? node7339 : node7334;
														assign node7334 = (inp[12]) ? 4'b1001 : node7335;
															assign node7335 = (inp[1]) ? 4'b0101 : 4'b1001;
														assign node7339 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node7342 = (inp[13]) ? 4'b0101 : node7343;
													assign node7343 = (inp[2]) ? node7345 : 4'b0001;
														assign node7345 = (inp[14]) ? 4'b0000 : node7346;
															assign node7346 = (inp[1]) ? 4'b0000 : 4'b1101;
									assign node7351 = (inp[10]) ? node7397 : node7352;
										assign node7352 = (inp[1]) ? node7378 : node7353;
											assign node7353 = (inp[13]) ? node7367 : node7354;
												assign node7354 = (inp[2]) ? node7362 : node7355;
													assign node7355 = (inp[4]) ? node7357 : 4'b1101;
														assign node7357 = (inp[7]) ? 4'b1001 : node7358;
															assign node7358 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node7362 = (inp[14]) ? node7364 : 4'b1001;
														assign node7364 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node7367 = (inp[7]) ? node7371 : node7368;
													assign node7368 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node7371 = (inp[2]) ? node7375 : node7372;
														assign node7372 = (inp[14]) ? 4'b0001 : 4'b1101;
														assign node7375 = (inp[4]) ? 4'b1001 : 4'b0001;
											assign node7378 = (inp[12]) ? node7390 : node7379;
												assign node7379 = (inp[4]) ? node7385 : node7380;
													assign node7380 = (inp[13]) ? 4'b0001 : node7381;
														assign node7381 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node7385 = (inp[14]) ? 4'b1100 : node7386;
														assign node7386 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node7390 = (inp[2]) ? 4'b1001 : node7391;
													assign node7391 = (inp[4]) ? 4'b1001 : node7392;
														assign node7392 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node7397 = (inp[4]) ? node7417 : node7398;
											assign node7398 = (inp[1]) ? node7408 : node7399;
												assign node7399 = (inp[14]) ? 4'b0001 : node7400;
													assign node7400 = (inp[7]) ? node7404 : node7401;
														assign node7401 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node7404 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node7408 = (inp[12]) ? 4'b0001 : node7409;
													assign node7409 = (inp[2]) ? node7413 : node7410;
														assign node7410 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node7413 = (inp[13]) ? 4'b1001 : 4'b0000;
											assign node7417 = (inp[13]) ? node7427 : node7418;
												assign node7418 = (inp[12]) ? node7422 : node7419;
													assign node7419 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7422 = (inp[1]) ? 4'b1000 : node7423;
														assign node7423 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node7427 = (inp[12]) ? node7429 : 4'b1101;
													assign node7429 = (inp[2]) ? 4'b0101 : node7430;
														assign node7430 = (inp[14]) ? node7434 : node7431;
															assign node7431 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node7434 = (inp[7]) ? 4'b1001 : 4'b0100;
								assign node7438 = (inp[1]) ? node7544 : node7439;
									assign node7439 = (inp[13]) ? node7489 : node7440;
										assign node7440 = (inp[3]) ? node7462 : node7441;
											assign node7441 = (inp[2]) ? node7455 : node7442;
												assign node7442 = (inp[10]) ? node7448 : node7443;
													assign node7443 = (inp[4]) ? node7445 : 4'b1101;
														assign node7445 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7448 = (inp[12]) ? 4'b0000 : node7449;
														assign node7449 = (inp[7]) ? 4'b1000 : node7450;
															assign node7450 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node7455 = (inp[4]) ? node7457 : 4'b1101;
													assign node7457 = (inp[7]) ? node7459 : 4'b1001;
														assign node7459 = (inp[14]) ? 4'b1101 : 4'b0001;
											assign node7462 = (inp[7]) ? node7474 : node7463;
												assign node7463 = (inp[4]) ? node7471 : node7464;
													assign node7464 = (inp[10]) ? node7468 : node7465;
														assign node7465 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node7468 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7471 = (inp[10]) ? 4'b1100 : 4'b0001;
												assign node7474 = (inp[12]) ? node7480 : node7475;
													assign node7475 = (inp[2]) ? 4'b0000 : node7476;
														assign node7476 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7480 = (inp[14]) ? node7486 : node7481;
														assign node7481 = (inp[4]) ? node7483 : 4'b1001;
															assign node7483 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node7486 = (inp[2]) ? 4'b0000 : 4'b0100;
										assign node7489 = (inp[4]) ? node7511 : node7490;
											assign node7490 = (inp[2]) ? node7502 : node7491;
												assign node7491 = (inp[3]) ? node7497 : node7492;
													assign node7492 = (inp[12]) ? 4'b0101 : node7493;
														assign node7493 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node7497 = (inp[10]) ? node7499 : 4'b1000;
														assign node7499 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node7502 = (inp[3]) ? node7508 : node7503;
													assign node7503 = (inp[12]) ? 4'b0001 : node7504;
														assign node7504 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node7508 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node7511 = (inp[2]) ? node7525 : node7512;
												assign node7512 = (inp[3]) ? node7518 : node7513;
													assign node7513 = (inp[10]) ? 4'b1100 : node7514;
														assign node7514 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node7518 = (inp[10]) ? 4'b0101 : node7519;
														assign node7519 = (inp[12]) ? 4'b0101 : node7520;
															assign node7520 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node7525 = (inp[3]) ? node7531 : node7526;
													assign node7526 = (inp[7]) ? 4'b0001 : node7527;
														assign node7527 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7531 = (inp[14]) ? node7539 : node7532;
														assign node7532 = (inp[10]) ? node7536 : node7533;
															assign node7533 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node7536 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7539 = (inp[12]) ? node7541 : 4'b0100;
															assign node7541 = (inp[10]) ? 4'b0100 : 4'b1100;
									assign node7544 = (inp[10]) ? node7590 : node7545;
										assign node7545 = (inp[4]) ? node7565 : node7546;
											assign node7546 = (inp[7]) ? node7554 : node7547;
												assign node7547 = (inp[13]) ? node7549 : 4'b0000;
													assign node7549 = (inp[14]) ? 4'b0000 : node7550;
														assign node7550 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node7554 = (inp[3]) ? node7560 : node7555;
													assign node7555 = (inp[12]) ? node7557 : 4'b0100;
														assign node7557 = (inp[2]) ? 4'b0100 : 4'b1100;
													assign node7560 = (inp[13]) ? 4'b0000 : node7561;
														assign node7561 = (inp[2]) ? 4'b0000 : 4'b0100;
											assign node7565 = (inp[13]) ? node7577 : node7566;
												assign node7566 = (inp[7]) ? 4'b0000 : node7567;
													assign node7567 = (inp[3]) ? node7571 : node7568;
														assign node7568 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node7571 = (inp[2]) ? 4'b0100 : node7572;
															assign node7572 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node7577 = (inp[3]) ? node7583 : node7578;
													assign node7578 = (inp[2]) ? node7580 : 4'b0100;
														assign node7580 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node7583 = (inp[2]) ? 4'b0100 : node7584;
														assign node7584 = (inp[12]) ? node7586 : 4'b0100;
															assign node7586 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node7590 = (inp[4]) ? node7614 : node7591;
											assign node7591 = (inp[13]) ? node7603 : node7592;
												assign node7592 = (inp[7]) ? node7596 : node7593;
													assign node7593 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node7596 = (inp[2]) ? node7600 : node7597;
														assign node7597 = (inp[3]) ? 4'b1100 : 4'b0100;
														assign node7600 = (inp[14]) ? 4'b0000 : 4'b0100;
												assign node7603 = (inp[14]) ? 4'b1000 : node7604;
													assign node7604 = (inp[3]) ? 4'b1000 : node7605;
														assign node7605 = (inp[12]) ? node7607 : 4'b1100;
															assign node7607 = (inp[2]) ? node7609 : 4'b1000;
																assign node7609 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node7614 = (inp[13]) ? node7630 : node7615;
												assign node7615 = (inp[7]) ? node7623 : node7616;
													assign node7616 = (inp[3]) ? node7620 : node7617;
														assign node7617 = (inp[14]) ? 4'b1100 : 4'b0000;
														assign node7620 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node7623 = (inp[12]) ? node7625 : 4'b0000;
														assign node7625 = (inp[14]) ? node7627 : 4'b1000;
															assign node7627 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node7630 = (inp[3]) ? 4'b1100 : node7631;
													assign node7631 = (inp[2]) ? 4'b1000 : 4'b1100;
							assign node7635 = (inp[2]) ? 4'b1100 : node7636;
								assign node7636 = (inp[1]) ? node7728 : node7637;
									assign node7637 = (inp[13]) ? node7679 : node7638;
										assign node7638 = (inp[12]) ? node7658 : node7639;
											assign node7639 = (inp[10]) ? node7651 : node7640;
												assign node7640 = (inp[3]) ? node7646 : node7641;
													assign node7641 = (inp[14]) ? 4'b1100 : node7642;
														assign node7642 = (inp[7]) ? 4'b1100 : 4'b1001;
													assign node7646 = (inp[14]) ? node7648 : 4'b1101;
														assign node7648 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node7651 = (inp[14]) ? node7653 : 4'b0001;
													assign node7653 = (inp[3]) ? node7655 : 4'b0000;
														assign node7655 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node7658 = (inp[3]) ? node7666 : node7659;
												assign node7659 = (inp[4]) ? node7661 : 4'b1100;
													assign node7661 = (inp[7]) ? 4'b1100 : node7662;
														assign node7662 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node7666 = (inp[7]) ? node7676 : node7667;
													assign node7667 = (inp[4]) ? node7671 : node7668;
														assign node7668 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7671 = (inp[14]) ? node7673 : 4'b1101;
															assign node7673 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node7676 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node7679 = (inp[10]) ? node7697 : node7680;
											assign node7680 = (inp[4]) ? node7690 : node7681;
												assign node7681 = (inp[12]) ? node7683 : 4'b0001;
													assign node7683 = (inp[7]) ? node7687 : node7684;
														assign node7684 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node7687 = (inp[3]) ? 4'b0000 : 4'b1100;
												assign node7690 = (inp[3]) ? node7692 : 4'b0001;
													assign node7692 = (inp[11]) ? 4'b0101 : node7693;
														assign node7693 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node7697 = (inp[12]) ? node7713 : node7698;
												assign node7698 = (inp[11]) ? node7706 : node7699;
													assign node7699 = (inp[3]) ? node7703 : node7700;
														assign node7700 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node7703 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7706 = (inp[7]) ? node7708 : 4'b1001;
														assign node7708 = (inp[4]) ? 4'b1001 : node7709;
															assign node7709 = (inp[3]) ? 4'b1001 : 4'b1100;
												assign node7713 = (inp[11]) ? node7723 : node7714;
													assign node7714 = (inp[14]) ? node7716 : 4'b0001;
														assign node7716 = (inp[3]) ? node7718 : 4'b0000;
															assign node7718 = (inp[4]) ? 4'b0100 : node7719;
																assign node7719 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7723 = (inp[14]) ? node7725 : 4'b1100;
														assign node7725 = (inp[3]) ? 4'b0101 : 4'b0001;
									assign node7728 = (inp[14]) ? node7760 : node7729;
										assign node7729 = (inp[13]) ? node7737 : node7730;
											assign node7730 = (inp[3]) ? node7732 : 4'b0000;
												assign node7732 = (inp[10]) ? 4'b0100 : node7733;
													assign node7733 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node7737 = (inp[3]) ? node7751 : node7738;
												assign node7738 = (inp[4]) ? node7746 : node7739;
													assign node7739 = (inp[7]) ? 4'b1100 : node7740;
														assign node7740 = (inp[12]) ? node7742 : 4'b1000;
															assign node7742 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node7746 = (inp[10]) ? 4'b1000 : node7747;
														assign node7747 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node7751 = (inp[12]) ? node7757 : node7752;
													assign node7752 = (inp[7]) ? node7754 : 4'b1100;
														assign node7754 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node7757 = (inp[7]) ? 4'b0100 : 4'b1100;
										assign node7760 = (inp[11]) ? node7782 : node7761;
											assign node7761 = (inp[13]) ? node7765 : node7762;
												assign node7762 = (inp[3]) ? 4'b1001 : 4'b1100;
												assign node7765 = (inp[12]) ? node7775 : node7766;
													assign node7766 = (inp[10]) ? node7768 : 4'b0001;
														assign node7768 = (inp[3]) ? node7770 : 4'b1001;
															assign node7770 = (inp[7]) ? node7772 : 4'b1101;
																assign node7772 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node7775 = (inp[3]) ? node7777 : 4'b0001;
														assign node7777 = (inp[7]) ? node7779 : 4'b0101;
															assign node7779 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node7782 = (inp[13]) ? node7792 : node7783;
												assign node7783 = (inp[10]) ? node7787 : node7784;
													assign node7784 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node7787 = (inp[7]) ? 4'b0000 : node7788;
														assign node7788 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node7792 = (inp[12]) ? node7804 : node7793;
													assign node7793 = (inp[4]) ? 4'b1000 : node7794;
														assign node7794 = (inp[10]) ? 4'b1100 : node7795;
															assign node7795 = (inp[7]) ? node7799 : node7796;
																assign node7796 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node7799 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node7804 = (inp[3]) ? node7810 : node7805;
														assign node7805 = (inp[7]) ? node7807 : 4'b0000;
															assign node7807 = (inp[4]) ? 4'b0000 : 4'b1100;
														assign node7810 = (inp[4]) ? 4'b1100 : node7811;
															assign node7811 = (inp[7]) ? 4'b1000 : 4'b1100;
						assign node7816 = (inp[3]) ? node8198 : node7817;
							assign node7817 = (inp[4]) ? node7995 : node7818;
								assign node7818 = (inp[7]) ? node7920 : node7819;
									assign node7819 = (inp[1]) ? node7863 : node7820;
										assign node7820 = (inp[2]) ? node7838 : node7821;
											assign node7821 = (inp[0]) ? node7827 : node7822;
												assign node7822 = (inp[13]) ? node7824 : 4'b0000;
													assign node7824 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node7827 = (inp[10]) ? node7833 : node7828;
													assign node7828 = (inp[14]) ? node7830 : 4'b1000;
														assign node7830 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node7833 = (inp[12]) ? node7835 : 4'b1000;
														assign node7835 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node7838 = (inp[13]) ? node7850 : node7839;
												assign node7839 = (inp[0]) ? 4'b1100 : node7840;
													assign node7840 = (inp[10]) ? node7844 : node7841;
														assign node7841 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node7844 = (inp[14]) ? 4'b1001 : node7845;
															assign node7845 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node7850 = (inp[10]) ? node7860 : node7851;
													assign node7851 = (inp[0]) ? node7855 : node7852;
														assign node7852 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7855 = (inp[11]) ? 4'b0001 : node7856;
															assign node7856 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node7860 = (inp[0]) ? 4'b0001 : 4'b0101;
										assign node7863 = (inp[11]) ? node7897 : node7864;
											assign node7864 = (inp[10]) ? node7884 : node7865;
												assign node7865 = (inp[2]) ? node7873 : node7866;
													assign node7866 = (inp[13]) ? node7870 : node7867;
														assign node7867 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7870 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node7873 = (inp[14]) ? node7879 : node7874;
														assign node7874 = (inp[13]) ? 4'b1001 : node7875;
															assign node7875 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node7879 = (inp[13]) ? node7881 : 4'b1100;
															assign node7881 = (inp[0]) ? 4'b0001 : 4'b1000;
												assign node7884 = (inp[12]) ? node7892 : node7885;
													assign node7885 = (inp[2]) ? node7889 : node7886;
														assign node7886 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7889 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node7892 = (inp[2]) ? node7894 : 4'b0001;
														assign node7894 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node7897 = (inp[10]) ? node7913 : node7898;
												assign node7898 = (inp[0]) ? node7906 : node7899;
													assign node7899 = (inp[13]) ? node7903 : node7900;
														assign node7900 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node7903 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node7906 = (inp[2]) ? node7908 : 4'b0000;
														assign node7908 = (inp[13]) ? 4'b0000 : node7909;
															assign node7909 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node7913 = (inp[2]) ? node7915 : 4'b1000;
													assign node7915 = (inp[13]) ? node7917 : 4'b0000;
														assign node7917 = (inp[0]) ? 4'b1000 : 4'b1100;
									assign node7920 = (inp[0]) ? node7974 : node7921;
										assign node7921 = (inp[2]) ? node7945 : node7922;
											assign node7922 = (inp[1]) ? node7934 : node7923;
												assign node7923 = (inp[11]) ? node7929 : node7924;
													assign node7924 = (inp[10]) ? node7926 : 4'b0100;
														assign node7926 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node7929 = (inp[13]) ? node7931 : 4'b0000;
														assign node7931 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node7934 = (inp[14]) ? node7938 : node7935;
													assign node7935 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node7938 = (inp[11]) ? 4'b1000 : node7939;
														assign node7939 = (inp[13]) ? 4'b1000 : node7940;
															assign node7940 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node7945 = (inp[13]) ? node7957 : node7946;
												assign node7946 = (inp[11]) ? node7954 : node7947;
													assign node7947 = (inp[10]) ? node7949 : 4'b1101;
														assign node7949 = (inp[1]) ? node7951 : 4'b0101;
															assign node7951 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node7954 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node7957 = (inp[14]) ? node7971 : node7958;
													assign node7958 = (inp[12]) ? node7968 : node7959;
														assign node7959 = (inp[10]) ? 4'b0001 : node7960;
															assign node7960 = (inp[1]) ? node7964 : node7961;
																assign node7961 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node7964 = (inp[11]) ? 4'b0000 : 4'b1001;
														assign node7968 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node7971 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node7974 = (inp[2]) ? 4'b1100 : node7975;
											assign node7975 = (inp[13]) ? node7985 : node7976;
												assign node7976 = (inp[1]) ? node7978 : 4'b1101;
													assign node7978 = (inp[10]) ? 4'b0100 : node7979;
														assign node7979 = (inp[14]) ? 4'b1101 : node7980;
															assign node7980 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node7985 = (inp[11]) ? node7991 : node7986;
													assign node7986 = (inp[12]) ? node7988 : 4'b0001;
														assign node7988 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node7991 = (inp[10]) ? 4'b1000 : 4'b0000;
								assign node7995 = (inp[11]) ? node8123 : node7996;
									assign node7996 = (inp[2]) ? node8056 : node7997;
										assign node7997 = (inp[10]) ? node8029 : node7998;
											assign node7998 = (inp[12]) ? node8012 : node7999;
												assign node7999 = (inp[0]) ? node8005 : node8000;
													assign node8000 = (inp[1]) ? 4'b1001 : node8001;
														assign node8001 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8005 = (inp[1]) ? node8007 : 4'b1001;
														assign node8007 = (inp[13]) ? node8009 : 4'b0101;
															assign node8009 = (inp[7]) ? 4'b0101 : 4'b1001;
												assign node8012 = (inp[14]) ? node8020 : node8013;
													assign node8013 = (inp[0]) ? 4'b0000 : node8014;
														assign node8014 = (inp[1]) ? node8016 : 4'b1001;
															assign node8016 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node8020 = (inp[0]) ? node8024 : node8021;
														assign node8021 = (inp[1]) ? 4'b0001 : 4'b1100;
														assign node8024 = (inp[7]) ? 4'b1001 : node8025;
															assign node8025 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node8029 = (inp[13]) ? node8041 : node8030;
												assign node8030 = (inp[7]) ? node8034 : node8031;
													assign node8031 = (inp[0]) ? 4'b0101 : 4'b0001;
													assign node8034 = (inp[1]) ? 4'b1001 : node8035;
														assign node8035 = (inp[14]) ? node8037 : 4'b0001;
															assign node8037 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node8041 = (inp[12]) ? node8049 : node8042;
													assign node8042 = (inp[1]) ? node8046 : node8043;
														assign node8043 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node8046 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node8049 = (inp[0]) ? node8051 : 4'b0001;
														assign node8051 = (inp[7]) ? node8053 : 4'b0000;
															assign node8053 = (inp[1]) ? 4'b0000 : 4'b0101;
										assign node8056 = (inp[10]) ? node8088 : node8057;
											assign node8057 = (inp[13]) ? node8079 : node8058;
												assign node8058 = (inp[0]) ? node8074 : node8059;
													assign node8059 = (inp[1]) ? node8069 : node8060;
														assign node8060 = (inp[14]) ? node8064 : node8061;
															assign node8061 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node8064 = (inp[12]) ? 4'b1101 : node8065;
																assign node8065 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node8069 = (inp[7]) ? node8071 : 4'b0000;
															assign node8071 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node8074 = (inp[7]) ? 4'b1100 : node8075;
														assign node8075 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node8079 = (inp[0]) ? node8083 : node8080;
													assign node8080 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node8083 = (inp[12]) ? node8085 : 4'b0001;
														assign node8085 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node8088 = (inp[1]) ? node8112 : node8089;
												assign node8089 = (inp[14]) ? node8097 : node8090;
													assign node8090 = (inp[7]) ? node8094 : node8091;
														assign node8091 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8094 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node8097 = (inp[7]) ? node8105 : node8098;
														assign node8098 = (inp[13]) ? node8100 : 4'b1000;
															assign node8100 = (inp[0]) ? node8102 : 4'b1000;
																assign node8102 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8105 = (inp[0]) ? node8109 : node8106;
															assign node8106 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node8109 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8112 = (inp[12]) ? node8114 : 4'b1000;
													assign node8114 = (inp[14]) ? node8116 : 4'b0000;
														assign node8116 = (inp[0]) ? node8120 : node8117;
															assign node8117 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node8120 = (inp[13]) ? 4'b0001 : 4'b1001;
									assign node8123 = (inp[1]) ? node8167 : node8124;
										assign node8124 = (inp[0]) ? node8150 : node8125;
											assign node8125 = (inp[13]) ? node8141 : node8126;
												assign node8126 = (inp[14]) ? node8132 : node8127;
													assign node8127 = (inp[2]) ? 4'b0000 : node8128;
														assign node8128 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node8132 = (inp[10]) ? 4'b0101 : node8133;
														assign node8133 = (inp[7]) ? node8137 : node8134;
															assign node8134 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node8137 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node8141 = (inp[10]) ? 4'b0100 : node8142;
													assign node8142 = (inp[7]) ? node8146 : node8143;
														assign node8143 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node8146 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node8150 = (inp[2]) ? node8160 : node8151;
												assign node8151 = (inp[10]) ? node8155 : node8152;
													assign node8152 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node8155 = (inp[13]) ? 4'b0001 : node8156;
														assign node8156 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node8160 = (inp[13]) ? 4'b0001 : node8161;
													assign node8161 = (inp[10]) ? node8163 : 4'b1001;
														assign node8163 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node8167 = (inp[7]) ? node8181 : node8168;
											assign node8168 = (inp[10]) ? node8176 : node8169;
												assign node8169 = (inp[2]) ? 4'b1000 : node8170;
													assign node8170 = (inp[14]) ? 4'b0100 : node8171;
														assign node8171 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8176 = (inp[13]) ? 4'b1000 : node8177;
													assign node8177 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node8181 = (inp[13]) ? node8193 : node8182;
												assign node8182 = (inp[0]) ? node8188 : node8183;
													assign node8183 = (inp[2]) ? node8185 : 4'b0100;
														assign node8185 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node8188 = (inp[2]) ? 4'b0000 : node8189;
														assign node8189 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node8193 = (inp[10]) ? 4'b1000 : node8194;
													assign node8194 = (inp[12]) ? 4'b0100 : 4'b0000;
							assign node8198 = (inp[4]) ? node8376 : node8199;
								assign node8199 = (inp[11]) ? node8303 : node8200;
									assign node8200 = (inp[7]) ? node8250 : node8201;
										assign node8201 = (inp[2]) ? node8217 : node8202;
											assign node8202 = (inp[13]) ? node8212 : node8203;
												assign node8203 = (inp[0]) ? node8207 : node8204;
													assign node8204 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node8207 = (inp[1]) ? node8209 : 4'b0000;
														assign node8209 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8212 = (inp[1]) ? 4'b0000 : node8213;
													assign node8213 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node8217 = (inp[13]) ? node8233 : node8218;
												assign node8218 = (inp[12]) ? node8226 : node8219;
													assign node8219 = (inp[0]) ? node8221 : 4'b1001;
														assign node8221 = (inp[1]) ? 4'b0001 : node8222;
															assign node8222 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node8226 = (inp[10]) ? node8230 : node8227;
														assign node8227 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node8230 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node8233 = (inp[0]) ? node8239 : node8234;
													assign node8234 = (inp[10]) ? node8236 : 4'b0000;
														assign node8236 = (inp[14]) ? 4'b0000 : 4'b1001;
													assign node8239 = (inp[10]) ? node8245 : node8240;
														assign node8240 = (inp[1]) ? node8242 : 4'b1001;
															assign node8242 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8245 = (inp[12]) ? node8247 : 4'b1000;
															assign node8247 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node8250 = (inp[1]) ? node8278 : node8251;
											assign node8251 = (inp[13]) ? node8261 : node8252;
												assign node8252 = (inp[12]) ? node8258 : node8253;
													assign node8253 = (inp[0]) ? node8255 : 4'b1001;
														assign node8255 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node8258 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node8261 = (inp[14]) ? node8273 : node8262;
													assign node8262 = (inp[2]) ? node8268 : node8263;
														assign node8263 = (inp[0]) ? node8265 : 4'b0001;
															assign node8265 = (inp[12]) ? 4'b1000 : 4'b1001;
														assign node8268 = (inp[10]) ? node8270 : 4'b1000;
															assign node8270 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node8273 = (inp[2]) ? node8275 : 4'b0001;
														assign node8275 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node8278 = (inp[13]) ? node8286 : node8279;
												assign node8279 = (inp[0]) ? 4'b0000 : node8280;
													assign node8280 = (inp[14]) ? node8282 : 4'b1000;
														assign node8282 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node8286 = (inp[10]) ? node8292 : node8287;
													assign node8287 = (inp[2]) ? node8289 : 4'b0001;
														assign node8289 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node8292 = (inp[14]) ? 4'b1001 : node8293;
														assign node8293 = (inp[0]) ? node8297 : node8294;
															assign node8294 = (inp[12]) ? 4'b1000 : 4'b0001;
															assign node8297 = (inp[2]) ? node8299 : 4'b0001;
																assign node8299 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node8303 = (inp[1]) ? node8357 : node8304;
										assign node8304 = (inp[0]) ? node8332 : node8305;
											assign node8305 = (inp[2]) ? node8321 : node8306;
												assign node8306 = (inp[7]) ? node8312 : node8307;
													assign node8307 = (inp[14]) ? 4'b1001 : node8308;
														assign node8308 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node8312 = (inp[12]) ? node8318 : node8313;
														assign node8313 = (inp[14]) ? node8315 : 4'b0000;
															assign node8315 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8318 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node8321 = (inp[10]) ? node8323 : 4'b0001;
													assign node8323 = (inp[13]) ? node8327 : node8324;
														assign node8324 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node8327 = (inp[7]) ? 4'b0001 : node8328;
															assign node8328 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node8332 = (inp[2]) ? node8342 : node8333;
												assign node8333 = (inp[7]) ? node8339 : node8334;
													assign node8334 = (inp[10]) ? node8336 : 4'b1001;
														assign node8336 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node8339 = (inp[10]) ? 4'b1001 : 4'b0000;
												assign node8342 = (inp[7]) ? node8352 : node8343;
													assign node8343 = (inp[10]) ? node8347 : node8344;
														assign node8344 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node8347 = (inp[13]) ? 4'b0001 : node8348;
															assign node8348 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node8352 = (inp[13]) ? node8354 : 4'b1001;
														assign node8354 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node8357 = (inp[2]) ? node8367 : node8358;
											assign node8358 = (inp[7]) ? 4'b1000 : node8359;
												assign node8359 = (inp[14]) ? 4'b1000 : node8360;
													assign node8360 = (inp[10]) ? node8362 : 4'b1000;
														assign node8362 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node8367 = (inp[10]) ? node8369 : 4'b0000;
												assign node8369 = (inp[13]) ? 4'b1000 : node8370;
													assign node8370 = (inp[7]) ? 4'b0000 : node8371;
														assign node8371 = (inp[0]) ? 4'b1000 : 4'b0000;
								assign node8376 = (inp[11]) ? node8474 : node8377;
									assign node8377 = (inp[13]) ? node8427 : node8378;
										assign node8378 = (inp[7]) ? node8408 : node8379;
											assign node8379 = (inp[2]) ? node8401 : node8380;
												assign node8380 = (inp[14]) ? node8390 : node8381;
													assign node8381 = (inp[10]) ? 4'b0000 : node8382;
														assign node8382 = (inp[0]) ? node8386 : node8383;
															assign node8383 = (inp[1]) ? 4'b0001 : 4'b1000;
															assign node8386 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node8390 = (inp[0]) ? node8392 : 4'b0000;
														assign node8392 = (inp[10]) ? node8396 : node8393;
															assign node8393 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node8396 = (inp[12]) ? node8398 : 4'b0001;
																assign node8398 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node8401 = (inp[1]) ? 4'b1000 : node8402;
													assign node8402 = (inp[14]) ? node8404 : 4'b0001;
														assign node8404 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node8408 = (inp[1]) ? node8410 : 4'b0001;
												assign node8410 = (inp[2]) ? node8416 : node8411;
													assign node8411 = (inp[14]) ? 4'b0001 : node8412;
														assign node8412 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node8416 = (inp[12]) ? node8422 : node8417;
														assign node8417 = (inp[0]) ? node8419 : 4'b0000;
															assign node8419 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8422 = (inp[0]) ? node8424 : 4'b0001;
															assign node8424 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node8427 = (inp[1]) ? node8459 : node8428;
											assign node8428 = (inp[2]) ? node8448 : node8429;
												assign node8429 = (inp[0]) ? node8435 : node8430;
													assign node8430 = (inp[14]) ? node8432 : 4'b0000;
														assign node8432 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node8435 = (inp[10]) ? node8443 : node8436;
														assign node8436 = (inp[7]) ? node8440 : node8437;
															assign node8437 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8440 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node8443 = (inp[14]) ? 4'b0001 : node8444;
															assign node8444 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node8448 = (inp[0]) ? 4'b0000 : node8449;
													assign node8449 = (inp[7]) ? node8455 : node8450;
														assign node8450 = (inp[14]) ? node8452 : 4'b0000;
															assign node8452 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8455 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node8459 = (inp[10]) ? 4'b0000 : node8460;
												assign node8460 = (inp[14]) ? 4'b0001 : node8461;
													assign node8461 = (inp[12]) ? node8463 : 4'b0000;
														assign node8463 = (inp[7]) ? node8467 : node8464;
															assign node8464 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node8467 = (inp[0]) ? 4'b0000 : node8468;
																assign node8468 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node8474 = (inp[13]) ? node8520 : node8475;
										assign node8475 = (inp[10]) ? node8503 : node8476;
											assign node8476 = (inp[0]) ? node8494 : node8477;
												assign node8477 = (inp[2]) ? node8487 : node8478;
													assign node8478 = (inp[12]) ? node8482 : node8479;
														assign node8479 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node8482 = (inp[14]) ? 4'b1000 : node8483;
															assign node8483 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node8487 = (inp[7]) ? 4'b0000 : node8488;
														assign node8488 = (inp[12]) ? node8490 : 4'b1000;
															assign node8490 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node8494 = (inp[1]) ? node8496 : 4'b1000;
													assign node8496 = (inp[2]) ? node8498 : 4'b0000;
														assign node8498 = (inp[12]) ? node8500 : 4'b1000;
															assign node8500 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node8503 = (inp[1]) ? 4'b0000 : node8504;
												assign node8504 = (inp[0]) ? node8512 : node8505;
													assign node8505 = (inp[12]) ? node8507 : 4'b0001;
														assign node8507 = (inp[2]) ? node8509 : 4'b0001;
															assign node8509 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node8512 = (inp[7]) ? 4'b0000 : node8513;
														assign node8513 = (inp[12]) ? node8515 : 4'b0000;
															assign node8515 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node8520 = (inp[14]) ? node8522 : 4'b0000;
											assign node8522 = (inp[10]) ? 4'b0000 : node8523;
												assign node8523 = (inp[0]) ? 4'b0000 : node8524;
													assign node8524 = (inp[2]) ? 4'b0000 : node8525;
														assign node8525 = (inp[1]) ? 4'b0000 : 4'b0001;
				assign node8531 = (inp[0]) ? node9697 : node8532;
					assign node8532 = (inp[6]) ? node8876 : node8533;
						assign node8533 = (inp[5]) ? node8609 : node8534;
							assign node8534 = (inp[3]) ? node8536 : 4'b1010;
								assign node8536 = (inp[2]) ? 4'b1010 : node8537;
									assign node8537 = (inp[7]) ? node8581 : node8538;
										assign node8538 = (inp[13]) ? node8560 : node8539;
											assign node8539 = (inp[4]) ? node8547 : node8540;
												assign node8540 = (inp[12]) ? 4'b1010 : node8541;
													assign node8541 = (inp[10]) ? node8543 : 4'b1010;
														assign node8543 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node8547 = (inp[11]) ? 4'b1001 : node8548;
													assign node8548 = (inp[10]) ? node8552 : node8549;
														assign node8549 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8552 = (inp[14]) ? node8554 : 4'b0000;
															assign node8554 = (inp[12]) ? 4'b1001 : node8555;
																assign node8555 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node8560 = (inp[12]) ? node8570 : node8561;
												assign node8561 = (inp[1]) ? node8565 : node8562;
													assign node8562 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8565 = (inp[14]) ? node8567 : 4'b1000;
														assign node8567 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node8570 = (inp[10]) ? 4'b0001 : node8571;
													assign node8571 = (inp[1]) ? node8577 : node8572;
														assign node8572 = (inp[11]) ? 4'b0001 : node8573;
															assign node8573 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node8577 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node8581 = (inp[4]) ? node8583 : 4'b1010;
											assign node8583 = (inp[1]) ? node8593 : node8584;
												assign node8584 = (inp[12]) ? 4'b1010 : node8585;
													assign node8585 = (inp[10]) ? node8587 : 4'b1010;
														assign node8587 = (inp[13]) ? node8589 : 4'b0001;
															assign node8589 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node8593 = (inp[11]) ? node8605 : node8594;
													assign node8594 = (inp[13]) ? node8602 : node8595;
														assign node8595 = (inp[12]) ? node8597 : 4'b0001;
															assign node8597 = (inp[14]) ? 4'b1010 : node8598;
																assign node8598 = (inp[10]) ? 4'b0000 : 4'b1010;
														assign node8602 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node8605 = (inp[13]) ? 4'b1000 : 4'b0000;
							assign node8609 = (inp[2]) ? node8787 : node8610;
								assign node8610 = (inp[1]) ? node8694 : node8611;
									assign node8611 = (inp[14]) ? node8651 : node8612;
										assign node8612 = (inp[13]) ? node8630 : node8613;
											assign node8613 = (inp[10]) ? node8619 : node8614;
												assign node8614 = (inp[3]) ? node8616 : 4'b1001;
													assign node8616 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8619 = (inp[12]) ? node8627 : node8620;
													assign node8620 = (inp[3]) ? 4'b0001 : node8621;
														assign node8621 = (inp[11]) ? 4'b0101 : node8622;
															assign node8622 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node8627 = (inp[3]) ? 4'b1101 : 4'b1001;
											assign node8630 = (inp[10]) ? node8642 : node8631;
												assign node8631 = (inp[3]) ? node8637 : node8632;
													assign node8632 = (inp[4]) ? 4'b0101 : node8633;
														assign node8633 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node8637 = (inp[7]) ? node8639 : 4'b0001;
														assign node8639 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node8642 = (inp[12]) ? node8646 : node8643;
													assign node8643 = (inp[11]) ? 4'b1001 : 4'b1101;
													assign node8646 = (inp[4]) ? node8648 : 4'b0001;
														assign node8648 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node8651 = (inp[11]) ? node8675 : node8652;
											assign node8652 = (inp[3]) ? node8668 : node8653;
												assign node8653 = (inp[4]) ? node8661 : node8654;
													assign node8654 = (inp[7]) ? 4'b0000 : node8655;
														assign node8655 = (inp[13]) ? 4'b0100 : node8656;
															assign node8656 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node8661 = (inp[7]) ? node8663 : 4'b1100;
														assign node8663 = (inp[10]) ? node8665 : 4'b0100;
															assign node8665 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node8668 = (inp[10]) ? node8670 : 4'b1100;
													assign node8670 = (inp[13]) ? node8672 : 4'b0000;
														assign node8672 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node8675 = (inp[13]) ? node8685 : node8676;
												assign node8676 = (inp[3]) ? node8680 : node8677;
													assign node8677 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node8680 = (inp[7]) ? 4'b1101 : node8681;
														assign node8681 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8685 = (inp[3]) ? 4'b0001 : node8686;
													assign node8686 = (inp[10]) ? 4'b1101 : node8687;
														assign node8687 = (inp[12]) ? node8689 : 4'b0101;
															assign node8689 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node8694 = (inp[11]) ? node8748 : node8695;
										assign node8695 = (inp[14]) ? node8727 : node8696;
											assign node8696 = (inp[3]) ? node8706 : node8697;
												assign node8697 = (inp[7]) ? node8703 : node8698;
													assign node8698 = (inp[13]) ? 4'b0100 : node8699;
														assign node8699 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node8703 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node8706 = (inp[4]) ? node8720 : node8707;
													assign node8707 = (inp[7]) ? node8715 : node8708;
														assign node8708 = (inp[10]) ? node8712 : node8709;
															assign node8709 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node8712 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node8715 = (inp[12]) ? 4'b1100 : node8716;
															assign node8716 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node8720 = (inp[10]) ? 4'b0000 : node8721;
														assign node8721 = (inp[7]) ? 4'b1000 : node8722;
															assign node8722 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node8727 = (inp[13]) ? node8739 : node8728;
												assign node8728 = (inp[10]) ? node8734 : node8729;
													assign node8729 = (inp[7]) ? node8731 : 4'b1001;
														assign node8731 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node8734 = (inp[12]) ? node8736 : 4'b0101;
														assign node8736 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node8739 = (inp[12]) ? 4'b0001 : node8740;
													assign node8740 = (inp[10]) ? node8744 : node8741;
														assign node8741 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node8744 = (inp[3]) ? 4'b1001 : 4'b1101;
										assign node8748 = (inp[13]) ? node8774 : node8749;
											assign node8749 = (inp[12]) ? node8761 : node8750;
												assign node8750 = (inp[3]) ? node8756 : node8751;
													assign node8751 = (inp[4]) ? 4'b0100 : node8752;
														assign node8752 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node8756 = (inp[4]) ? 4'b0000 : node8757;
														assign node8757 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node8761 = (inp[10]) ? node8767 : node8762;
													assign node8762 = (inp[3]) ? 4'b1100 : node8763;
														assign node8763 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node8767 = (inp[4]) ? 4'b0100 : node8768;
														assign node8768 = (inp[3]) ? node8770 : 4'b0000;
															assign node8770 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node8774 = (inp[3]) ? node8784 : node8775;
												assign node8775 = (inp[7]) ? node8781 : node8776;
													assign node8776 = (inp[12]) ? node8778 : 4'b1100;
														assign node8778 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node8781 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node8784 = (inp[12]) ? 4'b1100 : 4'b1000;
								assign node8787 = (inp[3]) ? node8789 : 4'b1010;
									assign node8789 = (inp[4]) ? node8819 : node8790;
										assign node8790 = (inp[7]) ? 4'b1010 : node8791;
											assign node8791 = (inp[13]) ? node8803 : node8792;
												assign node8792 = (inp[12]) ? node8798 : node8793;
													assign node8793 = (inp[10]) ? 4'b0001 : node8794;
														assign node8794 = (inp[14]) ? 4'b1010 : 4'b0000;
													assign node8798 = (inp[10]) ? node8800 : 4'b1010;
														assign node8800 = (inp[11]) ? 4'b0000 : 4'b1010;
												assign node8803 = (inp[1]) ? node8811 : node8804;
													assign node8804 = (inp[11]) ? node8806 : 4'b0000;
														assign node8806 = (inp[12]) ? 4'b0001 : node8807;
															assign node8807 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8811 = (inp[11]) ? node8813 : 4'b0001;
														assign node8813 = (inp[12]) ? node8815 : 4'b1000;
															assign node8815 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node8819 = (inp[1]) ? node8847 : node8820;
											assign node8820 = (inp[13]) ? node8836 : node8821;
												assign node8821 = (inp[7]) ? node8829 : node8822;
													assign node8822 = (inp[11]) ? node8826 : node8823;
														assign node8823 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8826 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node8829 = (inp[12]) ? 4'b1010 : node8830;
														assign node8830 = (inp[10]) ? node8832 : 4'b1010;
															assign node8832 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node8836 = (inp[10]) ? node8842 : node8837;
													assign node8837 = (inp[11]) ? 4'b0001 : node8838;
														assign node8838 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8842 = (inp[12]) ? 4'b0001 : node8843;
														assign node8843 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node8847 = (inp[11]) ? node8865 : node8848;
												assign node8848 = (inp[14]) ? node8856 : node8849;
													assign node8849 = (inp[10]) ? node8853 : node8850;
														assign node8850 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node8853 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8856 = (inp[13]) ? node8860 : node8857;
														assign node8857 = (inp[7]) ? 4'b1010 : 4'b1001;
														assign node8860 = (inp[12]) ? 4'b0001 : node8861;
															assign node8861 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node8865 = (inp[13]) ? node8871 : node8866;
													assign node8866 = (inp[12]) ? node8868 : 4'b0000;
														assign node8868 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node8871 = (inp[12]) ? node8873 : 4'b1000;
														assign node8873 = (inp[10]) ? 4'b1000 : 4'b0000;
						assign node8876 = (inp[5]) ? node9300 : node8877;
							assign node8877 = (inp[11]) ? node9109 : node8878;
								assign node8878 = (inp[2]) ? node8994 : node8879;
									assign node8879 = (inp[10]) ? node8931 : node8880;
										assign node8880 = (inp[3]) ? node8912 : node8881;
											assign node8881 = (inp[13]) ? node8903 : node8882;
												assign node8882 = (inp[7]) ? node8894 : node8883;
													assign node8883 = (inp[4]) ? 4'b1100 : node8884;
														assign node8884 = (inp[12]) ? node8888 : node8885;
															assign node8885 = (inp[1]) ? 4'b0100 : 4'b1001;
															assign node8888 = (inp[1]) ? node8890 : 4'b1000;
																assign node8890 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8894 = (inp[1]) ? node8898 : node8895;
														assign node8895 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8898 = (inp[14]) ? 4'b1001 : node8899;
															assign node8899 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node8903 = (inp[7]) ? node8907 : node8904;
													assign node8904 = (inp[14]) ? 4'b1001 : 4'b1100;
													assign node8907 = (inp[4]) ? node8909 : 4'b0000;
														assign node8909 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node8912 = (inp[1]) ? node8920 : node8913;
												assign node8913 = (inp[4]) ? 4'b1101 : node8914;
													assign node8914 = (inp[13]) ? node8916 : 4'b1001;
														assign node8916 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node8920 = (inp[12]) ? node8924 : node8921;
													assign node8921 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node8924 = (inp[7]) ? 4'b1101 : node8925;
														assign node8925 = (inp[4]) ? 4'b1001 : node8926;
															assign node8926 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node8931 = (inp[1]) ? node8963 : node8932;
											assign node8932 = (inp[3]) ? node8952 : node8933;
												assign node8933 = (inp[12]) ? node8947 : node8934;
													assign node8934 = (inp[14]) ? node8940 : node8935;
														assign node8935 = (inp[13]) ? 4'b1101 : node8936;
															assign node8936 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node8940 = (inp[13]) ? 4'b1000 : node8941;
															assign node8941 = (inp[4]) ? 4'b0100 : node8942;
																assign node8942 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node8947 = (inp[4]) ? 4'b0001 : node8948;
														assign node8948 = (inp[13]) ? 4'b0101 : 4'b1001;
												assign node8952 = (inp[4]) ? node8958 : node8953;
													assign node8953 = (inp[13]) ? 4'b0101 : node8954;
														assign node8954 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node8958 = (inp[7]) ? node8960 : 4'b0001;
														assign node8960 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node8963 = (inp[12]) ? node8981 : node8964;
												assign node8964 = (inp[4]) ? node8974 : node8965;
													assign node8965 = (inp[13]) ? node8969 : node8966;
														assign node8966 = (inp[3]) ? 4'b1001 : 4'b0001;
														assign node8969 = (inp[3]) ? 4'b1101 : node8970;
															assign node8970 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node8974 = (inp[7]) ? 4'b1101 : node8975;
														assign node8975 = (inp[14]) ? node8977 : 4'b1001;
															assign node8977 = (inp[3]) ? 4'b1000 : 4'b1001;
												assign node8981 = (inp[14]) ? node8985 : node8982;
													assign node8982 = (inp[3]) ? 4'b0101 : 4'b0100;
													assign node8985 = (inp[3]) ? node8991 : node8986;
														assign node8986 = (inp[7]) ? 4'b1001 : node8987;
															assign node8987 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node8991 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node8994 = (inp[13]) ? node9048 : node8995;
										assign node8995 = (inp[12]) ? node9023 : node8996;
											assign node8996 = (inp[10]) ? node9010 : node8997;
												assign node8997 = (inp[14]) ? node9003 : node8998;
													assign node8998 = (inp[1]) ? node9000 : 4'b1101;
														assign node9000 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node9003 = (inp[1]) ? node9007 : node9004;
														assign node9004 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9007 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node9010 = (inp[3]) ? node9018 : node9011;
													assign node9011 = (inp[1]) ? node9015 : node9012;
														assign node9012 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node9015 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node9018 = (inp[7]) ? node9020 : 4'b0001;
														assign node9020 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node9023 = (inp[3]) ? node9041 : node9024;
												assign node9024 = (inp[14]) ? node9034 : node9025;
													assign node9025 = (inp[1]) ? node9027 : 4'b1001;
														assign node9027 = (inp[10]) ? 4'b0100 : node9028;
															assign node9028 = (inp[7]) ? 4'b1000 : node9029;
																assign node9029 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9034 = (inp[1]) ? node9036 : 4'b1000;
														assign node9036 = (inp[7]) ? 4'b1001 : node9037;
															assign node9037 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node9041 = (inp[14]) ? node9045 : node9042;
													assign node9042 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node9045 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node9048 = (inp[10]) ? node9078 : node9049;
											assign node9049 = (inp[3]) ? node9065 : node9050;
												assign node9050 = (inp[14]) ? node9058 : node9051;
													assign node9051 = (inp[1]) ? 4'b1100 : node9052;
														assign node9052 = (inp[7]) ? node9054 : 4'b0101;
															assign node9054 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node9058 = (inp[1]) ? 4'b0101 : node9059;
														assign node9059 = (inp[4]) ? 4'b0100 : node9060;
															assign node9060 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node9065 = (inp[14]) ? node9073 : node9066;
													assign node9066 = (inp[12]) ? node9068 : 4'b1100;
														assign node9068 = (inp[7]) ? node9070 : 4'b0000;
															assign node9070 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node9073 = (inp[1]) ? 4'b0001 : node9074;
														assign node9074 = (inp[4]) ? 4'b1001 : 4'b0000;
											assign node9078 = (inp[12]) ? node9096 : node9079;
												assign node9079 = (inp[4]) ? node9087 : node9080;
													assign node9080 = (inp[14]) ? node9084 : node9081;
														assign node9081 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node9084 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node9087 = (inp[3]) ? 4'b1001 : node9088;
														assign node9088 = (inp[14]) ? node9092 : node9089;
															assign node9089 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node9092 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node9096 = (inp[14]) ? node9102 : node9097;
													assign node9097 = (inp[1]) ? 4'b1000 : node9098;
														assign node9098 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node9102 = (inp[1]) ? node9106 : node9103;
														assign node9103 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9106 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node9109 = (inp[1]) ? node9217 : node9110;
									assign node9110 = (inp[3]) ? node9154 : node9111;
										assign node9111 = (inp[13]) ? node9129 : node9112;
											assign node9112 = (inp[10]) ? node9120 : node9113;
												assign node9113 = (inp[4]) ? node9115 : 4'b1001;
													assign node9115 = (inp[7]) ? 4'b1001 : node9116;
														assign node9116 = (inp[12]) ? 4'b1101 : 4'b0000;
												assign node9120 = (inp[4]) ? node9124 : node9121;
													assign node9121 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9124 = (inp[7]) ? 4'b1001 : node9125;
														assign node9125 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node9129 = (inp[12]) ? node9147 : node9130;
												assign node9130 = (inp[10]) ? node9136 : node9131;
													assign node9131 = (inp[4]) ? 4'b0000 : node9132;
														assign node9132 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9136 = (inp[2]) ? node9142 : node9137;
														assign node9137 = (inp[4]) ? 4'b1000 : node9138;
															assign node9138 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node9142 = (inp[7]) ? node9144 : 4'b1101;
															assign node9144 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node9147 = (inp[10]) ? node9149 : 4'b0101;
													assign node9149 = (inp[4]) ? 4'b0000 : node9150;
														assign node9150 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node9154 = (inp[13]) ? node9182 : node9155;
											assign node9155 = (inp[2]) ? node9175 : node9156;
												assign node9156 = (inp[4]) ? node9168 : node9157;
													assign node9157 = (inp[7]) ? node9163 : node9158;
														assign node9158 = (inp[10]) ? 4'b0100 : node9159;
															assign node9159 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node9163 = (inp[12]) ? node9165 : 4'b0000;
															assign node9165 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node9168 = (inp[7]) ? node9170 : 4'b0000;
														assign node9170 = (inp[10]) ? 4'b1100 : node9171;
															assign node9171 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node9175 = (inp[4]) ? node9177 : 4'b1101;
													assign node9177 = (inp[7]) ? node9179 : 4'b0000;
														assign node9179 = (inp[14]) ? 4'b1101 : 4'b0001;
											assign node9182 = (inp[4]) ? node9194 : node9183;
												assign node9183 = (inp[2]) ? node9189 : node9184;
													assign node9184 = (inp[7]) ? 4'b1000 : node9185;
														assign node9185 = (inp[14]) ? 4'b1100 : 4'b0100;
													assign node9189 = (inp[7]) ? node9191 : 4'b0001;
														assign node9191 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node9194 = (inp[2]) ? node9202 : node9195;
													assign node9195 = (inp[7]) ? node9199 : node9196;
														assign node9196 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node9199 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node9202 = (inp[7]) ? node9210 : node9203;
														assign node9203 = (inp[10]) ? node9207 : node9204;
															assign node9204 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node9207 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9210 = (inp[12]) ? node9214 : node9211;
															assign node9211 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node9214 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node9217 = (inp[10]) ? node9265 : node9218;
										assign node9218 = (inp[12]) ? node9240 : node9219;
											assign node9219 = (inp[13]) ? node9231 : node9220;
												assign node9220 = (inp[4]) ? node9226 : node9221;
													assign node9221 = (inp[3]) ? 4'b0000 : node9222;
														assign node9222 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node9226 = (inp[14]) ? 4'b0100 : node9227;
														assign node9227 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node9231 = (inp[4]) ? node9235 : node9232;
													assign node9232 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node9235 = (inp[2]) ? node9237 : 4'b0000;
														assign node9237 = (inp[3]) ? 4'b0000 : 4'b1100;
											assign node9240 = (inp[13]) ? node9252 : node9241;
												assign node9241 = (inp[3]) ? node9247 : node9242;
													assign node9242 = (inp[4]) ? node9244 : 4'b1000;
														assign node9244 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node9247 = (inp[2]) ? 4'b1100 : node9248;
														assign node9248 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node9252 = (inp[4]) ? node9260 : node9253;
													assign node9253 = (inp[2]) ? node9255 : 4'b0100;
														assign node9255 = (inp[7]) ? 4'b0000 : node9256;
															assign node9256 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node9260 = (inp[7]) ? node9262 : 4'b1000;
														assign node9262 = (inp[2]) ? 4'b0100 : 4'b0000;
										assign node9265 = (inp[13]) ? node9287 : node9266;
											assign node9266 = (inp[3]) ? node9272 : node9267;
												assign node9267 = (inp[4]) ? 4'b0100 : node9268;
													assign node9268 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9272 = (inp[7]) ? node9282 : node9273;
													assign node9273 = (inp[12]) ? node9279 : node9274;
														assign node9274 = (inp[14]) ? 4'b0000 : node9275;
															assign node9275 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node9279 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node9282 = (inp[12]) ? 4'b0100 : node9283;
														assign node9283 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node9287 = (inp[4]) ? node9295 : node9288;
												assign node9288 = (inp[3]) ? node9292 : node9289;
													assign node9289 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9292 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node9295 = (inp[2]) ? node9297 : 4'b1000;
													assign node9297 = (inp[3]) ? 4'b1000 : 4'b1100;
							assign node9300 = (inp[3]) ? node9520 : node9301;
								assign node9301 = (inp[4]) ? node9417 : node9302;
									assign node9302 = (inp[11]) ? node9364 : node9303;
										assign node9303 = (inp[2]) ? node9337 : node9304;
											assign node9304 = (inp[13]) ? node9322 : node9305;
												assign node9305 = (inp[12]) ? node9317 : node9306;
													assign node9306 = (inp[1]) ? node9314 : node9307;
														assign node9307 = (inp[14]) ? 4'b1001 : node9308;
															assign node9308 = (inp[7]) ? node9310 : 4'b0100;
																assign node9310 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node9314 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node9317 = (inp[14]) ? 4'b0101 : node9318;
														assign node9318 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node9322 = (inp[7]) ? node9330 : node9323;
													assign node9323 = (inp[14]) ? 4'b1000 : node9324;
														assign node9324 = (inp[1]) ? node9326 : 4'b0100;
															assign node9326 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node9330 = (inp[1]) ? node9334 : node9331;
														assign node9331 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node9334 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node9337 = (inp[7]) ? node9353 : node9338;
												assign node9338 = (inp[10]) ? node9342 : node9339;
													assign node9339 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node9342 = (inp[13]) ? node9344 : 4'b0101;
														assign node9344 = (inp[1]) ? node9348 : node9345;
															assign node9345 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node9348 = (inp[14]) ? 4'b0000 : node9349;
																assign node9349 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9353 = (inp[10]) ? node9359 : node9354;
													assign node9354 = (inp[13]) ? 4'b1001 : node9355;
														assign node9355 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node9359 = (inp[12]) ? 4'b0101 : node9360;
														assign node9360 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node9364 = (inp[1]) ? node9392 : node9365;
											assign node9365 = (inp[2]) ? node9377 : node9366;
												assign node9366 = (inp[13]) ? node9372 : node9367;
													assign node9367 = (inp[7]) ? 4'b1001 : node9368;
														assign node9368 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node9372 = (inp[7]) ? node9374 : 4'b0000;
														assign node9374 = (inp[10]) ? 4'b0000 : 4'b1101;
												assign node9377 = (inp[10]) ? node9383 : node9378;
													assign node9378 = (inp[12]) ? node9380 : 4'b0100;
														assign node9380 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node9383 = (inp[7]) ? node9387 : node9384;
														assign node9384 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node9387 = (inp[12]) ? 4'b0100 : node9388;
															assign node9388 = (inp[13]) ? 4'b1100 : 4'b1000;
											assign node9392 = (inp[13]) ? node9410 : node9393;
												assign node9393 = (inp[7]) ? node9401 : node9394;
													assign node9394 = (inp[12]) ? 4'b0100 : node9395;
														assign node9395 = (inp[14]) ? node9397 : 4'b0100;
															assign node9397 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node9401 = (inp[2]) ? node9407 : node9402;
														assign node9402 = (inp[10]) ? 4'b0100 : node9403;
															assign node9403 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9407 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node9410 = (inp[7]) ? node9414 : node9411;
													assign node9411 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node9414 = (inp[2]) ? 4'b1100 : 4'b1000;
									assign node9417 = (inp[1]) ? node9471 : node9418;
										assign node9418 = (inp[10]) ? node9442 : node9419;
											assign node9419 = (inp[11]) ? node9433 : node9420;
												assign node9420 = (inp[13]) ? node9428 : node9421;
													assign node9421 = (inp[14]) ? node9425 : node9422;
														assign node9422 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node9425 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node9428 = (inp[2]) ? 4'b0100 : node9429;
														assign node9429 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node9433 = (inp[13]) ? node9439 : node9434;
													assign node9434 = (inp[2]) ? 4'b0001 : node9435;
														assign node9435 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node9439 = (inp[14]) ? 4'b0000 : 4'b1001;
											assign node9442 = (inp[13]) ? node9456 : node9443;
												assign node9443 = (inp[2]) ? node9451 : node9444;
													assign node9444 = (inp[7]) ? 4'b0100 : node9445;
														assign node9445 = (inp[12]) ? node9447 : 4'b1001;
															assign node9447 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9451 = (inp[7]) ? 4'b1001 : node9452;
														assign node9452 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node9456 = (inp[2]) ? node9468 : node9457;
													assign node9457 = (inp[12]) ? node9463 : node9458;
														assign node9458 = (inp[7]) ? node9460 : 4'b1001;
															assign node9460 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9463 = (inp[7]) ? node9465 : 4'b1000;
															assign node9465 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9468 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node9471 = (inp[13]) ? node9497 : node9472;
											assign node9472 = (inp[10]) ? node9484 : node9473;
												assign node9473 = (inp[12]) ? node9477 : node9474;
													assign node9474 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node9477 = (inp[7]) ? node9479 : 4'b0000;
														assign node9479 = (inp[14]) ? 4'b0000 : node9480;
															assign node9480 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node9484 = (inp[11]) ? node9494 : node9485;
													assign node9485 = (inp[7]) ? node9491 : node9486;
														assign node9486 = (inp[12]) ? 4'b1000 : node9487;
															assign node9487 = (inp[2]) ? 4'b0100 : 4'b1001;
														assign node9491 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node9494 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node9497 = (inp[11]) ? node9511 : node9498;
												assign node9498 = (inp[2]) ? node9506 : node9499;
													assign node9499 = (inp[14]) ? node9501 : 4'b0000;
														assign node9501 = (inp[12]) ? node9503 : 4'b0001;
															assign node9503 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node9506 = (inp[12]) ? node9508 : 4'b1000;
														assign node9508 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node9511 = (inp[2]) ? 4'b1000 : node9512;
													assign node9512 = (inp[10]) ? 4'b1000 : node9513;
														assign node9513 = (inp[12]) ? 4'b0000 : node9514;
															assign node9514 = (inp[7]) ? 4'b1000 : 4'b0000;
								assign node9520 = (inp[4]) ? node9626 : node9521;
									assign node9521 = (inp[11]) ? node9573 : node9522;
										assign node9522 = (inp[10]) ? node9558 : node9523;
											assign node9523 = (inp[1]) ? node9539 : node9524;
												assign node9524 = (inp[2]) ? node9534 : node9525;
													assign node9525 = (inp[13]) ? node9529 : node9526;
														assign node9526 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node9529 = (inp[7]) ? 4'b0000 : node9530;
															assign node9530 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node9534 = (inp[12]) ? node9536 : 4'b0001;
														assign node9536 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9539 = (inp[2]) ? node9549 : node9540;
													assign node9540 = (inp[12]) ? node9546 : node9541;
														assign node9541 = (inp[13]) ? 4'b0000 : node9542;
															assign node9542 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9546 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9549 = (inp[13]) ? node9553 : node9550;
														assign node9550 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9553 = (inp[14]) ? node9555 : 4'b1001;
															assign node9555 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node9558 = (inp[2]) ? node9560 : 4'b0000;
												assign node9560 = (inp[13]) ? node9568 : node9561;
													assign node9561 = (inp[14]) ? node9563 : 4'b0001;
														assign node9563 = (inp[1]) ? node9565 : 4'b0000;
															assign node9565 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9568 = (inp[14]) ? node9570 : 4'b0000;
														assign node9570 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node9573 = (inp[1]) ? node9607 : node9574;
											assign node9574 = (inp[12]) ? node9596 : node9575;
												assign node9575 = (inp[7]) ? node9589 : node9576;
													assign node9576 = (inp[10]) ? node9582 : node9577;
														assign node9577 = (inp[14]) ? 4'b1001 : node9578;
															assign node9578 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node9582 = (inp[2]) ? node9586 : node9583;
															assign node9583 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node9586 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node9589 = (inp[13]) ? node9591 : 4'b1000;
														assign node9591 = (inp[2]) ? node9593 : 4'b0001;
															assign node9593 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node9596 = (inp[10]) ? node9600 : node9597;
													assign node9597 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node9600 = (inp[7]) ? 4'b0001 : node9601;
														assign node9601 = (inp[2]) ? node9603 : 4'b1000;
															assign node9603 = (inp[13]) ? 4'b1000 : 4'b0001;
											assign node9607 = (inp[10]) ? node9619 : node9608;
												assign node9608 = (inp[13]) ? node9614 : node9609;
													assign node9609 = (inp[12]) ? 4'b0000 : node9610;
														assign node9610 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node9614 = (inp[2]) ? node9616 : 4'b0000;
														assign node9616 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node9619 = (inp[13]) ? 4'b1000 : node9620;
													assign node9620 = (inp[7]) ? 4'b1000 : node9621;
														assign node9621 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node9626 = (inp[13]) ? node9672 : node9627;
										assign node9627 = (inp[10]) ? node9659 : node9628;
											assign node9628 = (inp[1]) ? node9646 : node9629;
												assign node9629 = (inp[7]) ? node9635 : node9630;
													assign node9630 = (inp[11]) ? node9632 : 4'b0001;
														assign node9632 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node9635 = (inp[2]) ? node9641 : node9636;
														assign node9636 = (inp[12]) ? 4'b0000 : node9637;
															assign node9637 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9641 = (inp[12]) ? node9643 : 4'b0000;
															assign node9643 = (inp[11]) ? 4'b1001 : 4'b0000;
												assign node9646 = (inp[11]) ? node9652 : node9647;
													assign node9647 = (inp[2]) ? node9649 : 4'b1000;
														assign node9649 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node9652 = (inp[12]) ? 4'b1000 : node9653;
														assign node9653 = (inp[7]) ? node9655 : 4'b0000;
															assign node9655 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node9659 = (inp[1]) ? node9669 : node9660;
												assign node9660 = (inp[7]) ? node9664 : node9661;
													assign node9661 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node9664 = (inp[12]) ? node9666 : 4'b1000;
														assign node9666 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node9669 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node9672 = (inp[10]) ? 4'b0000 : node9673;
											assign node9673 = (inp[12]) ? node9681 : node9674;
												assign node9674 = (inp[2]) ? node9676 : 4'b0000;
													assign node9676 = (inp[7]) ? 4'b0000 : node9677;
														assign node9677 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node9681 = (inp[11]) ? node9687 : node9682;
													assign node9682 = (inp[2]) ? 4'b0001 : node9683;
														assign node9683 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node9687 = (inp[1]) ? 4'b0000 : node9688;
														assign node9688 = (inp[14]) ? node9690 : 4'b0000;
															assign node9690 = (inp[7]) ? node9692 : 4'b0001;
																assign node9692 = (inp[2]) ? 4'b0000 : 4'b0001;
					assign node9697 = (inp[6]) ? node9699 : 4'b1000;
						assign node9699 = (inp[5]) ? node9775 : node9700;
							assign node9700 = (inp[3]) ? node9702 : 4'b1000;
								assign node9702 = (inp[2]) ? 4'b1000 : node9703;
									assign node9703 = (inp[4]) ? node9719 : node9704;
										assign node9704 = (inp[7]) ? 4'b1000 : node9705;
											assign node9705 = (inp[12]) ? 4'b1000 : node9706;
												assign node9706 = (inp[1]) ? node9714 : node9707;
													assign node9707 = (inp[13]) ? node9711 : node9708;
														assign node9708 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node9711 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node9714 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node9719 = (inp[13]) ? node9753 : node9720;
											assign node9720 = (inp[7]) ? node9738 : node9721;
												assign node9721 = (inp[10]) ? node9729 : node9722;
													assign node9722 = (inp[14]) ? node9726 : node9723;
														assign node9723 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node9726 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node9729 = (inp[12]) ? node9733 : node9730;
														assign node9730 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9733 = (inp[1]) ? node9735 : 4'b1001;
															assign node9735 = (inp[14]) ? 4'b1001 : 4'b0000;
												assign node9738 = (inp[1]) ? node9744 : node9739;
													assign node9739 = (inp[14]) ? node9741 : 4'b1000;
														assign node9741 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node9744 = (inp[12]) ? node9746 : 4'b0000;
														assign node9746 = (inp[11]) ? 4'b0000 : node9747;
															assign node9747 = (inp[10]) ? node9749 : 4'b1000;
																assign node9749 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node9753 = (inp[12]) ? node9763 : node9754;
												assign node9754 = (inp[10]) ? node9758 : node9755;
													assign node9755 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node9758 = (inp[1]) ? node9760 : 4'b1001;
														assign node9760 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node9763 = (inp[11]) ? 4'b0000 : node9764;
													assign node9764 = (inp[1]) ? node9768 : node9765;
														assign node9765 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9768 = (inp[14]) ? 4'b0001 : node9769;
															assign node9769 = (inp[7]) ? 4'b0000 : 4'b1000;
							assign node9775 = (inp[2]) ? node9995 : node9776;
								assign node9776 = (inp[3]) ? node9896 : node9777;
									assign node9777 = (inp[1]) ? node9851 : node9778;
										assign node9778 = (inp[14]) ? node9816 : node9779;
											assign node9779 = (inp[11]) ? node9799 : node9780;
												assign node9780 = (inp[4]) ? node9792 : node9781;
													assign node9781 = (inp[7]) ? node9787 : node9782;
														assign node9782 = (inp[12]) ? 4'b1001 : node9783;
															assign node9783 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node9787 = (inp[12]) ? node9789 : 4'b1001;
															assign node9789 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node9792 = (inp[10]) ? 4'b0001 : node9793;
														assign node9793 = (inp[7]) ? 4'b0101 : node9794;
															assign node9794 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node9799 = (inp[13]) ? node9809 : node9800;
													assign node9800 = (inp[12]) ? node9804 : node9801;
														assign node9801 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node9804 = (inp[7]) ? 4'b1001 : node9805;
															assign node9805 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node9809 = (inp[4]) ? node9813 : node9810;
														assign node9810 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node9813 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node9816 = (inp[11]) ? node9838 : node9817;
												assign node9817 = (inp[4]) ? node9831 : node9818;
													assign node9818 = (inp[7]) ? node9824 : node9819;
														assign node9819 = (inp[12]) ? 4'b0100 : node9820;
															assign node9820 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node9824 = (inp[13]) ? node9826 : 4'b1000;
															assign node9826 = (inp[12]) ? 4'b0000 : node9827;
																assign node9827 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node9831 = (inp[10]) ? node9833 : 4'b1001;
														assign node9833 = (inp[7]) ? node9835 : 4'b0001;
															assign node9835 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node9838 = (inp[4]) ? node9844 : node9839;
													assign node9839 = (inp[7]) ? 4'b0001 : node9840;
														assign node9840 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node9844 = (inp[7]) ? 4'b1001 : node9845;
														assign node9845 = (inp[12]) ? 4'b1000 : node9846;
															assign node9846 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node9851 = (inp[11]) ? node9877 : node9852;
											assign node9852 = (inp[14]) ? node9868 : node9853;
												assign node9853 = (inp[13]) ? node9859 : node9854;
													assign node9854 = (inp[4]) ? node9856 : 4'b0100;
														assign node9856 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node9859 = (inp[4]) ? 4'b1001 : node9860;
														assign node9860 = (inp[7]) ? 4'b1000 : node9861;
															assign node9861 = (inp[10]) ? 4'b1100 : node9862;
																assign node9862 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node9868 = (inp[13]) ? node9872 : node9869;
													assign node9869 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node9872 = (inp[10]) ? node9874 : 4'b0001;
														assign node9874 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node9877 = (inp[4]) ? node9887 : node9878;
												assign node9878 = (inp[7]) ? node9884 : node9879;
													assign node9879 = (inp[12]) ? 4'b1000 : node9880;
														assign node9880 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node9884 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node9887 = (inp[14]) ? node9893 : node9888;
													assign node9888 = (inp[10]) ? 4'b1000 : node9889;
														assign node9889 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node9893 = (inp[10]) ? 4'b0100 : 4'b0000;
									assign node9896 = (inp[4]) ? node9956 : node9897;
										assign node9897 = (inp[1]) ? node9933 : node9898;
											assign node9898 = (inp[13]) ? node9922 : node9899;
												assign node9899 = (inp[7]) ? node9913 : node9900;
													assign node9900 = (inp[12]) ? node9904 : node9901;
														assign node9901 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9904 = (inp[14]) ? node9910 : node9905;
															assign node9905 = (inp[10]) ? node9907 : 4'b1001;
																assign node9907 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node9910 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node9913 = (inp[11]) ? node9917 : node9914;
														assign node9914 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9917 = (inp[10]) ? node9919 : 4'b0000;
															assign node9919 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node9922 = (inp[10]) ? node9930 : node9923;
													assign node9923 = (inp[7]) ? node9925 : 4'b0000;
														assign node9925 = (inp[12]) ? 4'b0001 : node9926;
															assign node9926 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node9930 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node9933 = (inp[13]) ? node9947 : node9934;
												assign node9934 = (inp[11]) ? node9942 : node9935;
													assign node9935 = (inp[12]) ? 4'b1000 : node9936;
														assign node9936 = (inp[7]) ? 4'b0001 : node9937;
															assign node9937 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9942 = (inp[10]) ? 4'b0000 : node9943;
														assign node9943 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node9947 = (inp[11]) ? 4'b1000 : node9948;
													assign node9948 = (inp[12]) ? node9950 : 4'b1000;
														assign node9950 = (inp[7]) ? 4'b1001 : node9951;
															assign node9951 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node9956 = (inp[13]) ? node9976 : node9957;
											assign node9957 = (inp[10]) ? node9969 : node9958;
												assign node9958 = (inp[12]) ? node9966 : node9959;
													assign node9959 = (inp[7]) ? 4'b0001 : node9960;
														assign node9960 = (inp[11]) ? 4'b1000 : node9961;
															assign node9961 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9966 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node9969 = (inp[7]) ? node9973 : node9970;
													assign node9970 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node9973 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node9976 = (inp[11]) ? 4'b0000 : node9977;
												assign node9977 = (inp[1]) ? 4'b0000 : node9978;
													assign node9978 = (inp[12]) ? node9980 : 4'b0000;
														assign node9980 = (inp[14]) ? node9988 : node9981;
															assign node9981 = (inp[10]) ? node9985 : node9982;
																assign node9982 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node9985 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node9988 = (inp[7]) ? node9990 : 4'b0000;
																assign node9990 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node9995 = (inp[3]) ? node9997 : 4'b1000;
									assign node9997 = (inp[4]) ? node10017 : node9998;
										assign node9998 = (inp[7]) ? 4'b1000 : node9999;
											assign node9999 = (inp[12]) ? node10011 : node10000;
												assign node10000 = (inp[1]) ? node10008 : node10001;
													assign node10001 = (inp[14]) ? 4'b0000 : node10002;
														assign node10002 = (inp[11]) ? node10004 : 4'b0001;
															assign node10004 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node10008 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node10011 = (inp[13]) ? node10013 : 4'b1000;
													assign node10013 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node10017 = (inp[13]) ? node10049 : node10018;
											assign node10018 = (inp[1]) ? node10030 : node10019;
												assign node10019 = (inp[10]) ? node10025 : node10020;
													assign node10020 = (inp[7]) ? 4'b1000 : node10021;
														assign node10021 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node10025 = (inp[11]) ? node10027 : 4'b0001;
														assign node10027 = (inp[7]) ? 4'b0001 : 4'b1000;
												assign node10030 = (inp[12]) ? node10038 : node10031;
													assign node10031 = (inp[11]) ? 4'b0000 : node10032;
														assign node10032 = (inp[10]) ? 4'b0000 : node10033;
															assign node10033 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10038 = (inp[10]) ? node10042 : node10039;
														assign node10039 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node10042 = (inp[7]) ? node10046 : node10043;
															assign node10043 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node10046 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node10049 = (inp[11]) ? node10061 : node10050;
												assign node10050 = (inp[14]) ? node10052 : 4'b0001;
													assign node10052 = (inp[10]) ? 4'b0000 : node10053;
														assign node10053 = (inp[7]) ? 4'b0001 : node10054;
															assign node10054 = (inp[1]) ? node10056 : 4'b0000;
																assign node10056 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node10061 = (inp[14]) ? 4'b0000 : node10062;
													assign node10062 = (inp[12]) ? node10064 : 4'b0000;
														assign node10064 = (inp[10]) ? 4'b0000 : node10065;
															assign node10065 = (inp[1]) ? 4'b0000 : 4'b0001;
			assign node10070 = (inp[15]) ? node11862 : node10071;
				assign node10071 = (inp[6]) ? node10529 : node10072;
					assign node10072 = (inp[0]) ? 4'b0100 : node10073;
						assign node10073 = (inp[2]) ? node10383 : node10074;
							assign node10074 = (inp[3]) ? node10228 : node10075;
								assign node10075 = (inp[5]) ? node10137 : node10076;
									assign node10076 = (inp[7]) ? node10126 : node10077;
										assign node10077 = (inp[4]) ? node10097 : node10078;
											assign node10078 = (inp[13]) ? node10080 : 4'b0110;
												assign node10080 = (inp[10]) ? node10082 : 4'b0110;
													assign node10082 = (inp[12]) ? node10090 : node10083;
														assign node10083 = (inp[1]) ? node10087 : node10084;
															assign node10084 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10087 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node10090 = (inp[1]) ? node10092 : 4'b0110;
															assign node10092 = (inp[14]) ? node10094 : 4'b0000;
																assign node10094 = (inp[11]) ? 4'b0000 : 4'b0110;
											assign node10097 = (inp[1]) ? node10111 : node10098;
												assign node10098 = (inp[11]) ? node10104 : node10099;
													assign node10099 = (inp[12]) ? 4'b0000 : node10100;
														assign node10100 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node10104 = (inp[13]) ? node10106 : 4'b0001;
														assign node10106 = (inp[12]) ? 4'b1001 : node10107;
															assign node10107 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node10111 = (inp[14]) ? node10119 : node10112;
													assign node10112 = (inp[11]) ? node10114 : 4'b0000;
														assign node10114 = (inp[13]) ? node10116 : 4'b1000;
															assign node10116 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node10119 = (inp[11]) ? 4'b0000 : node10120;
														assign node10120 = (inp[12]) ? node10122 : 4'b0001;
															assign node10122 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node10126 = (inp[13]) ? node10128 : 4'b0110;
											assign node10128 = (inp[4]) ? node10130 : 4'b0110;
												assign node10130 = (inp[10]) ? node10132 : 4'b0110;
													assign node10132 = (inp[12]) ? node10134 : 4'b0000;
														assign node10134 = (inp[11]) ? 4'b0000 : 4'b0110;
									assign node10137 = (inp[4]) ? node10175 : node10138;
										assign node10138 = (inp[1]) ? node10156 : node10139;
											assign node10139 = (inp[13]) ? node10149 : node10140;
												assign node10140 = (inp[10]) ? node10142 : 4'b0101;
													assign node10142 = (inp[12]) ? node10146 : node10143;
														assign node10143 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node10146 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node10149 = (inp[11]) ? 4'b1101 : node10150;
													assign node10150 = (inp[7]) ? node10152 : 4'b1101;
														assign node10152 = (inp[10]) ? 4'b0100 : 4'b1100;
											assign node10156 = (inp[14]) ? node10164 : node10157;
												assign node10157 = (inp[13]) ? node10159 : 4'b1100;
													assign node10159 = (inp[7]) ? 4'b0100 : node10160;
														assign node10160 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node10164 = (inp[11]) ? node10168 : node10165;
													assign node10165 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node10168 = (inp[7]) ? 4'b0100 : node10169;
														assign node10169 = (inp[10]) ? 4'b1100 : node10170;
															assign node10170 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node10175 = (inp[7]) ? node10205 : node10176;
											assign node10176 = (inp[1]) ? node10192 : node10177;
												assign node10177 = (inp[13]) ? node10187 : node10178;
													assign node10178 = (inp[11]) ? node10182 : node10179;
														assign node10179 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10182 = (inp[10]) ? node10184 : 4'b0001;
															assign node10184 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10187 = (inp[14]) ? node10189 : 4'b1001;
														assign node10189 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node10192 = (inp[14]) ? node10196 : node10193;
													assign node10193 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node10196 = (inp[11]) ? 4'b1000 : node10197;
														assign node10197 = (inp[12]) ? 4'b1001 : node10198;
															assign node10198 = (inp[13]) ? 4'b0001 : node10199;
																assign node10199 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node10205 = (inp[1]) ? node10215 : node10206;
												assign node10206 = (inp[14]) ? node10208 : 4'b1101;
													assign node10208 = (inp[11]) ? node10212 : node10209;
														assign node10209 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node10212 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node10215 = (inp[13]) ? node10223 : node10216;
													assign node10216 = (inp[11]) ? 4'b0100 : node10217;
														assign node10217 = (inp[14]) ? node10219 : 4'b1100;
															assign node10219 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node10223 = (inp[10]) ? 4'b0000 : node10224;
														assign node10224 = (inp[12]) ? 4'b1100 : 4'b0000;
								assign node10228 = (inp[4]) ? node10300 : node10229;
									assign node10229 = (inp[1]) ? node10265 : node10230;
										assign node10230 = (inp[14]) ? node10244 : node10231;
											assign node10231 = (inp[13]) ? node10237 : node10232;
												assign node10232 = (inp[10]) ? node10234 : 4'b0001;
													assign node10234 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node10237 = (inp[12]) ? 4'b1001 : node10238;
													assign node10238 = (inp[10]) ? node10240 : 4'b1001;
														assign node10240 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node10244 = (inp[11]) ? node10254 : node10245;
												assign node10245 = (inp[12]) ? node10251 : node10246;
													assign node10246 = (inp[10]) ? 4'b0100 : node10247;
														assign node10247 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node10251 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node10254 = (inp[10]) ? node10258 : node10255;
													assign node10255 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node10258 = (inp[12]) ? 4'b1001 : node10259;
														assign node10259 = (inp[13]) ? node10261 : 4'b1001;
															assign node10261 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node10265 = (inp[11]) ? node10283 : node10266;
											assign node10266 = (inp[14]) ? node10276 : node10267;
												assign node10267 = (inp[10]) ? 4'b1000 : node10268;
													assign node10268 = (inp[7]) ? node10270 : 4'b1000;
														assign node10270 = (inp[5]) ? 4'b0000 : node10271;
															assign node10271 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node10276 = (inp[13]) ? node10278 : 4'b0001;
													assign node10278 = (inp[10]) ? node10280 : 4'b1001;
														assign node10280 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node10283 = (inp[13]) ? node10291 : node10284;
												assign node10284 = (inp[7]) ? node10286 : 4'b1000;
													assign node10286 = (inp[12]) ? node10288 : 4'b1000;
														assign node10288 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node10291 = (inp[12]) ? node10295 : node10292;
													assign node10292 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node10295 = (inp[10]) ? node10297 : 4'b1000;
														assign node10297 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node10300 = (inp[7]) ? node10346 : node10301;
										assign node10301 = (inp[1]) ? node10323 : node10302;
											assign node10302 = (inp[14]) ? node10310 : node10303;
												assign node10303 = (inp[10]) ? node10305 : 4'b1101;
													assign node10305 = (inp[13]) ? node10307 : 4'b1101;
														assign node10307 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node10310 = (inp[11]) ? node10316 : node10311;
													assign node10311 = (inp[13]) ? 4'b0100 : node10312;
														assign node10312 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node10316 = (inp[5]) ? node10318 : 4'b1101;
														assign node10318 = (inp[12]) ? node10320 : 4'b0101;
															assign node10320 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node10323 = (inp[14]) ? node10333 : node10324;
												assign node10324 = (inp[13]) ? node10330 : node10325;
													assign node10325 = (inp[12]) ? node10327 : 4'b1100;
														assign node10327 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node10330 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node10333 = (inp[11]) ? node10337 : node10334;
													assign node10334 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node10337 = (inp[5]) ? 4'b1100 : node10338;
														assign node10338 = (inp[12]) ? node10340 : 4'b1100;
															assign node10340 = (inp[13]) ? 4'b0100 : node10341;
																assign node10341 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node10346 = (inp[13]) ? node10372 : node10347;
											assign node10347 = (inp[14]) ? node10355 : node10348;
												assign node10348 = (inp[1]) ? node10350 : 4'b0001;
													assign node10350 = (inp[10]) ? 4'b1000 : node10351;
														assign node10351 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10355 = (inp[12]) ? node10365 : node10356;
													assign node10356 = (inp[10]) ? node10362 : node10357;
														assign node10357 = (inp[1]) ? 4'b1000 : node10358;
															assign node10358 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node10362 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node10365 = (inp[10]) ? 4'b0001 : node10366;
														assign node10366 = (inp[1]) ? node10368 : 4'b0000;
															assign node10368 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node10372 = (inp[1]) ? node10380 : node10373;
												assign node10373 = (inp[14]) ? 4'b1000 : node10374;
													assign node10374 = (inp[10]) ? node10376 : 4'b1001;
														assign node10376 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node10380 = (inp[11]) ? 4'b0100 : 4'b1001;
							assign node10383 = (inp[5]) ? node10385 : 4'b0110;
								assign node10385 = (inp[3]) ? node10447 : node10386;
									assign node10386 = (inp[4]) ? node10408 : node10387;
										assign node10387 = (inp[13]) ? node10389 : 4'b0110;
											assign node10389 = (inp[12]) ? node10399 : node10390;
												assign node10390 = (inp[7]) ? 4'b0110 : node10391;
													assign node10391 = (inp[10]) ? node10395 : node10392;
														assign node10392 = (inp[1]) ? 4'b0000 : 4'b0110;
														assign node10395 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node10399 = (inp[10]) ? node10401 : 4'b0110;
													assign node10401 = (inp[1]) ? node10403 : 4'b0110;
														assign node10403 = (inp[7]) ? 4'b0110 : node10404;
															assign node10404 = (inp[14]) ? 4'b0110 : 4'b0000;
										assign node10408 = (inp[7]) ? node10436 : node10409;
											assign node10409 = (inp[13]) ? node10423 : node10410;
												assign node10410 = (inp[14]) ? node10418 : node10411;
													assign node10411 = (inp[1]) ? 4'b1000 : node10412;
														assign node10412 = (inp[10]) ? node10414 : 4'b0001;
															assign node10414 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10418 = (inp[1]) ? 4'b0001 : node10419;
														assign node10419 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node10423 = (inp[10]) ? node10433 : node10424;
													assign node10424 = (inp[11]) ? node10430 : node10425;
														assign node10425 = (inp[1]) ? 4'b1001 : node10426;
															assign node10426 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10430 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node10433 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node10436 = (inp[13]) ? node10438 : 4'b0110;
												assign node10438 = (inp[10]) ? node10440 : 4'b0110;
													assign node10440 = (inp[11]) ? node10444 : node10441;
														assign node10441 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node10444 = (inp[1]) ? 4'b0000 : 4'b0110;
									assign node10447 = (inp[1]) ? node10487 : node10448;
										assign node10448 = (inp[13]) ? node10464 : node10449;
											assign node10449 = (inp[14]) ? node10459 : node10450;
												assign node10450 = (inp[7]) ? node10454 : node10451;
													assign node10451 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node10454 = (inp[12]) ? 4'b0001 : node10455;
														assign node10455 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node10459 = (inp[11]) ? 4'b0001 : node10460;
													assign node10460 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node10464 = (inp[10]) ? node10472 : node10465;
												assign node10465 = (inp[12]) ? node10467 : 4'b1001;
													assign node10467 = (inp[7]) ? 4'b1001 : node10468;
														assign node10468 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node10472 = (inp[12]) ? node10482 : node10473;
													assign node10473 = (inp[11]) ? node10479 : node10474;
														assign node10474 = (inp[14]) ? node10476 : 4'b0101;
															assign node10476 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10479 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node10482 = (inp[14]) ? node10484 : 4'b1001;
														assign node10484 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node10487 = (inp[4]) ? node10515 : node10488;
											assign node10488 = (inp[11]) ? node10502 : node10489;
												assign node10489 = (inp[14]) ? node10495 : node10490;
													assign node10490 = (inp[13]) ? 4'b0000 : node10491;
														assign node10491 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node10495 = (inp[12]) ? 4'b1001 : node10496;
														assign node10496 = (inp[10]) ? node10498 : 4'b0001;
															assign node10498 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node10502 = (inp[13]) ? node10508 : node10503;
													assign node10503 = (inp[10]) ? 4'b1000 : node10504;
														assign node10504 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10508 = (inp[12]) ? node10512 : node10509;
														assign node10509 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10512 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node10515 = (inp[7]) ? node10523 : node10516;
												assign node10516 = (inp[13]) ? node10518 : 4'b1100;
													assign node10518 = (inp[11]) ? node10520 : 4'b0100;
														assign node10520 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node10523 = (inp[11]) ? 4'b0100 : node10524;
													assign node10524 = (inp[14]) ? 4'b1001 : 4'b1000;
					assign node10529 = (inp[5]) ? node11131 : node10530;
						assign node10530 = (inp[0]) ? node10984 : node10531;
							assign node10531 = (inp[11]) ? node10789 : node10532;
								assign node10532 = (inp[3]) ? node10674 : node10533;
									assign node10533 = (inp[4]) ? node10619 : node10534;
										assign node10534 = (inp[13]) ? node10574 : node10535;
											assign node10535 = (inp[10]) ? node10551 : node10536;
												assign node10536 = (inp[2]) ? node10546 : node10537;
													assign node10537 = (inp[14]) ? node10543 : node10538;
														assign node10538 = (inp[1]) ? node10540 : 4'b0101;
															assign node10540 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10543 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node10546 = (inp[14]) ? node10548 : 4'b0101;
														assign node10548 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node10551 = (inp[7]) ? node10563 : node10552;
													assign node10552 = (inp[1]) ? node10558 : node10553;
														assign node10553 = (inp[14]) ? 4'b1100 : node10554;
															assign node10554 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10558 = (inp[12]) ? node10560 : 4'b0001;
															assign node10560 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node10563 = (inp[12]) ? node10569 : node10564;
														assign node10564 = (inp[14]) ? 4'b1100 : node10565;
															assign node10565 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node10569 = (inp[14]) ? node10571 : 4'b1100;
															assign node10571 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node10574 = (inp[10]) ? node10602 : node10575;
												assign node10575 = (inp[2]) ? node10589 : node10576;
													assign node10576 = (inp[7]) ? node10582 : node10577;
														assign node10577 = (inp[12]) ? 4'b0001 : node10578;
															assign node10578 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node10582 = (inp[14]) ? node10586 : node10583;
															assign node10583 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node10586 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node10589 = (inp[12]) ? node10593 : node10590;
														assign node10590 = (inp[14]) ? 4'b1100 : 4'b0100;
														assign node10593 = (inp[7]) ? 4'b1101 : node10594;
															assign node10594 = (inp[1]) ? node10598 : node10595;
																assign node10595 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node10598 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node10602 = (inp[12]) ? node10614 : node10603;
													assign node10603 = (inp[7]) ? node10611 : node10604;
														assign node10604 = (inp[14]) ? node10608 : node10605;
															assign node10605 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node10608 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node10611 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node10614 = (inp[7]) ? 4'b0100 : node10615;
														assign node10615 = (inp[2]) ? 4'b1101 : 4'b1001;
										assign node10619 = (inp[2]) ? node10635 : node10620;
											assign node10620 = (inp[10]) ? node10630 : node10621;
												assign node10621 = (inp[13]) ? node10627 : node10622;
													assign node10622 = (inp[1]) ? node10624 : 4'b0001;
														assign node10624 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10627 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node10630 = (inp[7]) ? 4'b1001 : node10631;
													assign node10631 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node10635 = (inp[7]) ? node10653 : node10636;
												assign node10636 = (inp[13]) ? node10644 : node10637;
													assign node10637 = (inp[12]) ? node10639 : 4'b1000;
														assign node10639 = (inp[1]) ? 4'b1000 : node10640;
															assign node10640 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10644 = (inp[12]) ? node10650 : node10645;
														assign node10645 = (inp[14]) ? node10647 : 4'b0000;
															assign node10647 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node10650 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node10653 = (inp[10]) ? node10665 : node10654;
													assign node10654 = (inp[13]) ? node10660 : node10655;
														assign node10655 = (inp[1]) ? node10657 : 4'b0101;
															assign node10657 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10660 = (inp[14]) ? node10662 : 4'b1101;
															assign node10662 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node10665 = (inp[13]) ? node10669 : node10666;
														assign node10666 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node10669 = (inp[14]) ? node10671 : 4'b0000;
															assign node10671 = (inp[12]) ? 4'b1100 : 4'b0000;
									assign node10674 = (inp[10]) ? node10718 : node10675;
										assign node10675 = (inp[2]) ? node10699 : node10676;
											assign node10676 = (inp[4]) ? node10684 : node10677;
												assign node10677 = (inp[13]) ? node10681 : node10678;
													assign node10678 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node10681 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node10684 = (inp[7]) ? node10692 : node10685;
													assign node10685 = (inp[13]) ? node10689 : node10686;
														assign node10686 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node10689 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node10692 = (inp[13]) ? node10694 : 4'b0001;
														assign node10694 = (inp[1]) ? 4'b0001 : node10695;
															assign node10695 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node10699 = (inp[4]) ? node10707 : node10700;
												assign node10700 = (inp[7]) ? node10702 : 4'b0001;
													assign node10702 = (inp[1]) ? node10704 : 4'b1000;
														assign node10704 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node10707 = (inp[7]) ? 4'b0001 : node10708;
													assign node10708 = (inp[13]) ? node10714 : node10709;
														assign node10709 = (inp[14]) ? 4'b0001 : node10710;
															assign node10710 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10714 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node10718 = (inp[7]) ? node10754 : node10719;
											assign node10719 = (inp[13]) ? node10739 : node10720;
												assign node10720 = (inp[12]) ? node10730 : node10721;
													assign node10721 = (inp[2]) ? 4'b0101 : node10722;
														assign node10722 = (inp[14]) ? node10724 : 4'b1001;
															assign node10724 = (inp[1]) ? 4'b0001 : node10725;
																assign node10725 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node10730 = (inp[14]) ? node10736 : node10731;
														assign node10731 = (inp[4]) ? 4'b0001 : node10732;
															assign node10732 = (inp[2]) ? 4'b1000 : 4'b1101;
														assign node10736 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node10739 = (inp[4]) ? node10743 : node10740;
													assign node10740 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node10743 = (inp[2]) ? node10749 : node10744;
														assign node10744 = (inp[14]) ? node10746 : 4'b1100;
															assign node10746 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node10749 = (inp[1]) ? node10751 : 4'b1101;
															assign node10751 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node10754 = (inp[12]) ? node10772 : node10755;
												assign node10755 = (inp[14]) ? node10763 : node10756;
													assign node10756 = (inp[13]) ? node10760 : node10757;
														assign node10757 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node10760 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node10763 = (inp[4]) ? node10769 : node10764;
														assign node10764 = (inp[2]) ? node10766 : 4'b1101;
															assign node10766 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node10769 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node10772 = (inp[1]) ? node10774 : 4'b1001;
													assign node10774 = (inp[13]) ? node10780 : node10775;
														assign node10775 = (inp[2]) ? node10777 : 4'b0000;
															assign node10777 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node10780 = (inp[14]) ? node10784 : node10781;
															assign node10781 = (inp[2]) ? 4'b0000 : 4'b1001;
															assign node10784 = (inp[4]) ? 4'b1000 : node10785;
																assign node10785 = (inp[2]) ? 4'b1001 : 4'b1101;
								assign node10789 = (inp[1]) ? node10913 : node10790;
									assign node10790 = (inp[3]) ? node10840 : node10791;
										assign node10791 = (inp[2]) ? node10815 : node10792;
											assign node10792 = (inp[4]) ? node10810 : node10793;
												assign node10793 = (inp[13]) ? node10803 : node10794;
													assign node10794 = (inp[10]) ? node10796 : 4'b0101;
														assign node10796 = (inp[7]) ? node10800 : node10797;
															assign node10797 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node10800 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node10803 = (inp[10]) ? node10805 : 4'b1101;
														assign node10805 = (inp[12]) ? node10807 : 4'b0000;
															assign node10807 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node10810 = (inp[13]) ? 4'b0100 : node10811;
													assign node10811 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node10815 = (inp[7]) ? node10829 : node10816;
												assign node10816 = (inp[4]) ? node10822 : node10817;
													assign node10817 = (inp[14]) ? node10819 : 4'b1101;
														assign node10819 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node10822 = (inp[10]) ? node10824 : 4'b0001;
														assign node10824 = (inp[13]) ? node10826 : 4'b1001;
															assign node10826 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node10829 = (inp[10]) ? node10833 : node10830;
													assign node10830 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node10833 = (inp[13]) ? node10837 : node10834;
														assign node10834 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10837 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node10840 = (inp[2]) ? node10880 : node10841;
											assign node10841 = (inp[4]) ? node10861 : node10842;
												assign node10842 = (inp[7]) ? node10854 : node10843;
													assign node10843 = (inp[13]) ? 4'b1000 : node10844;
														assign node10844 = (inp[14]) ? node10848 : node10845;
															assign node10845 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node10848 = (inp[12]) ? node10850 : 4'b1100;
																assign node10850 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node10854 = (inp[12]) ? node10858 : node10855;
														assign node10855 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node10858 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node10861 = (inp[13]) ? node10871 : node10862;
													assign node10862 = (inp[10]) ? 4'b0001 : node10863;
														assign node10863 = (inp[7]) ? node10867 : node10864;
															assign node10864 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10867 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10871 = (inp[7]) ? node10875 : node10872;
														assign node10872 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node10875 = (inp[10]) ? 4'b1001 : node10876;
															assign node10876 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node10880 = (inp[4]) ? node10902 : node10881;
												assign node10881 = (inp[7]) ? node10895 : node10882;
													assign node10882 = (inp[13]) ? node10886 : node10883;
														assign node10883 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node10886 = (inp[14]) ? node10888 : 4'b0000;
															assign node10888 = (inp[12]) ? node10892 : node10889;
																assign node10889 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node10892 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node10895 = (inp[13]) ? node10897 : 4'b0001;
														assign node10897 = (inp[10]) ? node10899 : 4'b1001;
															assign node10899 = (inp[14]) ? 4'b0000 : 4'b1001;
												assign node10902 = (inp[7]) ? node10908 : node10903;
													assign node10903 = (inp[13]) ? node10905 : 4'b1000;
														assign node10905 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node10908 = (inp[10]) ? node10910 : 4'b0000;
														assign node10910 = (inp[14]) ? 4'b0000 : 4'b1000;
									assign node10913 = (inp[10]) ? node10951 : node10914;
										assign node10914 = (inp[2]) ? node10932 : node10915;
											assign node10915 = (inp[4]) ? node10923 : node10916;
												assign node10916 = (inp[7]) ? node10918 : 4'b1000;
													assign node10918 = (inp[3]) ? 4'b1100 : node10919;
														assign node10919 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node10923 = (inp[13]) ? node10929 : node10924;
													assign node10924 = (inp[7]) ? node10926 : 4'b1000;
														assign node10926 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node10929 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node10932 = (inp[3]) ? node10940 : node10933;
												assign node10933 = (inp[14]) ? node10935 : 4'b0100;
													assign node10935 = (inp[13]) ? 4'b0000 : node10936;
														assign node10936 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node10940 = (inp[4]) ? node10948 : node10941;
													assign node10941 = (inp[7]) ? node10943 : 4'b0000;
														assign node10943 = (inp[14]) ? 4'b1000 : node10944;
															assign node10944 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node10948 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node10951 = (inp[13]) ? node10973 : node10952;
											assign node10952 = (inp[4]) ? node10964 : node10953;
												assign node10953 = (inp[3]) ? node10959 : node10954;
													assign node10954 = (inp[2]) ? 4'b1100 : node10955;
														assign node10955 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node10959 = (inp[2]) ? node10961 : 4'b0100;
														assign node10961 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node10964 = (inp[7]) ? node10966 : 4'b1000;
													assign node10966 = (inp[14]) ? node10968 : 4'b0000;
														assign node10968 = (inp[2]) ? node10970 : 4'b0000;
															assign node10970 = (inp[3]) ? 4'b0000 : 4'b1100;
											assign node10973 = (inp[4]) ? node10979 : node10974;
												assign node10974 = (inp[7]) ? node10976 : 4'b0000;
													assign node10976 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node10979 = (inp[3]) ? 4'b0100 : node10980;
													assign node10980 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node10984 = (inp[2]) ? 4'b0100 : node10985;
								assign node10985 = (inp[3]) ? node11033 : node10986;
									assign node10986 = (inp[4]) ? node10996 : node10987;
										assign node10987 = (inp[10]) ? node10989 : 4'b0100;
											assign node10989 = (inp[12]) ? 4'b0100 : node10990;
												assign node10990 = (inp[14]) ? 4'b0100 : node10991;
													assign node10991 = (inp[1]) ? 4'b0100 : 4'b0001;
										assign node10996 = (inp[7]) ? node11024 : node10997;
											assign node10997 = (inp[12]) ? node11017 : node10998;
												assign node10998 = (inp[1]) ? node11008 : node10999;
													assign node10999 = (inp[11]) ? node11003 : node11000;
														assign node11000 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11003 = (inp[10]) ? node11005 : 4'b1001;
															assign node11005 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node11008 = (inp[11]) ? 4'b1000 : node11009;
														assign node11009 = (inp[14]) ? node11011 : 4'b1000;
															assign node11011 = (inp[13]) ? 4'b1001 : node11012;
																assign node11012 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node11017 = (inp[10]) ? node11019 : 4'b0000;
													assign node11019 = (inp[14]) ? 4'b1000 : node11020;
														assign node11020 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node11024 = (inp[13]) ? node11026 : 4'b0100;
												assign node11026 = (inp[11]) ? node11028 : 4'b0000;
													assign node11028 = (inp[12]) ? 4'b0100 : node11029;
														assign node11029 = (inp[10]) ? 4'b0001 : 4'b0100;
									assign node11033 = (inp[4]) ? node11085 : node11034;
										assign node11034 = (inp[1]) ? node11058 : node11035;
											assign node11035 = (inp[14]) ? node11047 : node11036;
												assign node11036 = (inp[7]) ? node11042 : node11037;
													assign node11037 = (inp[10]) ? 4'b0101 : node11038;
														assign node11038 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node11042 = (inp[10]) ? 4'b1001 : node11043;
														assign node11043 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node11047 = (inp[11]) ? node11055 : node11048;
													assign node11048 = (inp[7]) ? node11050 : 4'b1000;
														assign node11050 = (inp[13]) ? node11052 : 4'b0000;
															assign node11052 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node11055 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node11058 = (inp[11]) ? node11074 : node11059;
												assign node11059 = (inp[14]) ? node11063 : node11060;
													assign node11060 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node11063 = (inp[10]) ? node11067 : node11064;
														assign node11064 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node11067 = (inp[13]) ? node11071 : node11068;
															assign node11068 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11071 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node11074 = (inp[12]) ? node11078 : node11075;
													assign node11075 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node11078 = (inp[10]) ? node11082 : node11079;
														assign node11079 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node11082 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node11085 = (inp[7]) ? node11105 : node11086;
											assign node11086 = (inp[1]) ? node11096 : node11087;
												assign node11087 = (inp[13]) ? node11093 : node11088;
													assign node11088 = (inp[12]) ? 4'b0101 : node11089;
														assign node11089 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node11093 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node11096 = (inp[13]) ? node11102 : node11097;
													assign node11097 = (inp[11]) ? 4'b1100 : node11098;
														assign node11098 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node11102 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node11105 = (inp[10]) ? node11121 : node11106;
												assign node11106 = (inp[11]) ? node11114 : node11107;
													assign node11107 = (inp[13]) ? node11109 : 4'b0000;
														assign node11109 = (inp[14]) ? 4'b1001 : node11110;
															assign node11110 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node11114 = (inp[14]) ? node11118 : node11115;
														assign node11115 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node11118 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node11121 = (inp[13]) ? node11125 : node11122;
													assign node11122 = (inp[12]) ? 4'b0001 : 4'b1000;
													assign node11125 = (inp[1]) ? 4'b0100 : node11126;
														assign node11126 = (inp[11]) ? 4'b0101 : 4'b1001;
						assign node11131 = (inp[3]) ? node11495 : node11132;
							assign node11132 = (inp[4]) ? node11306 : node11133;
								assign node11133 = (inp[13]) ? node11205 : node11134;
									assign node11134 = (inp[0]) ? node11180 : node11135;
										assign node11135 = (inp[7]) ? node11159 : node11136;
											assign node11136 = (inp[10]) ? node11152 : node11137;
												assign node11137 = (inp[12]) ? node11145 : node11138;
													assign node11138 = (inp[1]) ? node11140 : 4'b1100;
														assign node11140 = (inp[2]) ? node11142 : 4'b0000;
															assign node11142 = (inp[11]) ? 4'b0000 : 4'b1101;
													assign node11145 = (inp[11]) ? 4'b0100 : node11146;
														assign node11146 = (inp[14]) ? node11148 : 4'b0101;
															assign node11148 = (inp[1]) ? 4'b1100 : 4'b0101;
												assign node11152 = (inp[2]) ? node11154 : 4'b0000;
													assign node11154 = (inp[1]) ? node11156 : 4'b0001;
														assign node11156 = (inp[12]) ? 4'b1000 : 4'b1001;
											assign node11159 = (inp[11]) ? node11167 : node11160;
												assign node11160 = (inp[14]) ? node11162 : 4'b0101;
													assign node11162 = (inp[10]) ? node11164 : 4'b0101;
														assign node11164 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node11167 = (inp[10]) ? node11171 : node11168;
													assign node11168 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node11171 = (inp[2]) ? node11175 : node11172;
														assign node11172 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node11175 = (inp[1]) ? 4'b0100 : node11176;
															assign node11176 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node11180 = (inp[2]) ? 4'b0100 : node11181;
											assign node11181 = (inp[1]) ? node11193 : node11182;
												assign node11182 = (inp[14]) ? node11188 : node11183;
													assign node11183 = (inp[12]) ? 4'b0101 : node11184;
														assign node11184 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node11188 = (inp[11]) ? node11190 : 4'b0100;
														assign node11190 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node11193 = (inp[11]) ? node11199 : node11194;
													assign node11194 = (inp[10]) ? 4'b0001 : node11195;
														assign node11195 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node11199 = (inp[12]) ? node11201 : 4'b1100;
														assign node11201 = (inp[10]) ? 4'b1100 : 4'b0100;
									assign node11205 = (inp[1]) ? node11255 : node11206;
										assign node11206 = (inp[0]) ? node11232 : node11207;
											assign node11207 = (inp[2]) ? node11219 : node11208;
												assign node11208 = (inp[10]) ? node11216 : node11209;
													assign node11209 = (inp[7]) ? node11211 : 4'b0000;
														assign node11211 = (inp[12]) ? node11213 : 4'b1000;
															assign node11213 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node11216 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node11219 = (inp[7]) ? node11227 : node11220;
													assign node11220 = (inp[11]) ? 4'b1001 : node11221;
														assign node11221 = (inp[14]) ? node11223 : 4'b1000;
															assign node11223 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node11227 = (inp[10]) ? 4'b1001 : node11228;
														assign node11228 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node11232 = (inp[2]) ? node11248 : node11233;
												assign node11233 = (inp[11]) ? node11243 : node11234;
													assign node11234 = (inp[7]) ? node11238 : node11235;
														assign node11235 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11238 = (inp[12]) ? node11240 : 4'b0101;
															assign node11240 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node11243 = (inp[12]) ? 4'b0000 : node11244;
														assign node11244 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node11248 = (inp[14]) ? node11250 : 4'b0100;
													assign node11250 = (inp[10]) ? node11252 : 4'b0100;
														assign node11252 = (inp[11]) ? 4'b0100 : 4'b0000;
										assign node11255 = (inp[11]) ? node11281 : node11256;
											assign node11256 = (inp[10]) ? node11264 : node11257;
												assign node11257 = (inp[14]) ? node11259 : 4'b0001;
													assign node11259 = (inp[12]) ? node11261 : 4'b1101;
														assign node11261 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node11264 = (inp[2]) ? node11272 : node11265;
													assign node11265 = (inp[0]) ? 4'b0001 : node11266;
														assign node11266 = (inp[12]) ? 4'b1000 : node11267;
															assign node11267 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node11272 = (inp[14]) ? node11276 : node11273;
														assign node11273 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node11276 = (inp[12]) ? 4'b0100 : node11277;
															assign node11277 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node11281 = (inp[10]) ? node11299 : node11282;
												assign node11282 = (inp[2]) ? node11292 : node11283;
													assign node11283 = (inp[12]) ? node11285 : 4'b0100;
														assign node11285 = (inp[0]) ? node11289 : node11286;
															assign node11286 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node11289 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node11292 = (inp[7]) ? node11296 : node11293;
														assign node11293 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node11296 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11299 = (inp[7]) ? 4'b0100 : node11300;
													assign node11300 = (inp[14]) ? 4'b0000 : node11301;
														assign node11301 = (inp[12]) ? 4'b0100 : 4'b0000;
								assign node11306 = (inp[1]) ? node11430 : node11307;
									assign node11307 = (inp[7]) ? node11373 : node11308;
										assign node11308 = (inp[13]) ? node11334 : node11309;
											assign node11309 = (inp[12]) ? node11323 : node11310;
												assign node11310 = (inp[2]) ? node11320 : node11311;
													assign node11311 = (inp[11]) ? node11315 : node11312;
														assign node11312 = (inp[0]) ? 4'b0001 : 4'b1000;
														assign node11315 = (inp[10]) ? node11317 : 4'b1000;
															assign node11317 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node11320 = (inp[10]) ? 4'b1001 : 4'b0101;
												assign node11323 = (inp[0]) ? node11331 : node11324;
													assign node11324 = (inp[11]) ? 4'b1001 : node11325;
														assign node11325 = (inp[2]) ? 4'b0100 : node11326;
															assign node11326 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node11331 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node11334 = (inp[10]) ? node11352 : node11335;
												assign node11335 = (inp[2]) ? node11345 : node11336;
													assign node11336 = (inp[14]) ? node11340 : node11337;
														assign node11337 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node11340 = (inp[12]) ? 4'b0001 : node11341;
															assign node11341 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node11345 = (inp[0]) ? node11347 : 4'b1000;
														assign node11347 = (inp[14]) ? node11349 : 4'b1001;
															assign node11349 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node11352 = (inp[0]) ? node11358 : node11353;
													assign node11353 = (inp[14]) ? node11355 : 4'b0001;
														assign node11355 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node11358 = (inp[11]) ? node11368 : node11359;
														assign node11359 = (inp[12]) ? node11363 : node11360;
															assign node11360 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node11363 = (inp[2]) ? node11365 : 4'b0001;
																assign node11365 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11368 = (inp[2]) ? node11370 : 4'b1001;
															assign node11370 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node11373 = (inp[13]) ? node11399 : node11374;
											assign node11374 = (inp[2]) ? node11388 : node11375;
												assign node11375 = (inp[11]) ? node11379 : node11376;
													assign node11376 = (inp[0]) ? 4'b0001 : 4'b0100;
													assign node11379 = (inp[10]) ? node11383 : node11380;
														assign node11380 = (inp[0]) ? 4'b1000 : 4'b1100;
														assign node11383 = (inp[12]) ? node11385 : 4'b0001;
															assign node11385 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node11388 = (inp[14]) ? node11392 : node11389;
													assign node11389 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node11392 = (inp[0]) ? 4'b0100 : node11393;
														assign node11393 = (inp[12]) ? node11395 : 4'b0101;
															assign node11395 = (inp[11]) ? 4'b0101 : 4'b1001;
											assign node11399 = (inp[0]) ? node11415 : node11400;
												assign node11400 = (inp[2]) ? node11410 : node11401;
													assign node11401 = (inp[11]) ? node11405 : node11402;
														assign node11402 = (inp[14]) ? 4'b1000 : 4'b0101;
														assign node11405 = (inp[14]) ? 4'b0000 : node11406;
															assign node11406 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11410 = (inp[11]) ? 4'b1000 : node11411;
														assign node11411 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11415 = (inp[2]) ? node11425 : node11416;
													assign node11416 = (inp[11]) ? node11420 : node11417;
														assign node11417 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11420 = (inp[10]) ? 4'b0100 : node11421;
															assign node11421 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11425 = (inp[10]) ? node11427 : 4'b0100;
														assign node11427 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node11430 = (inp[2]) ? node11472 : node11431;
										assign node11431 = (inp[11]) ? node11457 : node11432;
											assign node11432 = (inp[0]) ? node11442 : node11433;
												assign node11433 = (inp[14]) ? node11437 : node11434;
													assign node11434 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node11437 = (inp[12]) ? node11439 : 4'b0001;
														assign node11439 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node11442 = (inp[10]) ? node11448 : node11443;
													assign node11443 = (inp[12]) ? 4'b0001 : node11444;
														assign node11444 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node11448 = (inp[12]) ? node11452 : node11449;
														assign node11449 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11452 = (inp[13]) ? node11454 : 4'b1001;
															assign node11454 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node11457 = (inp[10]) ? node11465 : node11458;
												assign node11458 = (inp[12]) ? node11460 : 4'b1000;
													assign node11460 = (inp[13]) ? 4'b1000 : node11461;
														assign node11461 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node11465 = (inp[13]) ? 4'b0000 : node11466;
													assign node11466 = (inp[0]) ? node11468 : 4'b0000;
														assign node11468 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node11472 = (inp[0]) ? node11490 : node11473;
											assign node11473 = (inp[12]) ? node11483 : node11474;
												assign node11474 = (inp[7]) ? node11478 : node11475;
													assign node11475 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node11478 = (inp[13]) ? 4'b0000 : node11479;
														assign node11479 = (inp[14]) ? 4'b0000 : 4'b1001;
												assign node11483 = (inp[11]) ? node11485 : 4'b1000;
													assign node11485 = (inp[7]) ? node11487 : 4'b0000;
														assign node11487 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node11490 = (inp[7]) ? 4'b0100 : node11491;
												assign node11491 = (inp[11]) ? 4'b1000 : 4'b0000;
							assign node11495 = (inp[4]) ? node11701 : node11496;
								assign node11496 = (inp[11]) ? node11620 : node11497;
									assign node11497 = (inp[13]) ? node11549 : node11498;
										assign node11498 = (inp[14]) ? node11528 : node11499;
											assign node11499 = (inp[0]) ? node11517 : node11500;
												assign node11500 = (inp[1]) ? node11508 : node11501;
													assign node11501 = (inp[2]) ? node11503 : 4'b1000;
														assign node11503 = (inp[12]) ? 4'b1001 : node11504;
															assign node11504 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node11508 = (inp[7]) ? node11512 : node11509;
														assign node11509 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node11512 = (inp[10]) ? 4'b0000 : node11513;
															assign node11513 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node11517 = (inp[10]) ? 4'b1000 : node11518;
													assign node11518 = (inp[12]) ? 4'b0000 : node11519;
														assign node11519 = (inp[7]) ? node11523 : node11520;
															assign node11520 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node11523 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node11528 = (inp[1]) ? node11536 : node11529;
												assign node11529 = (inp[2]) ? 4'b0000 : node11530;
													assign node11530 = (inp[10]) ? node11532 : 4'b0001;
														assign node11532 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node11536 = (inp[0]) ? 4'b0001 : node11537;
													assign node11537 = (inp[12]) ? node11543 : node11538;
														assign node11538 = (inp[7]) ? node11540 : 4'b0001;
															assign node11540 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11543 = (inp[2]) ? 4'b1001 : node11544;
															assign node11544 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node11549 = (inp[7]) ? node11579 : node11550;
											assign node11550 = (inp[2]) ? node11560 : node11551;
												assign node11551 = (inp[1]) ? node11553 : 4'b0001;
													assign node11553 = (inp[10]) ? node11557 : node11554;
														assign node11554 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node11557 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node11560 = (inp[12]) ? node11574 : node11561;
													assign node11561 = (inp[10]) ? node11565 : node11562;
														assign node11562 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node11565 = (inp[14]) ? node11569 : node11566;
															assign node11566 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node11569 = (inp[0]) ? 4'b0000 : node11570;
																assign node11570 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node11574 = (inp[10]) ? 4'b0001 : node11575;
														assign node11575 = (inp[0]) ? 4'b0001 : 4'b1000;
											assign node11579 = (inp[10]) ? node11599 : node11580;
												assign node11580 = (inp[0]) ? node11590 : node11581;
													assign node11581 = (inp[12]) ? node11583 : 4'b0001;
														assign node11583 = (inp[1]) ? node11587 : node11584;
															assign node11584 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node11587 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node11590 = (inp[2]) ? node11594 : node11591;
														assign node11591 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node11594 = (inp[14]) ? 4'b1001 : node11595;
															assign node11595 = (inp[12]) ? 4'b1000 : 4'b1001;
												assign node11599 = (inp[2]) ? node11613 : node11600;
													assign node11600 = (inp[1]) ? node11606 : node11601;
														assign node11601 = (inp[0]) ? node11603 : 4'b0000;
															assign node11603 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11606 = (inp[14]) ? 4'b0001 : node11607;
															assign node11607 = (inp[0]) ? node11609 : 4'b1000;
																assign node11609 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node11613 = (inp[1]) ? node11615 : 4'b1000;
														assign node11615 = (inp[14]) ? 4'b0001 : node11616;
															assign node11616 = (inp[0]) ? 4'b0000 : 4'b1000;
									assign node11620 = (inp[1]) ? node11666 : node11621;
										assign node11621 = (inp[12]) ? node11645 : node11622;
											assign node11622 = (inp[10]) ? node11632 : node11623;
												assign node11623 = (inp[7]) ? node11627 : node11624;
													assign node11624 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node11627 = (inp[2]) ? node11629 : 4'b1000;
														assign node11629 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node11632 = (inp[2]) ? node11642 : node11633;
													assign node11633 = (inp[7]) ? node11637 : node11634;
														assign node11634 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node11637 = (inp[0]) ? node11639 : 4'b0000;
															assign node11639 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node11642 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node11645 = (inp[13]) ? node11653 : node11646;
												assign node11646 = (inp[0]) ? 4'b0001 : node11647;
													assign node11647 = (inp[10]) ? node11649 : 4'b1001;
														assign node11649 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node11653 = (inp[14]) ? node11659 : node11654;
													assign node11654 = (inp[7]) ? node11656 : 4'b1001;
														assign node11656 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node11659 = (inp[10]) ? node11663 : node11660;
														assign node11660 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node11663 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node11666 = (inp[2]) ? node11684 : node11667;
											assign node11667 = (inp[7]) ? node11669 : 4'b0000;
												assign node11669 = (inp[14]) ? node11675 : node11670;
													assign node11670 = (inp[0]) ? node11672 : 4'b0000;
														assign node11672 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node11675 = (inp[0]) ? 4'b0000 : node11676;
														assign node11676 = (inp[13]) ? node11680 : node11677;
															assign node11677 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node11680 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node11684 = (inp[13]) ? node11696 : node11685;
												assign node11685 = (inp[0]) ? node11689 : node11686;
													assign node11686 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node11689 = (inp[7]) ? 4'b1000 : node11690;
														assign node11690 = (inp[10]) ? 4'b0000 : node11691;
															assign node11691 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11696 = (inp[10]) ? 4'b0000 : node11697;
													assign node11697 = (inp[0]) ? 4'b1000 : 4'b0000;
								assign node11701 = (inp[13]) ? node11801 : node11702;
									assign node11702 = (inp[10]) ? node11760 : node11703;
										assign node11703 = (inp[1]) ? node11729 : node11704;
											assign node11704 = (inp[2]) ? node11718 : node11705;
												assign node11705 = (inp[0]) ? node11715 : node11706;
													assign node11706 = (inp[7]) ? node11710 : node11707;
														assign node11707 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node11710 = (inp[14]) ? node11712 : 4'b0000;
															assign node11712 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node11715 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node11718 = (inp[12]) ? node11722 : node11719;
													assign node11719 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node11722 = (inp[0]) ? node11726 : node11723;
														assign node11723 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node11726 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node11729 = (inp[11]) ? node11745 : node11730;
												assign node11730 = (inp[0]) ? node11736 : node11731;
													assign node11731 = (inp[7]) ? node11733 : 4'b0001;
														assign node11733 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11736 = (inp[2]) ? node11740 : node11737;
														assign node11737 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node11740 = (inp[12]) ? node11742 : 4'b1001;
															assign node11742 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node11745 = (inp[12]) ? node11747 : 4'b0000;
													assign node11747 = (inp[14]) ? node11753 : node11748;
														assign node11748 = (inp[7]) ? 4'b1000 : node11749;
															assign node11749 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node11753 = (inp[7]) ? 4'b0000 : node11754;
															assign node11754 = (inp[0]) ? 4'b0000 : node11755;
																assign node11755 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node11760 = (inp[12]) ? node11786 : node11761;
											assign node11761 = (inp[7]) ? node11771 : node11762;
												assign node11762 = (inp[0]) ? node11764 : 4'b0000;
													assign node11764 = (inp[2]) ? 4'b1000 : node11765;
														assign node11765 = (inp[14]) ? node11767 : 4'b0001;
															assign node11767 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node11771 = (inp[2]) ? node11777 : node11772;
													assign node11772 = (inp[0]) ? 4'b0000 : node11773;
														assign node11773 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node11777 = (inp[11]) ? node11783 : node11778;
														assign node11778 = (inp[0]) ? 4'b0000 : node11779;
															assign node11779 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node11783 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node11786 = (inp[7]) ? node11794 : node11787;
												assign node11787 = (inp[1]) ? node11789 : 4'b0000;
													assign node11789 = (inp[2]) ? node11791 : 4'b0000;
														assign node11791 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node11794 = (inp[11]) ? 4'b0000 : node11795;
													assign node11795 = (inp[2]) ? 4'b0001 : node11796;
														assign node11796 = (inp[0]) ? 4'b0001 : 4'b1000;
									assign node11801 = (inp[1]) ? node11851 : node11802;
										assign node11802 = (inp[10]) ? node11840 : node11803;
											assign node11803 = (inp[7]) ? node11821 : node11804;
												assign node11804 = (inp[11]) ? node11812 : node11805;
													assign node11805 = (inp[12]) ? node11807 : 4'b0000;
														assign node11807 = (inp[14]) ? node11809 : 4'b0001;
															assign node11809 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node11812 = (inp[12]) ? 4'b0000 : node11813;
														assign node11813 = (inp[14]) ? 4'b0001 : node11814;
															assign node11814 = (inp[2]) ? 4'b0000 : node11815;
																assign node11815 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node11821 = (inp[0]) ? node11829 : node11822;
													assign node11822 = (inp[11]) ? node11824 : 4'b0000;
														assign node11824 = (inp[12]) ? 4'b0001 : node11825;
															assign node11825 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node11829 = (inp[11]) ? node11835 : node11830;
														assign node11830 = (inp[2]) ? node11832 : 4'b0001;
															assign node11832 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11835 = (inp[12]) ? node11837 : 4'b0000;
															assign node11837 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node11840 = (inp[12]) ? node11842 : 4'b0000;
												assign node11842 = (inp[11]) ? 4'b0000 : node11843;
													assign node11843 = (inp[14]) ? node11845 : 4'b0001;
														assign node11845 = (inp[7]) ? 4'b0001 : node11846;
															assign node11846 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node11851 = (inp[7]) ? 4'b0000 : node11852;
											assign node11852 = (inp[11]) ? 4'b0000 : node11853;
												assign node11853 = (inp[10]) ? 4'b0000 : node11854;
													assign node11854 = (inp[0]) ? 4'b0001 : node11855;
														assign node11855 = (inp[12]) ? 4'b0001 : 4'b0000;
				assign node11862 = (inp[0]) ? node12906 : node11863;
					assign node11863 = (inp[6]) ? node12167 : node11864;
						assign node11864 = (inp[2]) ? node12134 : node11865;
							assign node11865 = (inp[5]) ? node11931 : node11866;
								assign node11866 = (inp[3]) ? node11868 : 4'b0010;
									assign node11868 = (inp[4]) ? node11886 : node11869;
										assign node11869 = (inp[7]) ? 4'b0010 : node11870;
											assign node11870 = (inp[13]) ? node11872 : 4'b0010;
												assign node11872 = (inp[10]) ? node11878 : node11873;
													assign node11873 = (inp[1]) ? node11875 : 4'b0010;
														assign node11875 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node11878 = (inp[1]) ? node11882 : node11879;
														assign node11879 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node11882 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node11886 = (inp[7]) ? node11918 : node11887;
											assign node11887 = (inp[11]) ? node11905 : node11888;
												assign node11888 = (inp[1]) ? node11896 : node11889;
													assign node11889 = (inp[14]) ? node11891 : 4'b1001;
														assign node11891 = (inp[13]) ? node11893 : 4'b0000;
															assign node11893 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node11896 = (inp[14]) ? node11898 : 4'b0000;
														assign node11898 = (inp[10]) ? node11900 : 4'b0001;
															assign node11900 = (inp[12]) ? 4'b1001 : node11901;
																assign node11901 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node11905 = (inp[1]) ? node11915 : node11906;
													assign node11906 = (inp[12]) ? node11912 : node11907;
														assign node11907 = (inp[10]) ? node11909 : 4'b1001;
															assign node11909 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node11912 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node11915 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node11918 = (inp[13]) ? node11920 : 4'b0010;
												assign node11920 = (inp[10]) ? node11924 : node11921;
													assign node11921 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node11924 = (inp[1]) ? node11926 : 4'b0001;
														assign node11926 = (inp[12]) ? node11928 : 4'b0000;
															assign node11928 = (inp[11]) ? 4'b0000 : 4'b0010;
								assign node11931 = (inp[1]) ? node12039 : node11932;
									assign node11932 = (inp[11]) ? node11992 : node11933;
										assign node11933 = (inp[14]) ? node11967 : node11934;
											assign node11934 = (inp[3]) ? node11948 : node11935;
												assign node11935 = (inp[7]) ? node11943 : node11936;
													assign node11936 = (inp[4]) ? node11938 : 4'b0001;
														assign node11938 = (inp[10]) ? node11940 : 4'b0101;
															assign node11940 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node11943 = (inp[13]) ? node11945 : 4'b0001;
														assign node11945 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node11948 = (inp[13]) ? node11958 : node11949;
													assign node11949 = (inp[12]) ? node11953 : node11950;
														assign node11950 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node11953 = (inp[7]) ? 4'b0101 : node11954;
															assign node11954 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node11958 = (inp[12]) ? node11962 : node11959;
														assign node11959 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node11962 = (inp[7]) ? 4'b1101 : node11963;
															assign node11963 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node11967 = (inp[13]) ? node11981 : node11968;
												assign node11968 = (inp[12]) ? node11976 : node11969;
													assign node11969 = (inp[10]) ? 4'b1000 : node11970;
														assign node11970 = (inp[3]) ? node11972 : 4'b0000;
															assign node11972 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node11976 = (inp[7]) ? 4'b0100 : node11977;
														assign node11977 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node11981 = (inp[10]) ? node11987 : node11982;
													assign node11982 = (inp[3]) ? 4'b1100 : node11983;
														assign node11983 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node11987 = (inp[12]) ? 4'b1000 : node11988;
														assign node11988 = (inp[3]) ? 4'b0100 : 4'b0000;
										assign node11992 = (inp[13]) ? node12014 : node11993;
											assign node11993 = (inp[3]) ? node12005 : node11994;
												assign node11994 = (inp[10]) ? node11996 : 4'b0001;
													assign node11996 = (inp[12]) ? node12000 : node11997;
														assign node11997 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node12000 = (inp[7]) ? 4'b0001 : node12001;
															assign node12001 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node12005 = (inp[4]) ? node12011 : node12006;
													assign node12006 = (inp[10]) ? node12008 : 4'b0101;
														assign node12008 = (inp[7]) ? 4'b0101 : 4'b1101;
													assign node12011 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node12014 = (inp[10]) ? node12022 : node12015;
												assign node12015 = (inp[3]) ? node12017 : 4'b1001;
													assign node12017 = (inp[14]) ? 4'b1101 : node12018;
														assign node12018 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node12022 = (inp[12]) ? node12032 : node12023;
													assign node12023 = (inp[14]) ? node12025 : 4'b0101;
														assign node12025 = (inp[7]) ? node12027 : 4'b0101;
															assign node12027 = (inp[4]) ? 4'b0001 : node12028;
																assign node12028 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node12032 = (inp[14]) ? 4'b1101 : node12033;
														assign node12033 = (inp[3]) ? node12035 : 4'b1001;
															assign node12035 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node12039 = (inp[11]) ? node12083 : node12040;
										assign node12040 = (inp[14]) ? node12062 : node12041;
											assign node12041 = (inp[13]) ? node12053 : node12042;
												assign node12042 = (inp[10]) ? node12048 : node12043;
													assign node12043 = (inp[4]) ? 4'b1000 : node12044;
														assign node12044 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node12048 = (inp[4]) ? 4'b1100 : node12049;
														assign node12049 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node12053 = (inp[3]) ? node12057 : node12054;
													assign node12054 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node12057 = (inp[4]) ? 4'b0000 : node12058;
														assign node12058 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node12062 = (inp[13]) ? node12072 : node12063;
												assign node12063 = (inp[3]) ? node12069 : node12064;
													assign node12064 = (inp[4]) ? node12066 : 4'b0001;
														assign node12066 = (inp[7]) ? 4'b0001 : 4'b1101;
													assign node12069 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node12072 = (inp[10]) ? node12078 : node12073;
													assign node12073 = (inp[3]) ? node12075 : 4'b1001;
														assign node12075 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12078 = (inp[3]) ? 4'b0001 : node12079;
														assign node12079 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node12083 = (inp[13]) ? node12103 : node12084;
											assign node12084 = (inp[10]) ? node12094 : node12085;
												assign node12085 = (inp[12]) ? node12089 : node12086;
													assign node12086 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node12089 = (inp[3]) ? node12091 : 4'b0000;
														assign node12091 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node12094 = (inp[3]) ? 4'b1100 : node12095;
													assign node12095 = (inp[12]) ? node12097 : 4'b1000;
														assign node12097 = (inp[4]) ? node12099 : 4'b1000;
															assign node12099 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node12103 = (inp[10]) ? node12117 : node12104;
												assign node12104 = (inp[12]) ? node12110 : node12105;
													assign node12105 = (inp[3]) ? node12107 : 4'b0100;
														assign node12107 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12110 = (inp[3]) ? 4'b1100 : node12111;
														assign node12111 = (inp[4]) ? node12113 : 4'b1000;
															assign node12113 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node12117 = (inp[14]) ? node12129 : node12118;
													assign node12118 = (inp[3]) ? node12124 : node12119;
														assign node12119 = (inp[4]) ? 4'b0100 : node12120;
															assign node12120 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node12124 = (inp[7]) ? node12126 : 4'b0000;
															assign node12126 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12129 = (inp[3]) ? 4'b0000 : node12130;
														assign node12130 = (inp[4]) ? 4'b0100 : 4'b0000;
							assign node12134 = (inp[5]) ? node12136 : 4'b0010;
								assign node12136 = (inp[3]) ? node12138 : 4'b0010;
									assign node12138 = (inp[7]) ? node12156 : node12139;
										assign node12139 = (inp[4]) ? node12145 : node12140;
											assign node12140 = (inp[13]) ? node12142 : 4'b0010;
												assign node12142 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node12145 = (inp[1]) ? node12149 : node12146;
												assign node12146 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node12149 = (inp[14]) ? node12153 : node12150;
													assign node12150 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node12153 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node12156 = (inp[1]) ? node12158 : 4'b0010;
											assign node12158 = (inp[14]) ? node12160 : 4'b0010;
												assign node12160 = (inp[4]) ? node12162 : 4'b0010;
													assign node12162 = (inp[12]) ? 4'b0010 : node12163;
														assign node12163 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node12167 = (inp[5]) ? node12527 : node12168;
							assign node12168 = (inp[11]) ? node12364 : node12169;
								assign node12169 = (inp[3]) ? node12269 : node12170;
									assign node12170 = (inp[4]) ? node12210 : node12171;
										assign node12171 = (inp[10]) ? node12187 : node12172;
											assign node12172 = (inp[13]) ? node12180 : node12173;
												assign node12173 = (inp[12]) ? 4'b0000 : node12174;
													assign node12174 = (inp[1]) ? 4'b0001 : node12175;
														assign node12175 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node12180 = (inp[2]) ? node12182 : 4'b1001;
													assign node12182 = (inp[1]) ? node12184 : 4'b1001;
														assign node12184 = (inp[14]) ? 4'b1001 : 4'b0000;
											assign node12187 = (inp[13]) ? node12201 : node12188;
												assign node12188 = (inp[12]) ? node12194 : node12189;
													assign node12189 = (inp[1]) ? node12191 : 4'b1000;
														assign node12191 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node12194 = (inp[14]) ? node12198 : node12195;
														assign node12195 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node12198 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node12201 = (inp[12]) ? 4'b1000 : node12202;
													assign node12202 = (inp[7]) ? node12206 : node12203;
														assign node12203 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node12206 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node12210 = (inp[7]) ? node12240 : node12211;
											assign node12211 = (inp[13]) ? node12227 : node12212;
												assign node12212 = (inp[10]) ? node12220 : node12213;
													assign node12213 = (inp[1]) ? node12217 : node12214;
														assign node12214 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node12217 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node12220 = (inp[14]) ? node12224 : node12221;
														assign node12221 = (inp[12]) ? 4'b1100 : 4'b1101;
														assign node12224 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node12227 = (inp[2]) ? node12233 : node12228;
													assign node12228 = (inp[10]) ? node12230 : 4'b0001;
														assign node12230 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12233 = (inp[14]) ? node12237 : node12234;
														assign node12234 = (inp[1]) ? 4'b0100 : 4'b1101;
														assign node12237 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node12240 = (inp[10]) ? node12252 : node12241;
												assign node12241 = (inp[14]) ? node12249 : node12242;
													assign node12242 = (inp[1]) ? node12244 : 4'b1001;
														assign node12244 = (inp[13]) ? node12246 : 4'b1000;
															assign node12246 = (inp[2]) ? 4'b0100 : 4'b1000;
													assign node12249 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node12252 = (inp[13]) ? node12258 : node12253;
													assign node12253 = (inp[2]) ? node12255 : 4'b0000;
														assign node12255 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node12258 = (inp[12]) ? node12266 : node12259;
														assign node12259 = (inp[1]) ? node12263 : node12260;
															assign node12260 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node12263 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node12266 = (inp[1]) ? 4'b0100 : 4'b1000;
									assign node12269 = (inp[2]) ? node12311 : node12270;
										assign node12270 = (inp[10]) ? node12298 : node12271;
											assign node12271 = (inp[4]) ? node12281 : node12272;
												assign node12272 = (inp[12]) ? node12276 : node12273;
													assign node12273 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node12276 = (inp[14]) ? node12278 : 4'b0001;
														assign node12278 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node12281 = (inp[7]) ? node12293 : node12282;
													assign node12282 = (inp[13]) ? node12284 : 4'b0101;
														assign node12284 = (inp[12]) ? node12290 : node12285;
															assign node12285 = (inp[14]) ? 4'b0000 : node12286;
																assign node12286 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node12290 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node12293 = (inp[12]) ? 4'b0101 : node12294;
														assign node12294 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node12298 = (inp[1]) ? node12304 : node12299;
												assign node12299 = (inp[7]) ? node12301 : 4'b1101;
													assign node12301 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node12304 = (inp[12]) ? node12306 : 4'b0001;
													assign node12306 = (inp[7]) ? node12308 : 4'b1000;
														assign node12308 = (inp[14]) ? 4'b1101 : 4'b1001;
										assign node12311 = (inp[13]) ? node12331 : node12312;
											assign node12312 = (inp[12]) ? node12320 : node12313;
												assign node12313 = (inp[10]) ? node12315 : 4'b0101;
													assign node12315 = (inp[7]) ? 4'b1100 : node12316;
														assign node12316 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node12320 = (inp[1]) ? node12328 : node12321;
													assign node12321 = (inp[14]) ? node12323 : 4'b0101;
														assign node12323 = (inp[7]) ? 4'b0100 : node12324;
															assign node12324 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12328 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node12331 = (inp[4]) ? node12347 : node12332;
												assign node12332 = (inp[10]) ? node12342 : node12333;
													assign node12333 = (inp[12]) ? node12339 : node12334;
														assign node12334 = (inp[7]) ? node12336 : 4'b1101;
															assign node12336 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node12339 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node12342 = (inp[12]) ? 4'b1101 : node12343;
														assign node12343 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node12347 = (inp[7]) ? node12357 : node12348;
													assign node12348 = (inp[10]) ? node12354 : node12349;
														assign node12349 = (inp[12]) ? 4'b0001 : node12350;
															assign node12350 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node12354 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12357 = (inp[10]) ? 4'b0001 : node12358;
														assign node12358 = (inp[1]) ? 4'b0000 : node12359;
															assign node12359 = (inp[14]) ? 4'b1100 : 4'b1101;
								assign node12364 = (inp[1]) ? node12438 : node12365;
									assign node12365 = (inp[3]) ? node12399 : node12366;
										assign node12366 = (inp[13]) ? node12372 : node12367;
											assign node12367 = (inp[4]) ? node12369 : 4'b0001;
												assign node12369 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node12372 = (inp[10]) ? node12380 : node12373;
												assign node12373 = (inp[7]) ? 4'b1001 : node12374;
													assign node12374 = (inp[12]) ? 4'b1101 : node12375;
														assign node12375 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node12380 = (inp[12]) ? node12392 : node12381;
													assign node12381 = (inp[2]) ? node12387 : node12382;
														assign node12382 = (inp[4]) ? 4'b0000 : node12383;
															assign node12383 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node12387 = (inp[4]) ? 4'b0101 : node12388;
															assign node12388 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node12392 = (inp[2]) ? node12396 : node12393;
														assign node12393 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node12396 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node12399 = (inp[2]) ? node12419 : node12400;
											assign node12400 = (inp[12]) ? node12412 : node12401;
												assign node12401 = (inp[10]) ? node12407 : node12402;
													assign node12402 = (inp[4]) ? 4'b1100 : node12403;
														assign node12403 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12407 = (inp[7]) ? 4'b0100 : node12408;
														assign node12408 = (inp[4]) ? 4'b1001 : 4'b0100;
												assign node12412 = (inp[10]) ? node12414 : 4'b0100;
													assign node12414 = (inp[4]) ? 4'b1100 : node12415;
														assign node12415 = (inp[13]) ? 4'b1100 : 4'b1000;
											assign node12419 = (inp[7]) ? node12431 : node12420;
												assign node12420 = (inp[4]) ? node12424 : node12421;
													assign node12421 = (inp[14]) ? 4'b0001 : 4'b1101;
													assign node12424 = (inp[13]) ? node12426 : 4'b0001;
														assign node12426 = (inp[12]) ? 4'b1000 : node12427;
															assign node12427 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node12431 = (inp[13]) ? 4'b1101 : node12432;
													assign node12432 = (inp[12]) ? 4'b0101 : node12433;
														assign node12433 = (inp[10]) ? 4'b1101 : 4'b0101;
									assign node12438 = (inp[10]) ? node12490 : node12439;
										assign node12439 = (inp[7]) ? node12477 : node12440;
											assign node12440 = (inp[12]) ? node12458 : node12441;
												assign node12441 = (inp[2]) ? node12449 : node12442;
													assign node12442 = (inp[13]) ? node12446 : node12443;
														assign node12443 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12446 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node12449 = (inp[13]) ? node12453 : node12450;
														assign node12450 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12453 = (inp[14]) ? node12455 : 4'b1000;
															assign node12455 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node12458 = (inp[13]) ? node12468 : node12459;
													assign node12459 = (inp[4]) ? node12465 : node12460;
														assign node12460 = (inp[3]) ? node12462 : 4'b0000;
															assign node12462 = (inp[2]) ? 4'b0100 : 4'b1000;
														assign node12465 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node12468 = (inp[2]) ? node12472 : node12469;
														assign node12469 = (inp[4]) ? 4'b0000 : 4'b1100;
														assign node12472 = (inp[4]) ? node12474 : 4'b1000;
															assign node12474 = (inp[14]) ? 4'b1100 : 4'b1000;
											assign node12477 = (inp[3]) ? node12483 : node12478;
												assign node12478 = (inp[13]) ? node12480 : 4'b1000;
													assign node12480 = (inp[2]) ? 4'b1000 : 4'b0100;
												assign node12483 = (inp[4]) ? 4'b1100 : node12484;
													assign node12484 = (inp[2]) ? node12486 : 4'b1000;
														assign node12486 = (inp[14]) ? 4'b1100 : 4'b0100;
										assign node12490 = (inp[13]) ? node12510 : node12491;
											assign node12491 = (inp[3]) ? node12499 : node12492;
												assign node12492 = (inp[7]) ? 4'b1000 : node12493;
													assign node12493 = (inp[2]) ? node12495 : 4'b0000;
														assign node12495 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node12499 = (inp[2]) ? node12507 : node12500;
													assign node12500 = (inp[4]) ? node12504 : node12501;
														assign node12501 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node12504 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node12507 = (inp[7]) ? 4'b1100 : 4'b0000;
											assign node12510 = (inp[7]) ? node12516 : node12511;
												assign node12511 = (inp[3]) ? 4'b0000 : node12512;
													assign node12512 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node12516 = (inp[12]) ? node12522 : node12517;
													assign node12517 = (inp[2]) ? 4'b0100 : node12518;
														assign node12518 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node12522 = (inp[4]) ? node12524 : 4'b0000;
														assign node12524 = (inp[14]) ? 4'b0100 : 4'b0000;
							assign node12527 = (inp[3]) ? node12727 : node12528;
								assign node12528 = (inp[1]) ? node12634 : node12529;
									assign node12529 = (inp[13]) ? node12583 : node12530;
										assign node12530 = (inp[4]) ? node12554 : node12531;
											assign node12531 = (inp[10]) ? node12541 : node12532;
												assign node12532 = (inp[11]) ? node12534 : 4'b0001;
													assign node12534 = (inp[12]) ? node12538 : node12535;
														assign node12535 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node12538 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node12541 = (inp[7]) ? node12549 : node12542;
													assign node12542 = (inp[12]) ? node12544 : 4'b0100;
														assign node12544 = (inp[2]) ? node12546 : 4'b0100;
															assign node12546 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node12549 = (inp[12]) ? 4'b1001 : node12550;
														assign node12550 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node12554 = (inp[2]) ? node12568 : node12555;
												assign node12555 = (inp[12]) ? node12561 : node12556;
													assign node12556 = (inp[7]) ? 4'b1000 : node12557;
														assign node12557 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node12561 = (inp[11]) ? 4'b1000 : node12562;
														assign node12562 = (inp[14]) ? node12564 : 4'b0000;
															assign node12564 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node12568 = (inp[10]) ? node12578 : node12569;
													assign node12569 = (inp[7]) ? node12575 : node12570;
														assign node12570 = (inp[14]) ? 4'b0001 : node12571;
															assign node12571 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12575 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node12578 = (inp[11]) ? 4'b0001 : node12579;
														assign node12579 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node12583 = (inp[4]) ? node12611 : node12584;
											assign node12584 = (inp[10]) ? node12592 : node12585;
												assign node12585 = (inp[7]) ? node12587 : 4'b1101;
													assign node12587 = (inp[2]) ? node12589 : 4'b1001;
														assign node12589 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node12592 = (inp[14]) ? node12600 : node12593;
													assign node12593 = (inp[12]) ? node12595 : 4'b1101;
														assign node12595 = (inp[7]) ? 4'b1100 : node12596;
															assign node12596 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node12600 = (inp[7]) ? node12606 : node12601;
														assign node12601 = (inp[11]) ? 4'b0100 : node12602;
															assign node12602 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node12606 = (inp[2]) ? 4'b1001 : node12607;
															assign node12607 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node12611 = (inp[2]) ? node12623 : node12612;
												assign node12612 = (inp[10]) ? node12618 : node12613;
													assign node12613 = (inp[14]) ? node12615 : 4'b0001;
														assign node12615 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node12618 = (inp[11]) ? node12620 : 4'b0000;
														assign node12620 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node12623 = (inp[12]) ? 4'b1001 : node12624;
													assign node12624 = (inp[7]) ? node12628 : node12625;
														assign node12625 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node12628 = (inp[10]) ? 4'b1001 : node12629;
															assign node12629 = (inp[11]) ? 4'b0001 : 4'b1001;
									assign node12634 = (inp[11]) ? node12684 : node12635;
										assign node12635 = (inp[4]) ? node12663 : node12636;
											assign node12636 = (inp[7]) ? node12644 : node12637;
												assign node12637 = (inp[13]) ? node12639 : 4'b1001;
													assign node12639 = (inp[12]) ? node12641 : 4'b0000;
														assign node12641 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node12644 = (inp[12]) ? node12654 : node12645;
													assign node12645 = (inp[10]) ? node12651 : node12646;
														assign node12646 = (inp[2]) ? 4'b1001 : node12647;
															assign node12647 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12651 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node12654 = (inp[2]) ? node12660 : node12655;
														assign node12655 = (inp[10]) ? node12657 : 4'b0101;
															assign node12657 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node12660 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node12663 = (inp[10]) ? node12679 : node12664;
												assign node12664 = (inp[14]) ? node12670 : node12665;
													assign node12665 = (inp[2]) ? node12667 : 4'b1000;
														assign node12667 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node12670 = (inp[13]) ? node12674 : node12671;
														assign node12671 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node12674 = (inp[2]) ? 4'b0000 : node12675;
															assign node12675 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node12679 = (inp[2]) ? node12681 : 4'b0100;
													assign node12681 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node12684 = (inp[13]) ? node12710 : node12685;
											assign node12685 = (inp[2]) ? node12697 : node12686;
												assign node12686 = (inp[4]) ? node12692 : node12687;
													assign node12687 = (inp[12]) ? 4'b1000 : node12688;
														assign node12688 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12692 = (inp[10]) ? node12694 : 4'b0100;
														assign node12694 = (inp[7]) ? 4'b0100 : 4'b1000;
												assign node12697 = (inp[7]) ? node12705 : node12698;
													assign node12698 = (inp[4]) ? node12702 : node12699;
														assign node12699 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node12702 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node12705 = (inp[10]) ? 4'b1000 : node12706;
														assign node12706 = (inp[14]) ? 4'b1000 : 4'b1100;
											assign node12710 = (inp[10]) ? node12722 : node12711;
												assign node12711 = (inp[2]) ? node12717 : node12712;
													assign node12712 = (inp[12]) ? node12714 : 4'b0000;
														assign node12714 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node12717 = (inp[7]) ? 4'b1000 : node12718;
														assign node12718 = (inp[12]) ? 4'b0000 : 4'b1100;
												assign node12722 = (inp[7]) ? node12724 : 4'b0000;
													assign node12724 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node12727 = (inp[4]) ? node12817 : node12728;
									assign node12728 = (inp[11]) ? node12776 : node12729;
										assign node12729 = (inp[13]) ? node12755 : node12730;
											assign node12730 = (inp[2]) ? node12744 : node12731;
												assign node12731 = (inp[7]) ? node12741 : node12732;
													assign node12732 = (inp[1]) ? node12736 : node12733;
														assign node12733 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12736 = (inp[10]) ? 4'b1000 : node12737;
															assign node12737 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node12741 = (inp[1]) ? 4'b0001 : 4'b1000;
												assign node12744 = (inp[1]) ? node12750 : node12745;
													assign node12745 = (inp[12]) ? node12747 : 4'b1000;
														assign node12747 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12750 = (inp[7]) ? node12752 : 4'b0000;
														assign node12752 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node12755 = (inp[10]) ? node12763 : node12756;
												assign node12756 = (inp[7]) ? node12758 : 4'b0001;
													assign node12758 = (inp[12]) ? 4'b1000 : node12759;
														assign node12759 = (inp[2]) ? 4'b0001 : 4'b1000;
												assign node12763 = (inp[1]) ? node12771 : node12764;
													assign node12764 = (inp[2]) ? node12768 : node12765;
														assign node12765 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node12768 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node12771 = (inp[12]) ? node12773 : 4'b1000;
														assign node12773 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node12776 = (inp[1]) ? node12800 : node12777;
											assign node12777 = (inp[12]) ? node12787 : node12778;
												assign node12778 = (inp[7]) ? node12784 : node12779;
													assign node12779 = (inp[2]) ? node12781 : 4'b1001;
														assign node12781 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node12784 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node12787 = (inp[13]) ? node12789 : 4'b1001;
													assign node12789 = (inp[2]) ? node12795 : node12790;
														assign node12790 = (inp[7]) ? node12792 : 4'b1001;
															assign node12792 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node12795 = (inp[10]) ? node12797 : 4'b1000;
															assign node12797 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node12800 = (inp[10]) ? node12810 : node12801;
												assign node12801 = (inp[13]) ? node12805 : node12802;
													assign node12802 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node12805 = (inp[7]) ? node12807 : 4'b1000;
														assign node12807 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node12810 = (inp[2]) ? node12812 : 4'b0000;
													assign node12812 = (inp[13]) ? 4'b0000 : node12813;
														assign node12813 = (inp[7]) ? 4'b1000 : 4'b0000;
									assign node12817 = (inp[13]) ? node12875 : node12818;
										assign node12818 = (inp[1]) ? node12848 : node12819;
											assign node12819 = (inp[14]) ? node12833 : node12820;
												assign node12820 = (inp[2]) ? node12826 : node12821;
													assign node12821 = (inp[12]) ? node12823 : 4'b0001;
														assign node12823 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node12826 = (inp[11]) ? 4'b1000 : node12827;
														assign node12827 = (inp[7]) ? 4'b1000 : node12828;
															assign node12828 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node12833 = (inp[12]) ? 4'b1000 : node12834;
													assign node12834 = (inp[11]) ? node12842 : node12835;
														assign node12835 = (inp[2]) ? node12839 : node12836;
															assign node12836 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node12839 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node12842 = (inp[7]) ? 4'b0001 : node12843;
															assign node12843 = (inp[10]) ? 4'b1000 : 4'b0001;
											assign node12848 = (inp[11]) ? node12866 : node12849;
												assign node12849 = (inp[7]) ? node12857 : node12850;
													assign node12850 = (inp[14]) ? 4'b0000 : node12851;
														assign node12851 = (inp[2]) ? 4'b0001 : node12852;
															assign node12852 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node12857 = (inp[12]) ? node12863 : node12858;
														assign node12858 = (inp[2]) ? 4'b0001 : node12859;
															assign node12859 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node12863 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node12866 = (inp[10]) ? 4'b0000 : node12867;
													assign node12867 = (inp[2]) ? node12869 : 4'b1000;
														assign node12869 = (inp[14]) ? node12871 : 4'b0000;
															assign node12871 = (inp[7]) ? 4'b1000 : 4'b0000;
										assign node12875 = (inp[1]) ? node12897 : node12876;
											assign node12876 = (inp[12]) ? node12890 : node12877;
												assign node12877 = (inp[7]) ? node12881 : node12878;
													assign node12878 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node12881 = (inp[11]) ? 4'b0000 : node12882;
														assign node12882 = (inp[10]) ? node12886 : node12883;
															assign node12883 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node12886 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node12890 = (inp[7]) ? node12892 : 4'b0000;
													assign node12892 = (inp[10]) ? 4'b0000 : node12893;
														assign node12893 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node12897 = (inp[2]) ? 4'b0000 : node12898;
												assign node12898 = (inp[7]) ? node12900 : 4'b0000;
													assign node12900 = (inp[10]) ? 4'b0000 : node12901;
														assign node12901 = (inp[11]) ? 4'b0000 : 4'b0001;
					assign node12906 = (inp[6]) ? node12908 : 4'b0000;
						assign node12908 = (inp[2]) ? node13136 : node12909;
							assign node12909 = (inp[5]) ? node12967 : node12910;
								assign node12910 = (inp[4]) ? node12924 : node12911;
									assign node12911 = (inp[12]) ? 4'b0000 : node12912;
										assign node12912 = (inp[1]) ? node12914 : 4'b0000;
											assign node12914 = (inp[14]) ? node12916 : 4'b0000;
												assign node12916 = (inp[3]) ? node12918 : 4'b0000;
													assign node12918 = (inp[11]) ? 4'b0000 : node12919;
														assign node12919 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node12924 = (inp[3]) ? node12926 : 4'b0000;
										assign node12926 = (inp[7]) ? node12960 : node12927;
											assign node12927 = (inp[1]) ? node12943 : node12928;
												assign node12928 = (inp[14]) ? node12936 : node12929;
													assign node12929 = (inp[13]) ? node12931 : 4'b0001;
														assign node12931 = (inp[12]) ? 4'b1001 : node12932;
															assign node12932 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node12936 = (inp[10]) ? node12938 : 4'b1000;
														assign node12938 = (inp[12]) ? 4'b1001 : node12939;
															assign node12939 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node12943 = (inp[14]) ? node12951 : node12944;
													assign node12944 = (inp[13]) ? node12946 : 4'b1000;
														assign node12946 = (inp[10]) ? 4'b0000 : node12947;
															assign node12947 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node12951 = (inp[11]) ? node12955 : node12952;
														assign node12952 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node12955 = (inp[10]) ? 4'b0000 : node12956;
															assign node12956 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node12960 = (inp[11]) ? 4'b0000 : node12961;
												assign node12961 = (inp[12]) ? 4'b0000 : node12962;
													assign node12962 = (inp[10]) ? 4'b0001 : 4'b0000;
								assign node12967 = (inp[1]) ? node13067 : node12968;
									assign node12968 = (inp[3]) ? node13018 : node12969;
										assign node12969 = (inp[13]) ? node12993 : node12970;
											assign node12970 = (inp[14]) ? node12980 : node12971;
												assign node12971 = (inp[7]) ? 4'b0001 : node12972;
													assign node12972 = (inp[4]) ? node12974 : 4'b0001;
														assign node12974 = (inp[11]) ? node12976 : 4'b0101;
															assign node12976 = (inp[10]) ? 4'b0000 : 4'b0101;
												assign node12980 = (inp[11]) ? node12988 : node12981;
													assign node12981 = (inp[12]) ? node12985 : node12982;
														assign node12982 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node12985 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node12988 = (inp[7]) ? 4'b0001 : node12989;
														assign node12989 = (inp[4]) ? 4'b0101 : 4'b1001;
											assign node12993 = (inp[4]) ? node12999 : node12994;
												assign node12994 = (inp[11]) ? 4'b1001 : node12995;
													assign node12995 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node12999 = (inp[12]) ? node13011 : node13000;
													assign node13000 = (inp[10]) ? node13004 : node13001;
														assign node13001 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node13004 = (inp[7]) ? node13006 : 4'b1001;
															assign node13006 = (inp[11]) ? 4'b0000 : node13007;
																assign node13007 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13011 = (inp[7]) ? 4'b1001 : node13012;
														assign node13012 = (inp[11]) ? node13014 : 4'b1001;
															assign node13014 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node13018 = (inp[11]) ? node13040 : node13019;
											assign node13019 = (inp[13]) ? node13031 : node13020;
												assign node13020 = (inp[4]) ? node13024 : node13021;
													assign node13021 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node13024 = (inp[14]) ? 4'b1000 : node13025;
														assign node13025 = (inp[12]) ? 4'b1001 : node13026;
															assign node13026 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node13031 = (inp[4]) ? node13033 : 4'b1000;
													assign node13033 = (inp[14]) ? node13035 : 4'b0000;
														assign node13035 = (inp[10]) ? 4'b0001 : node13036;
															assign node13036 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node13040 = (inp[4]) ? node13056 : node13041;
												assign node13041 = (inp[13]) ? node13047 : node13042;
													assign node13042 = (inp[10]) ? 4'b0001 : node13043;
														assign node13043 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13047 = (inp[10]) ? node13053 : node13048;
														assign node13048 = (inp[7]) ? 4'b0000 : node13049;
															assign node13049 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13053 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node13056 = (inp[13]) ? node13060 : node13057;
													assign node13057 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node13060 = (inp[12]) ? node13062 : 4'b0000;
														assign node13062 = (inp[14]) ? 4'b0000 : node13063;
															assign node13063 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node13067 = (inp[11]) ? node13097 : node13068;
										assign node13068 = (inp[3]) ? node13080 : node13069;
											assign node13069 = (inp[14]) ? node13077 : node13070;
												assign node13070 = (inp[10]) ? 4'b1001 : node13071;
													assign node13071 = (inp[7]) ? 4'b1000 : node13072;
														assign node13072 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node13077 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node13080 = (inp[13]) ? node13092 : node13081;
												assign node13081 = (inp[7]) ? node13087 : node13082;
													assign node13082 = (inp[10]) ? node13084 : 4'b0001;
														assign node13084 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node13087 = (inp[14]) ? 4'b0000 : node13088;
														assign node13088 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node13092 = (inp[10]) ? node13094 : 4'b0000;
													assign node13094 = (inp[4]) ? 4'b0000 : 4'b1001;
										assign node13097 = (inp[3]) ? node13121 : node13098;
											assign node13098 = (inp[7]) ? node13112 : node13099;
												assign node13099 = (inp[10]) ? node13107 : node13100;
													assign node13100 = (inp[13]) ? 4'b1000 : node13101;
														assign node13101 = (inp[12]) ? node13103 : 4'b1100;
															assign node13103 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node13107 = (inp[12]) ? 4'b0100 : node13108;
														assign node13108 = (inp[4]) ? 4'b0000 : 4'b1000;
												assign node13112 = (inp[10]) ? node13118 : node13113;
													assign node13113 = (inp[13]) ? 4'b1000 : node13114;
														assign node13114 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13118 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node13121 = (inp[13]) ? 4'b0000 : node13122;
												assign node13122 = (inp[4]) ? 4'b0000 : node13123;
													assign node13123 = (inp[12]) ? node13129 : node13124;
														assign node13124 = (inp[10]) ? 4'b1000 : node13125;
															assign node13125 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node13129 = (inp[7]) ? node13131 : 4'b1000;
															assign node13131 = (inp[10]) ? 4'b0000 : 4'b1000;
							assign node13136 = (inp[5]) ? node13138 : 4'b0000;
								assign node13138 = (inp[3]) ? node13140 : 4'b0000;
									assign node13140 = (inp[7]) ? node13184 : node13141;
										assign node13141 = (inp[1]) ? node13165 : node13142;
											assign node13142 = (inp[4]) ? node13148 : node13143;
												assign node13143 = (inp[14]) ? node13145 : 4'b0000;
													assign node13145 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node13148 = (inp[13]) ? node13160 : node13149;
													assign node13149 = (inp[10]) ? node13151 : 4'b0001;
														assign node13151 = (inp[14]) ? node13155 : node13152;
															assign node13152 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node13155 = (inp[12]) ? node13157 : 4'b0000;
																assign node13157 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node13160 = (inp[11]) ? 4'b0000 : node13161;
														assign node13161 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node13165 = (inp[12]) ? node13171 : node13166;
												assign node13166 = (inp[4]) ? node13168 : 4'b0000;
													assign node13168 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node13171 = (inp[11]) ? 4'b0000 : node13172;
													assign node13172 = (inp[4]) ? node13174 : 4'b0000;
														assign node13174 = (inp[14]) ? node13180 : node13175;
															assign node13175 = (inp[10]) ? 4'b0000 : node13176;
																assign node13176 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node13180 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node13184 = (inp[12]) ? 4'b0000 : node13185;
											assign node13185 = (inp[13]) ? node13187 : 4'b0000;
												assign node13187 = (inp[1]) ? 4'b0000 : node13188;
													assign node13188 = (inp[4]) ? 4'b0001 : 4'b0000;

endmodule