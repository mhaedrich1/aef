module dtc_split875_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node9;
	wire [15-1:0] node12;
	wire [15-1:0] node13;
	wire [15-1:0] node16;
	wire [15-1:0] node19;
	wire [15-1:0] node20;
	wire [15-1:0] node21;
	wire [15-1:0] node24;
	wire [15-1:0] node27;
	wire [15-1:0] node28;
	wire [15-1:0] node31;
	wire [15-1:0] node34;
	wire [15-1:0] node35;
	wire [15-1:0] node36;
	wire [15-1:0] node37;
	wire [15-1:0] node40;
	wire [15-1:0] node43;
	wire [15-1:0] node44;
	wire [15-1:0] node47;
	wire [15-1:0] node50;
	wire [15-1:0] node51;
	wire [15-1:0] node52;
	wire [15-1:0] node55;
	wire [15-1:0] node58;
	wire [15-1:0] node59;
	wire [15-1:0] node62;
	wire [15-1:0] node65;
	wire [15-1:0] node66;
	wire [15-1:0] node67;
	wire [15-1:0] node68;
	wire [15-1:0] node69;
	wire [15-1:0] node72;
	wire [15-1:0] node75;
	wire [15-1:0] node76;
	wire [15-1:0] node79;
	wire [15-1:0] node82;
	wire [15-1:0] node83;
	wire [15-1:0] node84;
	wire [15-1:0] node87;
	wire [15-1:0] node90;
	wire [15-1:0] node91;
	wire [15-1:0] node94;
	wire [15-1:0] node97;
	wire [15-1:0] node98;
	wire [15-1:0] node99;
	wire [15-1:0] node100;
	wire [15-1:0] node103;
	wire [15-1:0] node106;
	wire [15-1:0] node107;
	wire [15-1:0] node110;
	wire [15-1:0] node113;
	wire [15-1:0] node114;
	wire [15-1:0] node115;
	wire [15-1:0] node118;
	wire [15-1:0] node121;
	wire [15-1:0] node122;
	wire [15-1:0] node125;
	wire [15-1:0] node128;
	wire [15-1:0] node129;
	wire [15-1:0] node130;
	wire [15-1:0] node131;
	wire [15-1:0] node132;
	wire [15-1:0] node133;
	wire [15-1:0] node136;
	wire [15-1:0] node139;
	wire [15-1:0] node140;
	wire [15-1:0] node143;
	wire [15-1:0] node146;
	wire [15-1:0] node147;
	wire [15-1:0] node148;
	wire [15-1:0] node151;
	wire [15-1:0] node154;
	wire [15-1:0] node155;
	wire [15-1:0] node158;
	wire [15-1:0] node161;
	wire [15-1:0] node162;
	wire [15-1:0] node163;
	wire [15-1:0] node164;
	wire [15-1:0] node167;
	wire [15-1:0] node170;
	wire [15-1:0] node171;
	wire [15-1:0] node174;
	wire [15-1:0] node177;
	wire [15-1:0] node178;
	wire [15-1:0] node179;
	wire [15-1:0] node182;
	wire [15-1:0] node185;
	wire [15-1:0] node186;
	wire [15-1:0] node189;
	wire [15-1:0] node192;
	wire [15-1:0] node193;
	wire [15-1:0] node194;
	wire [15-1:0] node195;
	wire [15-1:0] node196;
	wire [15-1:0] node199;
	wire [15-1:0] node202;
	wire [15-1:0] node203;
	wire [15-1:0] node206;
	wire [15-1:0] node209;
	wire [15-1:0] node210;
	wire [15-1:0] node211;
	wire [15-1:0] node214;
	wire [15-1:0] node217;
	wire [15-1:0] node218;
	wire [15-1:0] node221;
	wire [15-1:0] node224;
	wire [15-1:0] node225;
	wire [15-1:0] node226;
	wire [15-1:0] node227;
	wire [15-1:0] node230;
	wire [15-1:0] node233;
	wire [15-1:0] node234;
	wire [15-1:0] node237;
	wire [15-1:0] node240;
	wire [15-1:0] node241;
	wire [15-1:0] node242;
	wire [15-1:0] node245;
	wire [15-1:0] node248;
	wire [15-1:0] node249;
	wire [15-1:0] node252;

	assign outp = (inp[10]) ? node128 : node1;
		assign node1 = (inp[8]) ? node65 : node2;
			assign node2 = (inp[1]) ? node34 : node3;
				assign node3 = (inp[7]) ? node19 : node4;
					assign node4 = (inp[2]) ? node12 : node5;
						assign node5 = (inp[3]) ? node9 : node6;
							assign node6 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
							assign node9 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
						assign node12 = (inp[13]) ? node16 : node13;
							assign node13 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node16 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
					assign node19 = (inp[0]) ? node27 : node20;
						assign node20 = (inp[3]) ? node24 : node21;
							assign node21 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node24 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node27 = (inp[14]) ? node31 : node28;
							assign node28 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node31 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
				assign node34 = (inp[13]) ? node50 : node35;
					assign node35 = (inp[4]) ? node43 : node36;
						assign node36 = (inp[14]) ? node40 : node37;
							assign node37 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node40 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node43 = (inp[7]) ? node47 : node44;
							assign node44 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node47 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
					assign node50 = (inp[3]) ? node58 : node51;
						assign node51 = (inp[7]) ? node55 : node52;
							assign node52 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node55 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node58 = (inp[12]) ? node62 : node59;
							assign node59 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node62 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
			assign node65 = (inp[9]) ? node97 : node66;
				assign node66 = (inp[7]) ? node82 : node67;
					assign node67 = (inp[12]) ? node75 : node68;
						assign node68 = (inp[11]) ? node72 : node69;
							assign node69 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node72 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node75 = (inp[14]) ? node79 : node76;
							assign node76 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node79 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
					assign node82 = (inp[3]) ? node90 : node83;
						assign node83 = (inp[4]) ? node87 : node84;
							assign node84 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node87 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node90 = (inp[0]) ? node94 : node91;
							assign node91 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node94 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
				assign node97 = (inp[14]) ? node113 : node98;
					assign node98 = (inp[11]) ? node106 : node99;
						assign node99 = (inp[0]) ? node103 : node100;
							assign node100 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node103 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node106 = (inp[12]) ? node110 : node107;
							assign node107 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node110 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node113 = (inp[5]) ? node121 : node114;
						assign node114 = (inp[0]) ? node118 : node115;
							assign node115 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node118 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node121 = (inp[4]) ? node125 : node122;
							assign node122 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node125 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
		assign node128 = (inp[3]) ? node192 : node129;
			assign node129 = (inp[0]) ? node161 : node130;
				assign node130 = (inp[14]) ? node146 : node131;
					assign node131 = (inp[13]) ? node139 : node132;
						assign node132 = (inp[8]) ? node136 : node133;
							assign node133 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node136 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node139 = (inp[1]) ? node143 : node140;
							assign node140 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node143 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
					assign node146 = (inp[4]) ? node154 : node147;
						assign node147 = (inp[7]) ? node151 : node148;
							assign node148 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node151 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node154 = (inp[5]) ? node158 : node155;
							assign node155 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node158 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
				assign node161 = (inp[7]) ? node177 : node162;
					assign node162 = (inp[5]) ? node170 : node163;
						assign node163 = (inp[11]) ? node167 : node164;
							assign node164 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node167 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node170 = (inp[13]) ? node174 : node171;
							assign node171 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node174 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node177 = (inp[2]) ? node185 : node178;
						assign node178 = (inp[9]) ? node182 : node179;
							assign node179 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node182 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node185 = (inp[5]) ? node189 : node186;
							assign node186 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node189 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
			assign node192 = (inp[12]) ? node224 : node193;
				assign node193 = (inp[4]) ? node209 : node194;
					assign node194 = (inp[2]) ? node202 : node195;
						assign node195 = (inp[6]) ? node199 : node196;
							assign node196 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node199 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node202 = (inp[6]) ? node206 : node203;
							assign node203 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node206 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node209 = (inp[0]) ? node217 : node210;
						assign node210 = (inp[9]) ? node214 : node211;
							assign node211 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node214 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node217 = (inp[7]) ? node221 : node218;
							assign node218 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node221 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
				assign node224 = (inp[11]) ? node240 : node225;
					assign node225 = (inp[6]) ? node233 : node226;
						assign node226 = (inp[0]) ? node230 : node227;
							assign node227 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node230 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node233 = (inp[8]) ? node237 : node234;
							assign node234 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node237 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node240 = (inp[13]) ? node248 : node241;
						assign node241 = (inp[1]) ? node245 : node242;
							assign node242 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node245 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node248 = (inp[8]) ? node252 : node249;
							assign node249 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node252 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;

endmodule