module dtc_split25_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node376;

	assign outp = (inp[0]) ? node138 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node43 : node4;
				assign node4 = (inp[3]) ? node30 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[1]) ? node21 : node8;
							assign node8 = (inp[7]) ? node10 : 3'b100;
								assign node10 = (inp[10]) ? node16 : node11;
									assign node11 = (inp[5]) ? 3'b100 : node12;
										assign node12 = (inp[2]) ? 3'b100 : 3'b000;
									assign node16 = (inp[11]) ? node18 : 3'b000;
										assign node18 = (inp[2]) ? 3'b000 : 3'b000;
							assign node21 = (inp[7]) ? node23 : 3'b000;
								assign node23 = (inp[2]) ? 3'b100 : node24;
									assign node24 = (inp[10]) ? node26 : 3'b101;
										assign node26 = (inp[8]) ? 3'b100 : 3'b101;
					assign node30 = (inp[4]) ? node32 : 3'b010;
						assign node32 = (inp[11]) ? node34 : 3'b010;
							assign node34 = (inp[1]) ? node36 : 3'b010;
								assign node36 = (inp[7]) ? node38 : 3'b010;
									assign node38 = (inp[2]) ? 3'b110 : node39;
										assign node39 = (inp[10]) ? 3'b010 : 3'b010;
				assign node43 = (inp[3]) ? node105 : node44;
					assign node44 = (inp[4]) ? node64 : node45;
						assign node45 = (inp[2]) ? node59 : node46;
							assign node46 = (inp[7]) ? 3'b001 : node47;
								assign node47 = (inp[1]) ? node53 : node48;
									assign node48 = (inp[5]) ? 3'b001 : node49;
										assign node49 = (inp[10]) ? 3'b001 : 3'b101;
									assign node53 = (inp[8]) ? 3'b001 : node54;
										assign node54 = (inp[11]) ? 3'b001 : 3'b100;
							assign node59 = (inp[7]) ? node61 : 3'b001;
								assign node61 = (inp[1]) ? 3'b100 : 3'b101;
						assign node64 = (inp[1]) ? node88 : node65;
							assign node65 = (inp[7]) ? node77 : node66;
								assign node66 = (inp[2]) ? node72 : node67;
									assign node67 = (inp[11]) ? 3'b101 : node68;
										assign node68 = (inp[8]) ? 3'b101 : 3'b111;
									assign node72 = (inp[11]) ? node74 : 3'b101;
										assign node74 = (inp[8]) ? 3'b011 : 3'b111;
								assign node77 = (inp[2]) ? node83 : node78;
									assign node78 = (inp[10]) ? 3'b011 : node79;
										assign node79 = (inp[5]) ? 3'b111 : 3'b011;
									assign node83 = (inp[5]) ? node85 : 3'b101;
										assign node85 = (inp[8]) ? 3'b001 : 3'b001;
							assign node88 = (inp[11]) ? node100 : node89;
								assign node89 = (inp[8]) ? node95 : node90;
									assign node90 = (inp[10]) ? node92 : 3'b001;
										assign node92 = (inp[7]) ? 3'b001 : 3'b100;
									assign node95 = (inp[5]) ? node97 : 3'b110;
										assign node97 = (inp[10]) ? 3'b001 : 3'b100;
								assign node100 = (inp[5]) ? node102 : 3'b110;
									assign node102 = (inp[7]) ? 3'b001 : 3'b110;
					assign node105 = (inp[1]) ? node107 : 3'b111;
						assign node107 = (inp[5]) ? node125 : node108;
							assign node108 = (inp[11]) ? node118 : node109;
								assign node109 = (inp[7]) ? node115 : node110;
									assign node110 = (inp[4]) ? node112 : 3'b111;
										assign node112 = (inp[10]) ? 3'b111 : 3'b011;
									assign node115 = (inp[2]) ? 3'b101 : 3'b111;
								assign node118 = (inp[10]) ? node120 : 3'b011;
									assign node120 = (inp[4]) ? node122 : 3'b101;
										assign node122 = (inp[7]) ? 3'b011 : 3'b001;
							assign node125 = (inp[7]) ? node133 : node126;
								assign node126 = (inp[4]) ? node128 : 3'b011;
									assign node128 = (inp[2]) ? node130 : 3'b001;
										assign node130 = (inp[8]) ? 3'b111 : 3'b001;
								assign node133 = (inp[10]) ? node135 : 3'b101;
									assign node135 = (inp[8]) ? 3'b001 : 3'b101;
		assign node138 = (inp[3]) ? node222 : node139;
			assign node139 = (inp[6]) ? node195 : node140;
				assign node140 = (inp[9]) ? node152 : node141;
					assign node141 = (inp[4]) ? node143 : 3'b010;
						assign node143 = (inp[1]) ? node149 : node144;
							assign node144 = (inp[11]) ? node146 : 3'b010;
								assign node146 = (inp[2]) ? 3'b010 : 3'b000;
							assign node149 = (inp[7]) ? 3'b010 : 3'b000;
					assign node152 = (inp[7]) ? node168 : node153;
						assign node153 = (inp[5]) ? node163 : node154;
							assign node154 = (inp[11]) ? 3'b010 : node155;
								assign node155 = (inp[4]) ? node157 : 3'b000;
									assign node157 = (inp[2]) ? node159 : 3'b010;
										assign node159 = (inp[1]) ? 3'b000 : 3'b000;
							assign node163 = (inp[10]) ? node165 : 3'b010;
								assign node165 = (inp[11]) ? 3'b000 : 3'b010;
						assign node168 = (inp[2]) ? node182 : node169;
							assign node169 = (inp[4]) ? node171 : 3'b000;
								assign node171 = (inp[10]) ? node177 : node172;
									assign node172 = (inp[5]) ? 3'b000 : node173;
										assign node173 = (inp[8]) ? 3'b010 : 3'b000;
									assign node177 = (inp[8]) ? node179 : 3'b010;
										assign node179 = (inp[5]) ? 3'b010 : 3'b000;
							assign node182 = (inp[4]) ? node184 : 3'b010;
								assign node184 = (inp[1]) ? node190 : node185;
									assign node185 = (inp[11]) ? node187 : 3'b000;
										assign node187 = (inp[8]) ? 3'b000 : 3'b010;
									assign node190 = (inp[10]) ? 3'b100 : node191;
										assign node191 = (inp[11]) ? 3'b000 : 3'b100;
				assign node195 = (inp[9]) ? node197 : 3'b000;
					assign node197 = (inp[4]) ? node199 : 3'b000;
						assign node199 = (inp[7]) ? node213 : node200;
							assign node200 = (inp[1]) ? 3'b100 : node201;
								assign node201 = (inp[11]) ? node207 : node202;
									assign node202 = (inp[5]) ? 3'b010 : node203;
										assign node203 = (inp[2]) ? 3'b110 : 3'b010;
									assign node207 = (inp[2]) ? 3'b100 : node208;
										assign node208 = (inp[5]) ? 3'b000 : 3'b100;
							assign node213 = (inp[1]) ? 3'b000 : node214;
								assign node214 = (inp[11]) ? node216 : 3'b010;
									assign node216 = (inp[2]) ? 3'b100 : node217;
										assign node217 = (inp[10]) ? 3'b100 : 3'b110;
			assign node222 = (inp[9]) ? node280 : node223;
				assign node223 = (inp[4]) ? node229 : node224;
					assign node224 = (inp[6]) ? 3'b000 : node225;
						assign node225 = (inp[1]) ? 3'b000 : 3'b001;
					assign node229 = (inp[1]) ? node253 : node230;
						assign node230 = (inp[7]) ? node240 : node231;
							assign node231 = (inp[6]) ? 3'b001 : node232;
								assign node232 = (inp[2]) ? node234 : 3'b011;
									assign node234 = (inp[11]) ? node236 : 3'b011;
										assign node236 = (inp[5]) ? 3'b011 : 3'b001;
							assign node240 = (inp[6]) ? node244 : node241;
								assign node241 = (inp[2]) ? 3'b001 : 3'b101;
								assign node244 = (inp[2]) ? node250 : node245;
									assign node245 = (inp[10]) ? 3'b100 : node246;
										assign node246 = (inp[5]) ? 3'b000 : 3'b100;
									assign node250 = (inp[11]) ? 3'b010 : 3'b000;
						assign node253 = (inp[7]) ? node267 : node254;
							assign node254 = (inp[6]) ? 3'b100 : node255;
								assign node255 = (inp[2]) ? node261 : node256;
									assign node256 = (inp[11]) ? 3'b001 : node257;
										assign node257 = (inp[10]) ? 3'b101 : 3'b001;
									assign node261 = (inp[11]) ? 3'b110 : node262;
										assign node262 = (inp[10]) ? 3'b001 : 3'b110;
							assign node267 = (inp[6]) ? 3'b000 : node268;
								assign node268 = (inp[2]) ? node274 : node269;
									assign node269 = (inp[8]) ? node271 : 3'b010;
										assign node271 = (inp[11]) ? 3'b010 : 3'b110;
									assign node274 = (inp[8]) ? node276 : 3'b100;
										assign node276 = (inp[11]) ? 3'b010 : 3'b100;
				assign node280 = (inp[6]) ? node324 : node281;
					assign node281 = (inp[1]) ? node283 : 3'b111;
						assign node283 = (inp[4]) ? node305 : node284;
							assign node284 = (inp[2]) ? node296 : node285;
								assign node285 = (inp[8]) ? node291 : node286;
									assign node286 = (inp[10]) ? 3'b001 : node287;
										assign node287 = (inp[7]) ? 3'b110 : 3'b010;
									assign node291 = (inp[7]) ? node293 : 3'b010;
										assign node293 = (inp[5]) ? 3'b001 : 3'b010;
								assign node296 = (inp[8]) ? node300 : node297;
									assign node297 = (inp[11]) ? 3'b101 : 3'b110;
									assign node300 = (inp[7]) ? 3'b001 : node301;
										assign node301 = (inp[10]) ? 3'b100 : 3'b010;
							assign node305 = (inp[7]) ? node313 : node306;
								assign node306 = (inp[10]) ? node308 : 3'b111;
									assign node308 = (inp[11]) ? node310 : 3'b011;
										assign node310 = (inp[2]) ? 3'b011 : 3'b111;
								assign node313 = (inp[2]) ? node319 : node314;
									assign node314 = (inp[8]) ? 3'b001 : node315;
										assign node315 = (inp[10]) ? 3'b011 : 3'b001;
									assign node319 = (inp[8]) ? 3'b101 : node320;
										assign node320 = (inp[10]) ? 3'b011 : 3'b101;
					assign node324 = (inp[1]) ? node350 : node325;
						assign node325 = (inp[7]) ? node341 : node326;
							assign node326 = (inp[4]) ? node334 : node327;
								assign node327 = (inp[10]) ? node329 : 3'b101;
									assign node329 = (inp[5]) ? 3'b001 : node330;
										assign node330 = (inp[11]) ? 3'b001 : 3'b101;
								assign node334 = (inp[2]) ? node336 : 3'b010;
									assign node336 = (inp[11]) ? node338 : 3'b101;
										assign node338 = (inp[10]) ? 3'b000 : 3'b001;
							assign node341 = (inp[4]) ? node345 : node342;
								assign node342 = (inp[2]) ? 3'b010 : 3'b110;
								assign node345 = (inp[11]) ? 3'b001 : node346;
									assign node346 = (inp[8]) ? 3'b001 : 3'b110;
						assign node350 = (inp[2]) ? node364 : node351;
							assign node351 = (inp[4]) ? node357 : node352;
								assign node352 = (inp[7]) ? 3'b100 : node353;
									assign node353 = (inp[5]) ? 3'b110 : 3'b010;
								assign node357 = (inp[7]) ? 3'b010 : node358;
									assign node358 = (inp[5]) ? 3'b000 : node359;
										assign node359 = (inp[10]) ? 3'b001 : 3'b000;
							assign node364 = (inp[7]) ? node372 : node365;
								assign node365 = (inp[10]) ? 3'b110 : node366;
									assign node366 = (inp[4]) ? 3'b010 : node367;
										assign node367 = (inp[5]) ? 3'b010 : 3'b110;
								assign node372 = (inp[8]) ? node374 : 3'b010;
									assign node374 = (inp[4]) ? node376 : 3'b000;
										assign node376 = (inp[11]) ? 3'b000 : 3'b100;

endmodule