module dtc_split75_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node11;
	wire [15-1:0] node14;
	wire [15-1:0] node15;
	wire [15-1:0] node18;
	wire [15-1:0] node21;
	wire [15-1:0] node22;
	wire [15-1:0] node23;
	wire [15-1:0] node26;
	wire [15-1:0] node29;
	wire [15-1:0] node30;
	wire [15-1:0] node33;
	wire [15-1:0] node36;
	wire [15-1:0] node37;
	wire [15-1:0] node38;
	wire [15-1:0] node39;
	wire [15-1:0] node42;
	wire [15-1:0] node45;
	wire [15-1:0] node46;
	wire [15-1:0] node49;
	wire [15-1:0] node52;
	wire [15-1:0] node53;
	wire [15-1:0] node54;
	wire [15-1:0] node57;
	wire [15-1:0] node60;
	wire [15-1:0] node61;
	wire [15-1:0] node64;
	wire [15-1:0] node67;
	wire [15-1:0] node68;
	wire [15-1:0] node69;
	wire [15-1:0] node70;
	wire [15-1:0] node71;
	wire [15-1:0] node74;
	wire [15-1:0] node77;
	wire [15-1:0] node78;
	wire [15-1:0] node81;
	wire [15-1:0] node84;
	wire [15-1:0] node85;
	wire [15-1:0] node86;
	wire [15-1:0] node89;
	wire [15-1:0] node92;
	wire [15-1:0] node93;
	wire [15-1:0] node96;
	wire [15-1:0] node99;
	wire [15-1:0] node100;
	wire [15-1:0] node101;
	wire [15-1:0] node102;
	wire [15-1:0] node105;
	wire [15-1:0] node108;
	wire [15-1:0] node109;
	wire [15-1:0] node112;
	wire [15-1:0] node115;
	wire [15-1:0] node116;
	wire [15-1:0] node117;
	wire [15-1:0] node120;
	wire [15-1:0] node123;
	wire [15-1:0] node124;
	wire [15-1:0] node127;
	wire [15-1:0] node130;
	wire [15-1:0] node131;
	wire [15-1:0] node132;
	wire [15-1:0] node133;
	wire [15-1:0] node134;
	wire [15-1:0] node135;
	wire [15-1:0] node138;
	wire [15-1:0] node141;
	wire [15-1:0] node142;
	wire [15-1:0] node145;
	wire [15-1:0] node148;
	wire [15-1:0] node149;
	wire [15-1:0] node150;
	wire [15-1:0] node153;
	wire [15-1:0] node156;
	wire [15-1:0] node157;
	wire [15-1:0] node160;
	wire [15-1:0] node163;
	wire [15-1:0] node164;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node169;
	wire [15-1:0] node172;
	wire [15-1:0] node173;
	wire [15-1:0] node176;
	wire [15-1:0] node179;
	wire [15-1:0] node180;
	wire [15-1:0] node181;
	wire [15-1:0] node184;
	wire [15-1:0] node187;
	wire [15-1:0] node188;
	wire [15-1:0] node191;
	wire [15-1:0] node194;
	wire [15-1:0] node195;
	wire [15-1:0] node196;
	wire [15-1:0] node197;
	wire [15-1:0] node198;
	wire [15-1:0] node201;
	wire [15-1:0] node204;
	wire [15-1:0] node205;
	wire [15-1:0] node208;
	wire [15-1:0] node211;
	wire [15-1:0] node212;
	wire [15-1:0] node213;
	wire [15-1:0] node216;
	wire [15-1:0] node219;
	wire [15-1:0] node220;
	wire [15-1:0] node223;
	wire [15-1:0] node226;
	wire [15-1:0] node227;
	wire [15-1:0] node228;
	wire [15-1:0] node229;
	wire [15-1:0] node232;
	wire [15-1:0] node235;
	wire [15-1:0] node236;
	wire [15-1:0] node239;
	wire [15-1:0] node242;
	wire [15-1:0] node243;
	wire [15-1:0] node244;
	wire [15-1:0] node247;
	wire [15-1:0] node250;
	wire [15-1:0] node251;
	wire [15-1:0] node254;
	wire [15-1:0] node257;
	wire [15-1:0] node258;
	wire [15-1:0] node259;
	wire [15-1:0] node260;
	wire [15-1:0] node261;
	wire [15-1:0] node262;
	wire [15-1:0] node263;
	wire [15-1:0] node266;
	wire [15-1:0] node269;
	wire [15-1:0] node270;
	wire [15-1:0] node273;
	wire [15-1:0] node276;
	wire [15-1:0] node277;
	wire [15-1:0] node278;
	wire [15-1:0] node281;
	wire [15-1:0] node284;
	wire [15-1:0] node285;
	wire [15-1:0] node288;
	wire [15-1:0] node291;
	wire [15-1:0] node292;
	wire [15-1:0] node293;
	wire [15-1:0] node294;
	wire [15-1:0] node297;
	wire [15-1:0] node300;
	wire [15-1:0] node301;
	wire [15-1:0] node304;
	wire [15-1:0] node307;
	wire [15-1:0] node308;
	wire [15-1:0] node309;
	wire [15-1:0] node312;
	wire [15-1:0] node315;
	wire [15-1:0] node316;
	wire [15-1:0] node319;
	wire [15-1:0] node322;
	wire [15-1:0] node323;
	wire [15-1:0] node324;
	wire [15-1:0] node325;
	wire [15-1:0] node326;
	wire [15-1:0] node329;
	wire [15-1:0] node332;
	wire [15-1:0] node333;
	wire [15-1:0] node336;
	wire [15-1:0] node339;
	wire [15-1:0] node340;
	wire [15-1:0] node341;
	wire [15-1:0] node344;
	wire [15-1:0] node347;
	wire [15-1:0] node348;
	wire [15-1:0] node351;
	wire [15-1:0] node354;
	wire [15-1:0] node355;
	wire [15-1:0] node356;
	wire [15-1:0] node357;
	wire [15-1:0] node360;
	wire [15-1:0] node363;
	wire [15-1:0] node364;
	wire [15-1:0] node367;
	wire [15-1:0] node370;
	wire [15-1:0] node371;
	wire [15-1:0] node372;
	wire [15-1:0] node375;
	wire [15-1:0] node378;
	wire [15-1:0] node379;
	wire [15-1:0] node382;
	wire [15-1:0] node385;
	wire [15-1:0] node386;
	wire [15-1:0] node387;
	wire [15-1:0] node388;
	wire [15-1:0] node389;
	wire [15-1:0] node390;
	wire [15-1:0] node393;
	wire [15-1:0] node396;
	wire [15-1:0] node397;
	wire [15-1:0] node400;
	wire [15-1:0] node403;
	wire [15-1:0] node404;
	wire [15-1:0] node405;
	wire [15-1:0] node408;
	wire [15-1:0] node411;
	wire [15-1:0] node412;
	wire [15-1:0] node415;
	wire [15-1:0] node418;
	wire [15-1:0] node419;
	wire [15-1:0] node420;
	wire [15-1:0] node421;
	wire [15-1:0] node424;
	wire [15-1:0] node427;
	wire [15-1:0] node428;
	wire [15-1:0] node431;
	wire [15-1:0] node434;
	wire [15-1:0] node435;
	wire [15-1:0] node436;
	wire [15-1:0] node439;
	wire [15-1:0] node442;
	wire [15-1:0] node443;
	wire [15-1:0] node446;
	wire [15-1:0] node449;
	wire [15-1:0] node450;
	wire [15-1:0] node451;
	wire [15-1:0] node452;
	wire [15-1:0] node453;
	wire [15-1:0] node456;
	wire [15-1:0] node459;
	wire [15-1:0] node460;
	wire [15-1:0] node463;
	wire [15-1:0] node466;
	wire [15-1:0] node467;
	wire [15-1:0] node468;
	wire [15-1:0] node471;
	wire [15-1:0] node474;
	wire [15-1:0] node475;
	wire [15-1:0] node478;
	wire [15-1:0] node481;
	wire [15-1:0] node482;
	wire [15-1:0] node483;
	wire [15-1:0] node484;
	wire [15-1:0] node487;
	wire [15-1:0] node490;
	wire [15-1:0] node491;
	wire [15-1:0] node494;
	wire [15-1:0] node497;
	wire [15-1:0] node498;
	wire [15-1:0] node499;
	wire [15-1:0] node502;
	wire [15-1:0] node505;
	wire [15-1:0] node506;
	wire [15-1:0] node509;
	wire [15-1:0] node512;
	wire [15-1:0] node513;
	wire [15-1:0] node514;
	wire [15-1:0] node515;
	wire [15-1:0] node516;
	wire [15-1:0] node517;
	wire [15-1:0] node518;
	wire [15-1:0] node519;
	wire [15-1:0] node522;
	wire [15-1:0] node525;
	wire [15-1:0] node526;
	wire [15-1:0] node529;
	wire [15-1:0] node532;
	wire [15-1:0] node533;
	wire [15-1:0] node534;
	wire [15-1:0] node537;
	wire [15-1:0] node540;
	wire [15-1:0] node541;
	wire [15-1:0] node544;
	wire [15-1:0] node547;
	wire [15-1:0] node548;
	wire [15-1:0] node549;
	wire [15-1:0] node550;
	wire [15-1:0] node553;
	wire [15-1:0] node556;
	wire [15-1:0] node557;
	wire [15-1:0] node560;
	wire [15-1:0] node563;
	wire [15-1:0] node564;
	wire [15-1:0] node565;
	wire [15-1:0] node568;
	wire [15-1:0] node571;
	wire [15-1:0] node572;
	wire [15-1:0] node575;
	wire [15-1:0] node578;
	wire [15-1:0] node579;
	wire [15-1:0] node580;
	wire [15-1:0] node581;
	wire [15-1:0] node582;
	wire [15-1:0] node585;
	wire [15-1:0] node588;
	wire [15-1:0] node589;
	wire [15-1:0] node592;
	wire [15-1:0] node595;
	wire [15-1:0] node596;
	wire [15-1:0] node597;
	wire [15-1:0] node600;
	wire [15-1:0] node603;
	wire [15-1:0] node604;
	wire [15-1:0] node607;
	wire [15-1:0] node610;
	wire [15-1:0] node611;
	wire [15-1:0] node612;
	wire [15-1:0] node613;
	wire [15-1:0] node616;
	wire [15-1:0] node619;
	wire [15-1:0] node620;
	wire [15-1:0] node623;
	wire [15-1:0] node626;
	wire [15-1:0] node627;
	wire [15-1:0] node628;
	wire [15-1:0] node631;
	wire [15-1:0] node634;
	wire [15-1:0] node635;
	wire [15-1:0] node638;
	wire [15-1:0] node641;
	wire [15-1:0] node642;
	wire [15-1:0] node643;
	wire [15-1:0] node644;
	wire [15-1:0] node645;
	wire [15-1:0] node646;
	wire [15-1:0] node649;
	wire [15-1:0] node652;
	wire [15-1:0] node653;
	wire [15-1:0] node656;
	wire [15-1:0] node659;
	wire [15-1:0] node660;
	wire [15-1:0] node661;
	wire [15-1:0] node664;
	wire [15-1:0] node667;
	wire [15-1:0] node668;
	wire [15-1:0] node671;
	wire [15-1:0] node674;
	wire [15-1:0] node675;
	wire [15-1:0] node676;
	wire [15-1:0] node677;
	wire [15-1:0] node680;
	wire [15-1:0] node683;
	wire [15-1:0] node684;
	wire [15-1:0] node687;
	wire [15-1:0] node690;
	wire [15-1:0] node691;
	wire [15-1:0] node692;
	wire [15-1:0] node695;
	wire [15-1:0] node698;
	wire [15-1:0] node699;
	wire [15-1:0] node702;
	wire [15-1:0] node705;
	wire [15-1:0] node706;
	wire [15-1:0] node707;
	wire [15-1:0] node708;
	wire [15-1:0] node709;
	wire [15-1:0] node712;
	wire [15-1:0] node715;
	wire [15-1:0] node716;
	wire [15-1:0] node719;
	wire [15-1:0] node722;
	wire [15-1:0] node723;
	wire [15-1:0] node724;
	wire [15-1:0] node727;
	wire [15-1:0] node730;
	wire [15-1:0] node731;
	wire [15-1:0] node734;
	wire [15-1:0] node737;
	wire [15-1:0] node738;
	wire [15-1:0] node739;
	wire [15-1:0] node740;
	wire [15-1:0] node743;
	wire [15-1:0] node746;
	wire [15-1:0] node747;
	wire [15-1:0] node750;
	wire [15-1:0] node753;
	wire [15-1:0] node754;
	wire [15-1:0] node755;
	wire [15-1:0] node758;
	wire [15-1:0] node761;
	wire [15-1:0] node762;
	wire [15-1:0] node765;
	wire [15-1:0] node768;
	wire [15-1:0] node769;
	wire [15-1:0] node770;
	wire [15-1:0] node771;
	wire [15-1:0] node772;
	wire [15-1:0] node773;
	wire [15-1:0] node774;
	wire [15-1:0] node777;
	wire [15-1:0] node780;
	wire [15-1:0] node781;
	wire [15-1:0] node784;
	wire [15-1:0] node787;
	wire [15-1:0] node788;
	wire [15-1:0] node789;
	wire [15-1:0] node792;
	wire [15-1:0] node795;
	wire [15-1:0] node796;
	wire [15-1:0] node799;
	wire [15-1:0] node802;
	wire [15-1:0] node803;
	wire [15-1:0] node804;
	wire [15-1:0] node805;
	wire [15-1:0] node808;
	wire [15-1:0] node811;
	wire [15-1:0] node812;
	wire [15-1:0] node815;
	wire [15-1:0] node818;
	wire [15-1:0] node819;
	wire [15-1:0] node820;
	wire [15-1:0] node823;
	wire [15-1:0] node826;
	wire [15-1:0] node827;
	wire [15-1:0] node830;
	wire [15-1:0] node833;
	wire [15-1:0] node834;
	wire [15-1:0] node835;
	wire [15-1:0] node836;
	wire [15-1:0] node837;
	wire [15-1:0] node840;
	wire [15-1:0] node843;
	wire [15-1:0] node844;
	wire [15-1:0] node847;
	wire [15-1:0] node850;
	wire [15-1:0] node851;
	wire [15-1:0] node852;
	wire [15-1:0] node855;
	wire [15-1:0] node858;
	wire [15-1:0] node859;
	wire [15-1:0] node862;
	wire [15-1:0] node865;
	wire [15-1:0] node866;
	wire [15-1:0] node867;
	wire [15-1:0] node868;
	wire [15-1:0] node871;
	wire [15-1:0] node874;
	wire [15-1:0] node875;
	wire [15-1:0] node878;
	wire [15-1:0] node881;
	wire [15-1:0] node882;
	wire [15-1:0] node883;
	wire [15-1:0] node886;
	wire [15-1:0] node889;
	wire [15-1:0] node890;
	wire [15-1:0] node893;
	wire [15-1:0] node896;
	wire [15-1:0] node897;
	wire [15-1:0] node898;
	wire [15-1:0] node899;
	wire [15-1:0] node900;
	wire [15-1:0] node901;
	wire [15-1:0] node904;
	wire [15-1:0] node907;
	wire [15-1:0] node908;
	wire [15-1:0] node911;
	wire [15-1:0] node914;
	wire [15-1:0] node915;
	wire [15-1:0] node916;
	wire [15-1:0] node919;
	wire [15-1:0] node922;
	wire [15-1:0] node923;
	wire [15-1:0] node926;
	wire [15-1:0] node929;
	wire [15-1:0] node930;
	wire [15-1:0] node931;
	wire [15-1:0] node932;
	wire [15-1:0] node935;
	wire [15-1:0] node938;
	wire [15-1:0] node939;
	wire [15-1:0] node942;
	wire [15-1:0] node945;
	wire [15-1:0] node946;
	wire [15-1:0] node947;
	wire [15-1:0] node950;
	wire [15-1:0] node953;
	wire [15-1:0] node954;
	wire [15-1:0] node957;
	wire [15-1:0] node960;
	wire [15-1:0] node961;
	wire [15-1:0] node962;
	wire [15-1:0] node963;
	wire [15-1:0] node964;
	wire [15-1:0] node967;
	wire [15-1:0] node970;
	wire [15-1:0] node971;
	wire [15-1:0] node974;
	wire [15-1:0] node977;
	wire [15-1:0] node978;
	wire [15-1:0] node979;
	wire [15-1:0] node982;
	wire [15-1:0] node985;
	wire [15-1:0] node986;
	wire [15-1:0] node989;
	wire [15-1:0] node992;
	wire [15-1:0] node993;
	wire [15-1:0] node994;
	wire [15-1:0] node995;
	wire [15-1:0] node998;
	wire [15-1:0] node1001;
	wire [15-1:0] node1002;
	wire [15-1:0] node1005;
	wire [15-1:0] node1008;
	wire [15-1:0] node1009;
	wire [15-1:0] node1010;
	wire [15-1:0] node1013;
	wire [15-1:0] node1016;
	wire [15-1:0] node1017;
	wire [15-1:0] node1020;

	assign outp = (inp[4]) ? node512 : node1;
		assign node1 = (inp[9]) ? node257 : node2;
			assign node2 = (inp[7]) ? node130 : node3;
				assign node3 = (inp[13]) ? node67 : node4;
					assign node4 = (inp[11]) ? node36 : node5;
						assign node5 = (inp[12]) ? node21 : node6;
							assign node6 = (inp[0]) ? node14 : node7;
								assign node7 = (inp[14]) ? node11 : node8;
									assign node8 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
									assign node11 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
								assign node14 = (inp[6]) ? node18 : node15;
									assign node15 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node18 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node21 = (inp[2]) ? node29 : node22;
								assign node22 = (inp[6]) ? node26 : node23;
									assign node23 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node26 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node29 = (inp[0]) ? node33 : node30;
									assign node30 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node33 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node36 = (inp[10]) ? node52 : node37;
							assign node37 = (inp[8]) ? node45 : node38;
								assign node38 = (inp[6]) ? node42 : node39;
									assign node39 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node42 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node45 = (inp[3]) ? node49 : node46;
									assign node46 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node49 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node52 = (inp[5]) ? node60 : node53;
								assign node53 = (inp[3]) ? node57 : node54;
									assign node54 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node57 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node60 = (inp[12]) ? node64 : node61;
									assign node61 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node64 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
					assign node67 = (inp[3]) ? node99 : node68;
						assign node68 = (inp[2]) ? node84 : node69;
							assign node69 = (inp[6]) ? node77 : node70;
								assign node70 = (inp[1]) ? node74 : node71;
									assign node71 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node74 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node77 = (inp[14]) ? node81 : node78;
									assign node78 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node81 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node84 = (inp[8]) ? node92 : node85;
								assign node85 = (inp[0]) ? node89 : node86;
									assign node86 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node89 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node92 = (inp[12]) ? node96 : node93;
									assign node93 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node96 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node99 = (inp[8]) ? node115 : node100;
							assign node100 = (inp[0]) ? node108 : node101;
								assign node101 = (inp[14]) ? node105 : node102;
									assign node102 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node105 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node108 = (inp[11]) ? node112 : node109;
									assign node109 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node112 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node115 = (inp[1]) ? node123 : node116;
								assign node116 = (inp[12]) ? node120 : node117;
									assign node117 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node120 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node123 = (inp[12]) ? node127 : node124;
									assign node124 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node127 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
				assign node130 = (inp[5]) ? node194 : node131;
					assign node131 = (inp[14]) ? node163 : node132;
						assign node132 = (inp[11]) ? node148 : node133;
							assign node133 = (inp[2]) ? node141 : node134;
								assign node134 = (inp[10]) ? node138 : node135;
									assign node135 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node138 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node141 = (inp[0]) ? node145 : node142;
									assign node142 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node145 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node148 = (inp[6]) ? node156 : node149;
								assign node149 = (inp[3]) ? node153 : node150;
									assign node150 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node153 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node156 = (inp[12]) ? node160 : node157;
									assign node157 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node160 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node163 = (inp[12]) ? node179 : node164;
							assign node164 = (inp[2]) ? node172 : node165;
								assign node165 = (inp[3]) ? node169 : node166;
									assign node166 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node169 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node172 = (inp[6]) ? node176 : node173;
									assign node173 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node176 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node179 = (inp[13]) ? node187 : node180;
								assign node180 = (inp[8]) ? node184 : node181;
									assign node181 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node184 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node187 = (inp[11]) ? node191 : node188;
									assign node188 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node191 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node194 = (inp[2]) ? node226 : node195;
						assign node195 = (inp[3]) ? node211 : node196;
							assign node196 = (inp[1]) ? node204 : node197;
								assign node197 = (inp[14]) ? node201 : node198;
									assign node198 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node201 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node204 = (inp[13]) ? node208 : node205;
									assign node205 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node208 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node211 = (inp[12]) ? node219 : node212;
								assign node212 = (inp[11]) ? node216 : node213;
									assign node213 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node216 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node219 = (inp[6]) ? node223 : node220;
									assign node220 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node223 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node226 = (inp[3]) ? node242 : node227;
							assign node227 = (inp[6]) ? node235 : node228;
								assign node228 = (inp[11]) ? node232 : node229;
									assign node229 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node232 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node235 = (inp[12]) ? node239 : node236;
									assign node236 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node239 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node242 = (inp[12]) ? node250 : node243;
								assign node243 = (inp[14]) ? node247 : node244;
									assign node244 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node247 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node250 = (inp[13]) ? node254 : node251;
									assign node251 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node254 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
			assign node257 = (inp[1]) ? node385 : node258;
				assign node258 = (inp[3]) ? node322 : node259;
					assign node259 = (inp[7]) ? node291 : node260;
						assign node260 = (inp[13]) ? node276 : node261;
							assign node261 = (inp[11]) ? node269 : node262;
								assign node262 = (inp[6]) ? node266 : node263;
									assign node263 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node266 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node269 = (inp[12]) ? node273 : node270;
									assign node270 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node273 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node276 = (inp[5]) ? node284 : node277;
								assign node277 = (inp[2]) ? node281 : node278;
									assign node278 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node281 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node284 = (inp[8]) ? node288 : node285;
									assign node285 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node288 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node291 = (inp[0]) ? node307 : node292;
							assign node292 = (inp[2]) ? node300 : node293;
								assign node293 = (inp[6]) ? node297 : node294;
									assign node294 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node297 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node300 = (inp[12]) ? node304 : node301;
									assign node301 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node304 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node307 = (inp[8]) ? node315 : node308;
								assign node308 = (inp[5]) ? node312 : node309;
									assign node309 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node312 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node315 = (inp[5]) ? node319 : node316;
									assign node316 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node319 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node322 = (inp[14]) ? node354 : node323;
						assign node323 = (inp[12]) ? node339 : node324;
							assign node324 = (inp[10]) ? node332 : node325;
								assign node325 = (inp[2]) ? node329 : node326;
									assign node326 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node329 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node332 = (inp[13]) ? node336 : node333;
									assign node333 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node336 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node339 = (inp[8]) ? node347 : node340;
								assign node340 = (inp[10]) ? node344 : node341;
									assign node341 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node344 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node347 = (inp[0]) ? node351 : node348;
									assign node348 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node351 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node354 = (inp[11]) ? node370 : node355;
							assign node355 = (inp[0]) ? node363 : node356;
								assign node356 = (inp[10]) ? node360 : node357;
									assign node357 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node360 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node363 = (inp[12]) ? node367 : node364;
									assign node364 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node367 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node370 = (inp[8]) ? node378 : node371;
								assign node371 = (inp[6]) ? node375 : node372;
									assign node372 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node375 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node378 = (inp[12]) ? node382 : node379;
									assign node379 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node382 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
				assign node385 = (inp[14]) ? node449 : node386;
					assign node386 = (inp[11]) ? node418 : node387;
						assign node387 = (inp[6]) ? node403 : node388;
							assign node388 = (inp[5]) ? node396 : node389;
								assign node389 = (inp[7]) ? node393 : node390;
									assign node390 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node393 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node396 = (inp[3]) ? node400 : node397;
									assign node397 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node400 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node403 = (inp[13]) ? node411 : node404;
								assign node404 = (inp[12]) ? node408 : node405;
									assign node405 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node408 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node411 = (inp[3]) ? node415 : node412;
									assign node412 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node415 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node418 = (inp[5]) ? node434 : node419;
							assign node419 = (inp[7]) ? node427 : node420;
								assign node420 = (inp[10]) ? node424 : node421;
									assign node421 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node424 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node427 = (inp[12]) ? node431 : node428;
									assign node428 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node431 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node434 = (inp[8]) ? node442 : node435;
								assign node435 = (inp[7]) ? node439 : node436;
									assign node436 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node439 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node442 = (inp[0]) ? node446 : node443;
									assign node443 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node446 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node449 = (inp[3]) ? node481 : node450;
						assign node450 = (inp[12]) ? node466 : node451;
							assign node451 = (inp[11]) ? node459 : node452;
								assign node452 = (inp[0]) ? node456 : node453;
									assign node453 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node456 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node459 = (inp[7]) ? node463 : node460;
									assign node460 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node463 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node466 = (inp[10]) ? node474 : node467;
								assign node467 = (inp[2]) ? node471 : node468;
									assign node468 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node471 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node474 = (inp[7]) ? node478 : node475;
									assign node475 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node478 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node481 = (inp[5]) ? node497 : node482;
							assign node482 = (inp[11]) ? node490 : node483;
								assign node483 = (inp[2]) ? node487 : node484;
									assign node484 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node487 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node490 = (inp[0]) ? node494 : node491;
									assign node491 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node494 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node497 = (inp[10]) ? node505 : node498;
								assign node498 = (inp[8]) ? node502 : node499;
									assign node499 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node502 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node505 = (inp[6]) ? node509 : node506;
									assign node506 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node509 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
		assign node512 = (inp[8]) ? node768 : node513;
			assign node513 = (inp[13]) ? node641 : node514;
				assign node514 = (inp[3]) ? node578 : node515;
					assign node515 = (inp[9]) ? node547 : node516;
						assign node516 = (inp[6]) ? node532 : node517;
							assign node517 = (inp[5]) ? node525 : node518;
								assign node518 = (inp[2]) ? node522 : node519;
									assign node519 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node522 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node525 = (inp[12]) ? node529 : node526;
									assign node526 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node529 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node532 = (inp[1]) ? node540 : node533;
								assign node533 = (inp[5]) ? node537 : node534;
									assign node534 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node537 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node540 = (inp[11]) ? node544 : node541;
									assign node541 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node544 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node547 = (inp[2]) ? node563 : node548;
							assign node548 = (inp[12]) ? node556 : node549;
								assign node549 = (inp[11]) ? node553 : node550;
									assign node550 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node553 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node556 = (inp[0]) ? node560 : node557;
									assign node557 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node560 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node563 = (inp[7]) ? node571 : node564;
								assign node564 = (inp[11]) ? node568 : node565;
									assign node565 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node568 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node571 = (inp[6]) ? node575 : node572;
									assign node572 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node575 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node578 = (inp[1]) ? node610 : node579;
						assign node579 = (inp[5]) ? node595 : node580;
							assign node580 = (inp[2]) ? node588 : node581;
								assign node581 = (inp[11]) ? node585 : node582;
									assign node582 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node585 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node588 = (inp[12]) ? node592 : node589;
									assign node589 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node592 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node595 = (inp[6]) ? node603 : node596;
								assign node596 = (inp[2]) ? node600 : node597;
									assign node597 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node600 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node603 = (inp[0]) ? node607 : node604;
									assign node604 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node607 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node610 = (inp[11]) ? node626 : node611;
							assign node611 = (inp[0]) ? node619 : node612;
								assign node612 = (inp[6]) ? node616 : node613;
									assign node613 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node616 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node619 = (inp[12]) ? node623 : node620;
									assign node620 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node623 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node626 = (inp[2]) ? node634 : node627;
								assign node627 = (inp[6]) ? node631 : node628;
									assign node628 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node631 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node634 = (inp[7]) ? node638 : node635;
									assign node635 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node638 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
				assign node641 = (inp[10]) ? node705 : node642;
					assign node642 = (inp[1]) ? node674 : node643;
						assign node643 = (inp[5]) ? node659 : node644;
							assign node644 = (inp[9]) ? node652 : node645;
								assign node645 = (inp[14]) ? node649 : node646;
									assign node646 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node649 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node652 = (inp[0]) ? node656 : node653;
									assign node653 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node656 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node659 = (inp[11]) ? node667 : node660;
								assign node660 = (inp[7]) ? node664 : node661;
									assign node661 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node664 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node667 = (inp[2]) ? node671 : node668;
									assign node668 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node671 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node674 = (inp[12]) ? node690 : node675;
							assign node675 = (inp[3]) ? node683 : node676;
								assign node676 = (inp[9]) ? node680 : node677;
									assign node677 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node680 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node683 = (inp[0]) ? node687 : node684;
									assign node684 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node687 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node690 = (inp[11]) ? node698 : node691;
								assign node691 = (inp[0]) ? node695 : node692;
									assign node692 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node695 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node698 = (inp[9]) ? node702 : node699;
									assign node699 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node702 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node705 = (inp[9]) ? node737 : node706;
						assign node706 = (inp[11]) ? node722 : node707;
							assign node707 = (inp[7]) ? node715 : node708;
								assign node708 = (inp[2]) ? node712 : node709;
									assign node709 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node712 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node715 = (inp[1]) ? node719 : node716;
									assign node716 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node719 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node722 = (inp[6]) ? node730 : node723;
								assign node723 = (inp[5]) ? node727 : node724;
									assign node724 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node727 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node730 = (inp[14]) ? node734 : node731;
									assign node731 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node734 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node737 = (inp[0]) ? node753 : node738;
							assign node738 = (inp[14]) ? node746 : node739;
								assign node739 = (inp[11]) ? node743 : node740;
									assign node740 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node743 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node746 = (inp[7]) ? node750 : node747;
									assign node747 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node750 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node753 = (inp[11]) ? node761 : node754;
								assign node754 = (inp[3]) ? node758 : node755;
									assign node755 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node758 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node761 = (inp[14]) ? node765 : node762;
									assign node762 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node765 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
			assign node768 = (inp[11]) ? node896 : node769;
				assign node769 = (inp[7]) ? node833 : node770;
					assign node770 = (inp[1]) ? node802 : node771;
						assign node771 = (inp[0]) ? node787 : node772;
							assign node772 = (inp[3]) ? node780 : node773;
								assign node773 = (inp[13]) ? node777 : node774;
									assign node774 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node777 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node780 = (inp[2]) ? node784 : node781;
									assign node781 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node784 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node787 = (inp[6]) ? node795 : node788;
								assign node788 = (inp[9]) ? node792 : node789;
									assign node789 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node792 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node795 = (inp[14]) ? node799 : node796;
									assign node796 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node799 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node802 = (inp[14]) ? node818 : node803;
							assign node803 = (inp[13]) ? node811 : node804;
								assign node804 = (inp[6]) ? node808 : node805;
									assign node805 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node808 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node811 = (inp[6]) ? node815 : node812;
									assign node812 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node815 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node818 = (inp[6]) ? node826 : node819;
								assign node819 = (inp[12]) ? node823 : node820;
									assign node820 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node823 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node826 = (inp[12]) ? node830 : node827;
									assign node827 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node830 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node833 = (inp[6]) ? node865 : node834;
						assign node834 = (inp[13]) ? node850 : node835;
							assign node835 = (inp[1]) ? node843 : node836;
								assign node836 = (inp[12]) ? node840 : node837;
									assign node837 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node840 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node843 = (inp[2]) ? node847 : node844;
									assign node844 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node847 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node850 = (inp[0]) ? node858 : node851;
								assign node851 = (inp[2]) ? node855 : node852;
									assign node852 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node855 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node858 = (inp[9]) ? node862 : node859;
									assign node859 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node862 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node865 = (inp[3]) ? node881 : node866;
							assign node866 = (inp[1]) ? node874 : node867;
								assign node867 = (inp[12]) ? node871 : node868;
									assign node868 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node871 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node874 = (inp[9]) ? node878 : node875;
									assign node875 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node878 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node881 = (inp[0]) ? node889 : node882;
								assign node882 = (inp[2]) ? node886 : node883;
									assign node883 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node886 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node889 = (inp[13]) ? node893 : node890;
									assign node890 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node893 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node896 = (inp[6]) ? node960 : node897;
					assign node897 = (inp[13]) ? node929 : node898;
						assign node898 = (inp[14]) ? node914 : node899;
							assign node899 = (inp[2]) ? node907 : node900;
								assign node900 = (inp[9]) ? node904 : node901;
									assign node901 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node904 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node907 = (inp[5]) ? node911 : node908;
									assign node908 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node911 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node914 = (inp[3]) ? node922 : node915;
								assign node915 = (inp[2]) ? node919 : node916;
									assign node916 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node919 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node922 = (inp[0]) ? node926 : node923;
									assign node923 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node926 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node929 = (inp[5]) ? node945 : node930;
							assign node930 = (inp[10]) ? node938 : node931;
								assign node931 = (inp[7]) ? node935 : node932;
									assign node932 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node935 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node938 = (inp[9]) ? node942 : node939;
									assign node939 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node942 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node945 = (inp[7]) ? node953 : node946;
								assign node946 = (inp[10]) ? node950 : node947;
									assign node947 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node950 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node953 = (inp[1]) ? node957 : node954;
									assign node954 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node957 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node960 = (inp[12]) ? node992 : node961;
						assign node961 = (inp[0]) ? node977 : node962;
							assign node962 = (inp[9]) ? node970 : node963;
								assign node963 = (inp[3]) ? node967 : node964;
									assign node964 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node967 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node970 = (inp[7]) ? node974 : node971;
									assign node971 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node974 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node977 = (inp[14]) ? node985 : node978;
								assign node978 = (inp[3]) ? node982 : node979;
									assign node979 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node982 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node985 = (inp[7]) ? node989 : node986;
									assign node986 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node989 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node992 = (inp[7]) ? node1008 : node993;
							assign node993 = (inp[0]) ? node1001 : node994;
								assign node994 = (inp[5]) ? node998 : node995;
									assign node995 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node998 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1001 = (inp[10]) ? node1005 : node1002;
									assign node1002 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1005 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node1008 = (inp[9]) ? node1016 : node1009;
								assign node1009 = (inp[1]) ? node1013 : node1010;
									assign node1010 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1013 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1016 = (inp[2]) ? node1020 : node1017;
									assign node1017 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node1020 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;

endmodule