module dtc_split25_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node8;
	wire [13-1:0] node9;
	wire [13-1:0] node10;
	wire [13-1:0] node14;
	wire [13-1:0] node15;
	wire [13-1:0] node18;
	wire [13-1:0] node21;
	wire [13-1:0] node22;
	wire [13-1:0] node23;
	wire [13-1:0] node26;
	wire [13-1:0] node29;
	wire [13-1:0] node30;
	wire [13-1:0] node34;
	wire [13-1:0] node35;
	wire [13-1:0] node36;
	wire [13-1:0] node37;
	wire [13-1:0] node41;
	wire [13-1:0] node43;
	wire [13-1:0] node46;
	wire [13-1:0] node47;
	wire [13-1:0] node48;
	wire [13-1:0] node51;
	wire [13-1:0] node54;
	wire [13-1:0] node57;
	wire [13-1:0] node58;
	wire [13-1:0] node59;
	wire [13-1:0] node60;
	wire [13-1:0] node61;
	wire [13-1:0] node65;
	wire [13-1:0] node66;
	wire [13-1:0] node69;
	wire [13-1:0] node72;
	wire [13-1:0] node73;
	wire [13-1:0] node76;
	wire [13-1:0] node77;
	wire [13-1:0] node80;
	wire [13-1:0] node83;
	wire [13-1:0] node84;
	wire [13-1:0] node85;
	wire [13-1:0] node87;
	wire [13-1:0] node91;
	wire [13-1:0] node92;
	wire [13-1:0] node93;
	wire [13-1:0] node97;
	wire [13-1:0] node100;
	wire [13-1:0] node101;
	wire [13-1:0] node102;
	wire [13-1:0] node103;
	wire [13-1:0] node104;
	wire [13-1:0] node106;
	wire [13-1:0] node109;
	wire [13-1:0] node110;
	wire [13-1:0] node114;
	wire [13-1:0] node115;
	wire [13-1:0] node116;
	wire [13-1:0] node119;
	wire [13-1:0] node122;
	wire [13-1:0] node125;
	wire [13-1:0] node126;
	wire [13-1:0] node128;
	wire [13-1:0] node131;
	wire [13-1:0] node132;
	wire [13-1:0] node133;
	wire [13-1:0] node136;
	wire [13-1:0] node139;
	wire [13-1:0] node140;
	wire [13-1:0] node143;
	wire [13-1:0] node146;
	wire [13-1:0] node147;
	wire [13-1:0] node148;
	wire [13-1:0] node149;
	wire [13-1:0] node151;
	wire [13-1:0] node155;
	wire [13-1:0] node157;
	wire [13-1:0] node160;
	wire [13-1:0] node161;
	wire [13-1:0] node162;
	wire [13-1:0] node164;
	wire [13-1:0] node168;
	wire [13-1:0] node170;
	wire [13-1:0] node173;
	wire [13-1:0] node174;
	wire [13-1:0] node175;
	wire [13-1:0] node176;
	wire [13-1:0] node177;
	wire [13-1:0] node178;
	wire [13-1:0] node179;
	wire [13-1:0] node182;
	wire [13-1:0] node185;
	wire [13-1:0] node186;
	wire [13-1:0] node189;
	wire [13-1:0] node192;
	wire [13-1:0] node193;
	wire [13-1:0] node194;
	wire [13-1:0] node198;
	wire [13-1:0] node199;
	wire [13-1:0] node202;
	wire [13-1:0] node205;
	wire [13-1:0] node206;
	wire [13-1:0] node208;
	wire [13-1:0] node211;
	wire [13-1:0] node212;
	wire [13-1:0] node213;
	wire [13-1:0] node216;
	wire [13-1:0] node219;
	wire [13-1:0] node220;
	wire [13-1:0] node224;
	wire [13-1:0] node225;
	wire [13-1:0] node226;
	wire [13-1:0] node227;
	wire [13-1:0] node228;
	wire [13-1:0] node232;
	wire [13-1:0] node233;
	wire [13-1:0] node237;
	wire [13-1:0] node238;
	wire [13-1:0] node239;
	wire [13-1:0] node243;
	wire [13-1:0] node245;
	wire [13-1:0] node248;
	wire [13-1:0] node249;
	wire [13-1:0] node251;
	wire [13-1:0] node252;
	wire [13-1:0] node255;
	wire [13-1:0] node258;
	wire [13-1:0] node259;
	wire [13-1:0] node260;
	wire [13-1:0] node264;
	wire [13-1:0] node266;
	wire [13-1:0] node269;
	wire [13-1:0] node270;
	wire [13-1:0] node271;
	wire [13-1:0] node272;
	wire [13-1:0] node273;
	wire [13-1:0] node276;
	wire [13-1:0] node278;
	wire [13-1:0] node281;
	wire [13-1:0] node282;
	wire [13-1:0] node284;
	wire [13-1:0] node288;
	wire [13-1:0] node289;
	wire [13-1:0] node291;
	wire [13-1:0] node292;
	wire [13-1:0] node295;
	wire [13-1:0] node298;
	wire [13-1:0] node299;
	wire [13-1:0] node300;
	wire [13-1:0] node304;
	wire [13-1:0] node306;
	wire [13-1:0] node309;
	wire [13-1:0] node310;
	wire [13-1:0] node311;
	wire [13-1:0] node312;
	wire [13-1:0] node315;
	wire [13-1:0] node316;
	wire [13-1:0] node319;
	wire [13-1:0] node322;
	wire [13-1:0] node323;
	wire [13-1:0] node324;
	wire [13-1:0] node328;
	wire [13-1:0] node329;
	wire [13-1:0] node332;
	wire [13-1:0] node335;
	wire [13-1:0] node336;
	wire [13-1:0] node337;
	wire [13-1:0] node338;
	wire [13-1:0] node342;
	wire [13-1:0] node344;
	wire [13-1:0] node347;
	wire [13-1:0] node348;
	wire [13-1:0] node352;
	wire [13-1:0] node353;
	wire [13-1:0] node354;
	wire [13-1:0] node355;
	wire [13-1:0] node356;
	wire [13-1:0] node357;
	wire [13-1:0] node358;
	wire [13-1:0] node359;
	wire [13-1:0] node363;
	wire [13-1:0] node364;
	wire [13-1:0] node367;
	wire [13-1:0] node370;
	wire [13-1:0] node371;
	wire [13-1:0] node372;
	wire [13-1:0] node375;
	wire [13-1:0] node378;
	wire [13-1:0] node379;
	wire [13-1:0] node383;
	wire [13-1:0] node384;
	wire [13-1:0] node385;
	wire [13-1:0] node386;
	wire [13-1:0] node391;
	wire [13-1:0] node392;
	wire [13-1:0] node395;
	wire [13-1:0] node396;
	wire [13-1:0] node400;
	wire [13-1:0] node401;
	wire [13-1:0] node402;
	wire [13-1:0] node403;
	wire [13-1:0] node406;
	wire [13-1:0] node409;
	wire [13-1:0] node410;
	wire [13-1:0] node412;
	wire [13-1:0] node416;
	wire [13-1:0] node417;
	wire [13-1:0] node419;
	wire [13-1:0] node420;
	wire [13-1:0] node423;
	wire [13-1:0] node426;
	wire [13-1:0] node427;
	wire [13-1:0] node429;
	wire [13-1:0] node432;
	wire [13-1:0] node434;
	wire [13-1:0] node437;
	wire [13-1:0] node438;
	wire [13-1:0] node439;
	wire [13-1:0] node440;
	wire [13-1:0] node441;
	wire [13-1:0] node444;
	wire [13-1:0] node445;
	wire [13-1:0] node448;
	wire [13-1:0] node451;
	wire [13-1:0] node452;
	wire [13-1:0] node454;
	wire [13-1:0] node458;
	wire [13-1:0] node459;
	wire [13-1:0] node460;
	wire [13-1:0] node462;
	wire [13-1:0] node465;
	wire [13-1:0] node466;
	wire [13-1:0] node469;
	wire [13-1:0] node472;
	wire [13-1:0] node474;
	wire [13-1:0] node475;
	wire [13-1:0] node479;
	wire [13-1:0] node480;
	wire [13-1:0] node481;
	wire [13-1:0] node482;
	wire [13-1:0] node483;
	wire [13-1:0] node486;
	wire [13-1:0] node489;
	wire [13-1:0] node490;
	wire [13-1:0] node493;
	wire [13-1:0] node496;
	wire [13-1:0] node497;
	wire [13-1:0] node498;
	wire [13-1:0] node501;
	wire [13-1:0] node504;
	wire [13-1:0] node505;
	wire [13-1:0] node509;
	wire [13-1:0] node510;
	wire [13-1:0] node511;
	wire [13-1:0] node512;
	wire [13-1:0] node515;
	wire [13-1:0] node518;
	wire [13-1:0] node521;
	wire [13-1:0] node522;
	wire [13-1:0] node525;
	wire [13-1:0] node526;
	wire [13-1:0] node529;
	wire [13-1:0] node532;
	wire [13-1:0] node533;
	wire [13-1:0] node534;
	wire [13-1:0] node535;
	wire [13-1:0] node536;
	wire [13-1:0] node537;
	wire [13-1:0] node538;
	wire [13-1:0] node543;
	wire [13-1:0] node544;
	wire [13-1:0] node545;
	wire [13-1:0] node550;
	wire [13-1:0] node551;
	wire [13-1:0] node552;
	wire [13-1:0] node554;
	wire [13-1:0] node557;
	wire [13-1:0] node560;
	wire [13-1:0] node562;
	wire [13-1:0] node563;
	wire [13-1:0] node567;
	wire [13-1:0] node568;
	wire [13-1:0] node569;
	wire [13-1:0] node570;
	wire [13-1:0] node572;
	wire [13-1:0] node575;
	wire [13-1:0] node576;
	wire [13-1:0] node579;
	wire [13-1:0] node582;
	wire [13-1:0] node583;
	wire [13-1:0] node584;
	wire [13-1:0] node589;
	wire [13-1:0] node590;
	wire [13-1:0] node591;
	wire [13-1:0] node592;
	wire [13-1:0] node596;
	wire [13-1:0] node597;
	wire [13-1:0] node601;
	wire [13-1:0] node602;
	wire [13-1:0] node604;
	wire [13-1:0] node607;
	wire [13-1:0] node610;
	wire [13-1:0] node611;
	wire [13-1:0] node612;
	wire [13-1:0] node613;
	wire [13-1:0] node614;
	wire [13-1:0] node616;
	wire [13-1:0] node620;
	wire [13-1:0] node622;
	wire [13-1:0] node623;
	wire [13-1:0] node627;
	wire [13-1:0] node628;
	wire [13-1:0] node629;
	wire [13-1:0] node631;
	wire [13-1:0] node634;
	wire [13-1:0] node635;
	wire [13-1:0] node639;
	wire [13-1:0] node640;
	wire [13-1:0] node641;
	wire [13-1:0] node646;
	wire [13-1:0] node647;
	wire [13-1:0] node648;
	wire [13-1:0] node650;
	wire [13-1:0] node651;
	wire [13-1:0] node655;
	wire [13-1:0] node657;
	wire [13-1:0] node658;
	wire [13-1:0] node662;
	wire [13-1:0] node663;
	wire [13-1:0] node665;
	wire [13-1:0] node667;
	wire [13-1:0] node670;
	wire [13-1:0] node672;
	wire [13-1:0] node675;
	wire [13-1:0] node676;
	wire [13-1:0] node677;
	wire [13-1:0] node678;
	wire [13-1:0] node679;
	wire [13-1:0] node680;
	wire [13-1:0] node681;
	wire [13-1:0] node682;
	wire [13-1:0] node683;
	wire [13-1:0] node686;
	wire [13-1:0] node689;
	wire [13-1:0] node690;
	wire [13-1:0] node694;
	wire [13-1:0] node695;
	wire [13-1:0] node696;
	wire [13-1:0] node699;
	wire [13-1:0] node702;
	wire [13-1:0] node703;
	wire [13-1:0] node706;
	wire [13-1:0] node709;
	wire [13-1:0] node710;
	wire [13-1:0] node711;
	wire [13-1:0] node712;
	wire [13-1:0] node715;
	wire [13-1:0] node718;
	wire [13-1:0] node719;
	wire [13-1:0] node723;
	wire [13-1:0] node726;
	wire [13-1:0] node727;
	wire [13-1:0] node728;
	wire [13-1:0] node729;
	wire [13-1:0] node730;
	wire [13-1:0] node734;
	wire [13-1:0] node737;
	wire [13-1:0] node738;
	wire [13-1:0] node741;
	wire [13-1:0] node743;
	wire [13-1:0] node746;
	wire [13-1:0] node747;
	wire [13-1:0] node749;
	wire [13-1:0] node752;
	wire [13-1:0] node755;
	wire [13-1:0] node756;
	wire [13-1:0] node757;
	wire [13-1:0] node758;
	wire [13-1:0] node759;
	wire [13-1:0] node760;
	wire [13-1:0] node764;
	wire [13-1:0] node767;
	wire [13-1:0] node768;
	wire [13-1:0] node771;
	wire [13-1:0] node772;
	wire [13-1:0] node776;
	wire [13-1:0] node777;
	wire [13-1:0] node778;
	wire [13-1:0] node780;
	wire [13-1:0] node784;
	wire [13-1:0] node786;
	wire [13-1:0] node789;
	wire [13-1:0] node790;
	wire [13-1:0] node791;
	wire [13-1:0] node793;
	wire [13-1:0] node794;
	wire [13-1:0] node798;
	wire [13-1:0] node799;
	wire [13-1:0] node800;
	wire [13-1:0] node803;
	wire [13-1:0] node806;
	wire [13-1:0] node807;
	wire [13-1:0] node811;
	wire [13-1:0] node812;
	wire [13-1:0] node813;
	wire [13-1:0] node814;
	wire [13-1:0] node819;
	wire [13-1:0] node820;
	wire [13-1:0] node821;
	wire [13-1:0] node825;
	wire [13-1:0] node827;
	wire [13-1:0] node830;
	wire [13-1:0] node831;
	wire [13-1:0] node832;
	wire [13-1:0] node833;
	wire [13-1:0] node834;
	wire [13-1:0] node835;
	wire [13-1:0] node836;
	wire [13-1:0] node841;
	wire [13-1:0] node842;
	wire [13-1:0] node843;
	wire [13-1:0] node846;
	wire [13-1:0] node849;
	wire [13-1:0] node850;
	wire [13-1:0] node853;
	wire [13-1:0] node856;
	wire [13-1:0] node857;
	wire [13-1:0] node858;
	wire [13-1:0] node859;
	wire [13-1:0] node862;
	wire [13-1:0] node866;
	wire [13-1:0] node867;
	wire [13-1:0] node871;
	wire [13-1:0] node872;
	wire [13-1:0] node873;
	wire [13-1:0] node874;
	wire [13-1:0] node878;
	wire [13-1:0] node879;
	wire [13-1:0] node880;
	wire [13-1:0] node883;
	wire [13-1:0] node887;
	wire [13-1:0] node888;
	wire [13-1:0] node889;
	wire [13-1:0] node893;
	wire [13-1:0] node894;
	wire [13-1:0] node896;
	wire [13-1:0] node899;
	wire [13-1:0] node901;
	wire [13-1:0] node904;
	wire [13-1:0] node905;
	wire [13-1:0] node906;
	wire [13-1:0] node907;
	wire [13-1:0] node908;
	wire [13-1:0] node909;
	wire [13-1:0] node914;
	wire [13-1:0] node915;
	wire [13-1:0] node916;
	wire [13-1:0] node920;
	wire [13-1:0] node922;
	wire [13-1:0] node925;
	wire [13-1:0] node926;
	wire [13-1:0] node927;
	wire [13-1:0] node928;
	wire [13-1:0] node932;
	wire [13-1:0] node933;
	wire [13-1:0] node937;
	wire [13-1:0] node938;
	wire [13-1:0] node940;
	wire [13-1:0] node943;
	wire [13-1:0] node944;
	wire [13-1:0] node947;
	wire [13-1:0] node950;
	wire [13-1:0] node951;
	wire [13-1:0] node952;
	wire [13-1:0] node953;
	wire [13-1:0] node955;
	wire [13-1:0] node958;
	wire [13-1:0] node959;
	wire [13-1:0] node963;
	wire [13-1:0] node964;
	wire [13-1:0] node966;
	wire [13-1:0] node970;
	wire [13-1:0] node971;
	wire [13-1:0] node972;
	wire [13-1:0] node973;
	wire [13-1:0] node976;
	wire [13-1:0] node979;
	wire [13-1:0] node980;
	wire [13-1:0] node983;
	wire [13-1:0] node986;
	wire [13-1:0] node987;
	wire [13-1:0] node989;
	wire [13-1:0] node992;
	wire [13-1:0] node993;
	wire [13-1:0] node997;
	wire [13-1:0] node998;
	wire [13-1:0] node999;
	wire [13-1:0] node1000;
	wire [13-1:0] node1001;
	wire [13-1:0] node1002;
	wire [13-1:0] node1003;
	wire [13-1:0] node1007;
	wire [13-1:0] node1009;
	wire [13-1:0] node1012;
	wire [13-1:0] node1013;
	wire [13-1:0] node1014;
	wire [13-1:0] node1017;
	wire [13-1:0] node1018;
	wire [13-1:0] node1022;
	wire [13-1:0] node1023;
	wire [13-1:0] node1024;
	wire [13-1:0] node1028;
	wire [13-1:0] node1031;
	wire [13-1:0] node1032;
	wire [13-1:0] node1033;
	wire [13-1:0] node1034;
	wire [13-1:0] node1035;
	wire [13-1:0] node1039;
	wire [13-1:0] node1042;
	wire [13-1:0] node1044;
	wire [13-1:0] node1045;
	wire [13-1:0] node1049;
	wire [13-1:0] node1050;
	wire [13-1:0] node1051;
	wire [13-1:0] node1052;
	wire [13-1:0] node1056;
	wire [13-1:0] node1057;
	wire [13-1:0] node1061;
	wire [13-1:0] node1062;
	wire [13-1:0] node1063;
	wire [13-1:0] node1066;
	wire [13-1:0] node1070;
	wire [13-1:0] node1071;
	wire [13-1:0] node1072;
	wire [13-1:0] node1073;
	wire [13-1:0] node1075;
	wire [13-1:0] node1076;
	wire [13-1:0] node1080;
	wire [13-1:0] node1082;
	wire [13-1:0] node1083;
	wire [13-1:0] node1087;
	wire [13-1:0] node1088;
	wire [13-1:0] node1089;
	wire [13-1:0] node1092;
	wire [13-1:0] node1093;
	wire [13-1:0] node1097;
	wire [13-1:0] node1098;
	wire [13-1:0] node1100;
	wire [13-1:0] node1104;
	wire [13-1:0] node1105;
	wire [13-1:0] node1106;
	wire [13-1:0] node1108;
	wire [13-1:0] node1109;
	wire [13-1:0] node1113;
	wire [13-1:0] node1115;
	wire [13-1:0] node1117;
	wire [13-1:0] node1120;
	wire [13-1:0] node1121;
	wire [13-1:0] node1122;
	wire [13-1:0] node1123;
	wire [13-1:0] node1127;
	wire [13-1:0] node1130;
	wire [13-1:0] node1131;
	wire [13-1:0] node1132;
	wire [13-1:0] node1135;
	wire [13-1:0] node1139;
	wire [13-1:0] node1140;
	wire [13-1:0] node1141;
	wire [13-1:0] node1142;
	wire [13-1:0] node1143;
	wire [13-1:0] node1144;
	wire [13-1:0] node1146;
	wire [13-1:0] node1149;
	wire [13-1:0] node1152;
	wire [13-1:0] node1154;
	wire [13-1:0] node1157;
	wire [13-1:0] node1158;
	wire [13-1:0] node1159;
	wire [13-1:0] node1160;
	wire [13-1:0] node1163;
	wire [13-1:0] node1166;
	wire [13-1:0] node1167;
	wire [13-1:0] node1171;
	wire [13-1:0] node1172;
	wire [13-1:0] node1173;
	wire [13-1:0] node1177;
	wire [13-1:0] node1179;
	wire [13-1:0] node1182;
	wire [13-1:0] node1183;
	wire [13-1:0] node1184;
	wire [13-1:0] node1187;
	wire [13-1:0] node1189;
	wire [13-1:0] node1190;
	wire [13-1:0] node1194;
	wire [13-1:0] node1195;
	wire [13-1:0] node1196;
	wire [13-1:0] node1198;
	wire [13-1:0] node1201;
	wire [13-1:0] node1202;
	wire [13-1:0] node1205;
	wire [13-1:0] node1208;
	wire [13-1:0] node1209;
	wire [13-1:0] node1210;
	wire [13-1:0] node1213;
	wire [13-1:0] node1216;
	wire [13-1:0] node1217;
	wire [13-1:0] node1220;
	wire [13-1:0] node1223;
	wire [13-1:0] node1224;
	wire [13-1:0] node1225;
	wire [13-1:0] node1226;
	wire [13-1:0] node1228;
	wire [13-1:0] node1231;
	wire [13-1:0] node1232;
	wire [13-1:0] node1233;
	wire [13-1:0] node1236;
	wire [13-1:0] node1239;
	wire [13-1:0] node1241;
	wire [13-1:0] node1244;
	wire [13-1:0] node1245;
	wire [13-1:0] node1247;
	wire [13-1:0] node1248;
	wire [13-1:0] node1252;
	wire [13-1:0] node1253;
	wire [13-1:0] node1254;
	wire [13-1:0] node1257;
	wire [13-1:0] node1261;
	wire [13-1:0] node1262;
	wire [13-1:0] node1263;
	wire [13-1:0] node1265;
	wire [13-1:0] node1268;
	wire [13-1:0] node1270;
	wire [13-1:0] node1272;
	wire [13-1:0] node1275;
	wire [13-1:0] node1276;
	wire [13-1:0] node1277;
	wire [13-1:0] node1278;
	wire [13-1:0] node1281;
	wire [13-1:0] node1284;
	wire [13-1:0] node1286;
	wire [13-1:0] node1289;
	wire [13-1:0] node1290;
	wire [13-1:0] node1291;
	wire [13-1:0] node1294;
	wire [13-1:0] node1297;
	wire [13-1:0] node1298;
	wire [13-1:0] node1301;
	wire [13-1:0] node1304;
	wire [13-1:0] node1305;
	wire [13-1:0] node1306;
	wire [13-1:0] node1307;
	wire [13-1:0] node1308;
	wire [13-1:0] node1309;
	wire [13-1:0] node1310;
	wire [13-1:0] node1311;
	wire [13-1:0] node1312;
	wire [13-1:0] node1313;
	wire [13-1:0] node1316;
	wire [13-1:0] node1319;
	wire [13-1:0] node1321;
	wire [13-1:0] node1324;
	wire [13-1:0] node1325;
	wire [13-1:0] node1326;
	wire [13-1:0] node1329;
	wire [13-1:0] node1332;
	wire [13-1:0] node1335;
	wire [13-1:0] node1336;
	wire [13-1:0] node1337;
	wire [13-1:0] node1340;
	wire [13-1:0] node1341;
	wire [13-1:0] node1345;
	wire [13-1:0] node1346;
	wire [13-1:0] node1350;
	wire [13-1:0] node1351;
	wire [13-1:0] node1352;
	wire [13-1:0] node1353;
	wire [13-1:0] node1355;
	wire [13-1:0] node1358;
	wire [13-1:0] node1361;
	wire [13-1:0] node1363;
	wire [13-1:0] node1365;
	wire [13-1:0] node1368;
	wire [13-1:0] node1369;
	wire [13-1:0] node1370;
	wire [13-1:0] node1371;
	wire [13-1:0] node1376;
	wire [13-1:0] node1377;
	wire [13-1:0] node1378;
	wire [13-1:0] node1381;
	wire [13-1:0] node1385;
	wire [13-1:0] node1386;
	wire [13-1:0] node1387;
	wire [13-1:0] node1388;
	wire [13-1:0] node1390;
	wire [13-1:0] node1391;
	wire [13-1:0] node1394;
	wire [13-1:0] node1397;
	wire [13-1:0] node1399;
	wire [13-1:0] node1402;
	wire [13-1:0] node1403;
	wire [13-1:0] node1404;
	wire [13-1:0] node1407;
	wire [13-1:0] node1408;
	wire [13-1:0] node1412;
	wire [13-1:0] node1414;
	wire [13-1:0] node1417;
	wire [13-1:0] node1418;
	wire [13-1:0] node1419;
	wire [13-1:0] node1421;
	wire [13-1:0] node1424;
	wire [13-1:0] node1425;
	wire [13-1:0] node1427;
	wire [13-1:0] node1431;
	wire [13-1:0] node1432;
	wire [13-1:0] node1433;
	wire [13-1:0] node1436;
	wire [13-1:0] node1438;
	wire [13-1:0] node1441;
	wire [13-1:0] node1442;
	wire [13-1:0] node1443;
	wire [13-1:0] node1446;
	wire [13-1:0] node1449;
	wire [13-1:0] node1451;
	wire [13-1:0] node1454;
	wire [13-1:0] node1455;
	wire [13-1:0] node1456;
	wire [13-1:0] node1457;
	wire [13-1:0] node1458;
	wire [13-1:0] node1459;
	wire [13-1:0] node1462;
	wire [13-1:0] node1463;
	wire [13-1:0] node1467;
	wire [13-1:0] node1468;
	wire [13-1:0] node1470;
	wire [13-1:0] node1473;
	wire [13-1:0] node1475;
	wire [13-1:0] node1478;
	wire [13-1:0] node1479;
	wire [13-1:0] node1480;
	wire [13-1:0] node1483;
	wire [13-1:0] node1484;
	wire [13-1:0] node1488;
	wire [13-1:0] node1489;
	wire [13-1:0] node1490;
	wire [13-1:0] node1493;
	wire [13-1:0] node1496;
	wire [13-1:0] node1499;
	wire [13-1:0] node1500;
	wire [13-1:0] node1501;
	wire [13-1:0] node1503;
	wire [13-1:0] node1506;
	wire [13-1:0] node1507;
	wire [13-1:0] node1509;
	wire [13-1:0] node1512;
	wire [13-1:0] node1513;
	wire [13-1:0] node1517;
	wire [13-1:0] node1518;
	wire [13-1:0] node1520;
	wire [13-1:0] node1521;
	wire [13-1:0] node1525;
	wire [13-1:0] node1526;
	wire [13-1:0] node1528;
	wire [13-1:0] node1531;
	wire [13-1:0] node1532;
	wire [13-1:0] node1535;
	wire [13-1:0] node1538;
	wire [13-1:0] node1539;
	wire [13-1:0] node1540;
	wire [13-1:0] node1541;
	wire [13-1:0] node1544;
	wire [13-1:0] node1545;
	wire [13-1:0] node1548;
	wire [13-1:0] node1549;
	wire [13-1:0] node1553;
	wire [13-1:0] node1554;
	wire [13-1:0] node1555;
	wire [13-1:0] node1556;
	wire [13-1:0] node1561;
	wire [13-1:0] node1562;
	wire [13-1:0] node1564;
	wire [13-1:0] node1567;
	wire [13-1:0] node1570;
	wire [13-1:0] node1571;
	wire [13-1:0] node1572;
	wire [13-1:0] node1573;
	wire [13-1:0] node1576;
	wire [13-1:0] node1578;
	wire [13-1:0] node1581;
	wire [13-1:0] node1582;
	wire [13-1:0] node1584;
	wire [13-1:0] node1587;
	wire [13-1:0] node1590;
	wire [13-1:0] node1591;
	wire [13-1:0] node1592;
	wire [13-1:0] node1594;
	wire [13-1:0] node1597;
	wire [13-1:0] node1598;
	wire [13-1:0] node1602;
	wire [13-1:0] node1603;
	wire [13-1:0] node1604;
	wire [13-1:0] node1607;
	wire [13-1:0] node1610;
	wire [13-1:0] node1613;
	wire [13-1:0] node1614;
	wire [13-1:0] node1615;
	wire [13-1:0] node1616;
	wire [13-1:0] node1617;
	wire [13-1:0] node1618;
	wire [13-1:0] node1620;
	wire [13-1:0] node1623;
	wire [13-1:0] node1624;
	wire [13-1:0] node1625;
	wire [13-1:0] node1628;
	wire [13-1:0] node1632;
	wire [13-1:0] node1633;
	wire [13-1:0] node1634;
	wire [13-1:0] node1635;
	wire [13-1:0] node1639;
	wire [13-1:0] node1640;
	wire [13-1:0] node1644;
	wire [13-1:0] node1645;
	wire [13-1:0] node1646;
	wire [13-1:0] node1650;
	wire [13-1:0] node1651;
	wire [13-1:0] node1655;
	wire [13-1:0] node1656;
	wire [13-1:0] node1657;
	wire [13-1:0] node1658;
	wire [13-1:0] node1659;
	wire [13-1:0] node1662;
	wire [13-1:0] node1665;
	wire [13-1:0] node1666;
	wire [13-1:0] node1669;
	wire [13-1:0] node1672;
	wire [13-1:0] node1674;
	wire [13-1:0] node1677;
	wire [13-1:0] node1678;
	wire [13-1:0] node1679;
	wire [13-1:0] node1680;
	wire [13-1:0] node1683;
	wire [13-1:0] node1687;
	wire [13-1:0] node1689;
	wire [13-1:0] node1690;
	wire [13-1:0] node1693;
	wire [13-1:0] node1696;
	wire [13-1:0] node1697;
	wire [13-1:0] node1698;
	wire [13-1:0] node1699;
	wire [13-1:0] node1700;
	wire [13-1:0] node1701;
	wire [13-1:0] node1704;
	wire [13-1:0] node1707;
	wire [13-1:0] node1708;
	wire [13-1:0] node1711;
	wire [13-1:0] node1714;
	wire [13-1:0] node1715;
	wire [13-1:0] node1716;
	wire [13-1:0] node1720;
	wire [13-1:0] node1722;
	wire [13-1:0] node1725;
	wire [13-1:0] node1726;
	wire [13-1:0] node1727;
	wire [13-1:0] node1728;
	wire [13-1:0] node1731;
	wire [13-1:0] node1734;
	wire [13-1:0] node1736;
	wire [13-1:0] node1739;
	wire [13-1:0] node1740;
	wire [13-1:0] node1743;
	wire [13-1:0] node1745;
	wire [13-1:0] node1748;
	wire [13-1:0] node1749;
	wire [13-1:0] node1750;
	wire [13-1:0] node1751;
	wire [13-1:0] node1753;
	wire [13-1:0] node1756;
	wire [13-1:0] node1757;
	wire [13-1:0] node1760;
	wire [13-1:0] node1763;
	wire [13-1:0] node1764;
	wire [13-1:0] node1766;
	wire [13-1:0] node1769;
	wire [13-1:0] node1770;
	wire [13-1:0] node1773;
	wire [13-1:0] node1776;
	wire [13-1:0] node1777;
	wire [13-1:0] node1778;
	wire [13-1:0] node1779;
	wire [13-1:0] node1782;
	wire [13-1:0] node1785;
	wire [13-1:0] node1786;
	wire [13-1:0] node1789;
	wire [13-1:0] node1792;
	wire [13-1:0] node1793;
	wire [13-1:0] node1795;
	wire [13-1:0] node1799;
	wire [13-1:0] node1800;
	wire [13-1:0] node1801;
	wire [13-1:0] node1802;
	wire [13-1:0] node1804;
	wire [13-1:0] node1805;
	wire [13-1:0] node1806;
	wire [13-1:0] node1810;
	wire [13-1:0] node1813;
	wire [13-1:0] node1814;
	wire [13-1:0] node1815;
	wire [13-1:0] node1816;
	wire [13-1:0] node1820;
	wire [13-1:0] node1821;
	wire [13-1:0] node1825;
	wire [13-1:0] node1826;
	wire [13-1:0] node1827;
	wire [13-1:0] node1830;
	wire [13-1:0] node1834;
	wire [13-1:0] node1835;
	wire [13-1:0] node1836;
	wire [13-1:0] node1837;
	wire [13-1:0] node1838;
	wire [13-1:0] node1841;
	wire [13-1:0] node1844;
	wire [13-1:0] node1845;
	wire [13-1:0] node1848;
	wire [13-1:0] node1851;
	wire [13-1:0] node1852;
	wire [13-1:0] node1853;
	wire [13-1:0] node1857;
	wire [13-1:0] node1858;
	wire [13-1:0] node1862;
	wire [13-1:0] node1863;
	wire [13-1:0] node1864;
	wire [13-1:0] node1866;
	wire [13-1:0] node1869;
	wire [13-1:0] node1870;
	wire [13-1:0] node1873;
	wire [13-1:0] node1876;
	wire [13-1:0] node1877;
	wire [13-1:0] node1880;
	wire [13-1:0] node1881;
	wire [13-1:0] node1885;
	wire [13-1:0] node1886;
	wire [13-1:0] node1887;
	wire [13-1:0] node1888;
	wire [13-1:0] node1889;
	wire [13-1:0] node1891;
	wire [13-1:0] node1894;
	wire [13-1:0] node1895;
	wire [13-1:0] node1898;
	wire [13-1:0] node1901;
	wire [13-1:0] node1902;
	wire [13-1:0] node1903;
	wire [13-1:0] node1906;
	wire [13-1:0] node1909;
	wire [13-1:0] node1912;
	wire [13-1:0] node1913;
	wire [13-1:0] node1914;
	wire [13-1:0] node1915;
	wire [13-1:0] node1918;
	wire [13-1:0] node1922;
	wire [13-1:0] node1924;
	wire [13-1:0] node1925;
	wire [13-1:0] node1928;
	wire [13-1:0] node1931;
	wire [13-1:0] node1932;
	wire [13-1:0] node1933;
	wire [13-1:0] node1934;
	wire [13-1:0] node1937;
	wire [13-1:0] node1938;
	wire [13-1:0] node1941;
	wire [13-1:0] node1944;
	wire [13-1:0] node1945;
	wire [13-1:0] node1947;
	wire [13-1:0] node1951;
	wire [13-1:0] node1952;
	wire [13-1:0] node1953;
	wire [13-1:0] node1954;
	wire [13-1:0] node1959;
	wire [13-1:0] node1960;
	wire [13-1:0] node1962;
	wire [13-1:0] node1965;
	wire [13-1:0] node1967;
	wire [13-1:0] node1970;
	wire [13-1:0] node1971;
	wire [13-1:0] node1972;
	wire [13-1:0] node1973;
	wire [13-1:0] node1974;
	wire [13-1:0] node1975;
	wire [13-1:0] node1976;
	wire [13-1:0] node1978;
	wire [13-1:0] node1979;
	wire [13-1:0] node1983;
	wire [13-1:0] node1984;
	wire [13-1:0] node1985;
	wire [13-1:0] node1988;
	wire [13-1:0] node1992;
	wire [13-1:0] node1993;
	wire [13-1:0] node1994;
	wire [13-1:0] node1997;
	wire [13-1:0] node1999;
	wire [13-1:0] node2002;
	wire [13-1:0] node2003;
	wire [13-1:0] node2005;
	wire [13-1:0] node2008;
	wire [13-1:0] node2011;
	wire [13-1:0] node2012;
	wire [13-1:0] node2013;
	wire [13-1:0] node2014;
	wire [13-1:0] node2015;
	wire [13-1:0] node2018;
	wire [13-1:0] node2021;
	wire [13-1:0] node2022;
	wire [13-1:0] node2025;
	wire [13-1:0] node2028;
	wire [13-1:0] node2029;
	wire [13-1:0] node2030;
	wire [13-1:0] node2033;
	wire [13-1:0] node2037;
	wire [13-1:0] node2038;
	wire [13-1:0] node2039;
	wire [13-1:0] node2040;
	wire [13-1:0] node2044;
	wire [13-1:0] node2045;
	wire [13-1:0] node2049;
	wire [13-1:0] node2051;
	wire [13-1:0] node2053;
	wire [13-1:0] node2056;
	wire [13-1:0] node2057;
	wire [13-1:0] node2058;
	wire [13-1:0] node2059;
	wire [13-1:0] node2060;
	wire [13-1:0] node2062;
	wire [13-1:0] node2065;
	wire [13-1:0] node2066;
	wire [13-1:0] node2070;
	wire [13-1:0] node2072;
	wire [13-1:0] node2075;
	wire [13-1:0] node2076;
	wire [13-1:0] node2077;
	wire [13-1:0] node2078;
	wire [13-1:0] node2081;
	wire [13-1:0] node2084;
	wire [13-1:0] node2086;
	wire [13-1:0] node2089;
	wire [13-1:0] node2090;
	wire [13-1:0] node2091;
	wire [13-1:0] node2095;
	wire [13-1:0] node2097;
	wire [13-1:0] node2100;
	wire [13-1:0] node2101;
	wire [13-1:0] node2102;
	wire [13-1:0] node2103;
	wire [13-1:0] node2105;
	wire [13-1:0] node2108;
	wire [13-1:0] node2110;
	wire [13-1:0] node2113;
	wire [13-1:0] node2114;
	wire [13-1:0] node2115;
	wire [13-1:0] node2118;
	wire [13-1:0] node2121;
	wire [13-1:0] node2122;
	wire [13-1:0] node2125;
	wire [13-1:0] node2128;
	wire [13-1:0] node2129;
	wire [13-1:0] node2130;
	wire [13-1:0] node2132;
	wire [13-1:0] node2135;
	wire [13-1:0] node2138;
	wire [13-1:0] node2139;
	wire [13-1:0] node2142;
	wire [13-1:0] node2145;
	wire [13-1:0] node2146;
	wire [13-1:0] node2147;
	wire [13-1:0] node2148;
	wire [13-1:0] node2149;
	wire [13-1:0] node2150;
	wire [13-1:0] node2151;
	wire [13-1:0] node2154;
	wire [13-1:0] node2158;
	wire [13-1:0] node2160;
	wire [13-1:0] node2161;
	wire [13-1:0] node2165;
	wire [13-1:0] node2166;
	wire [13-1:0] node2167;
	wire [13-1:0] node2169;
	wire [13-1:0] node2172;
	wire [13-1:0] node2175;
	wire [13-1:0] node2177;
	wire [13-1:0] node2178;
	wire [13-1:0] node2182;
	wire [13-1:0] node2183;
	wire [13-1:0] node2184;
	wire [13-1:0] node2185;
	wire [13-1:0] node2187;
	wire [13-1:0] node2190;
	wire [13-1:0] node2191;
	wire [13-1:0] node2195;
	wire [13-1:0] node2197;
	wire [13-1:0] node2200;
	wire [13-1:0] node2201;
	wire [13-1:0] node2202;
	wire [13-1:0] node2203;
	wire [13-1:0] node2206;
	wire [13-1:0] node2209;
	wire [13-1:0] node2210;
	wire [13-1:0] node2213;
	wire [13-1:0] node2216;
	wire [13-1:0] node2218;
	wire [13-1:0] node2220;
	wire [13-1:0] node2223;
	wire [13-1:0] node2224;
	wire [13-1:0] node2225;
	wire [13-1:0] node2226;
	wire [13-1:0] node2227;
	wire [13-1:0] node2229;
	wire [13-1:0] node2232;
	wire [13-1:0] node2233;
	wire [13-1:0] node2236;
	wire [13-1:0] node2239;
	wire [13-1:0] node2240;
	wire [13-1:0] node2242;
	wire [13-1:0] node2245;
	wire [13-1:0] node2247;
	wire [13-1:0] node2250;
	wire [13-1:0] node2251;
	wire [13-1:0] node2252;
	wire [13-1:0] node2255;
	wire [13-1:0] node2256;
	wire [13-1:0] node2259;
	wire [13-1:0] node2262;
	wire [13-1:0] node2263;
	wire [13-1:0] node2266;
	wire [13-1:0] node2267;
	wire [13-1:0] node2271;
	wire [13-1:0] node2272;
	wire [13-1:0] node2273;
	wire [13-1:0] node2274;
	wire [13-1:0] node2275;
	wire [13-1:0] node2279;
	wire [13-1:0] node2282;
	wire [13-1:0] node2283;
	wire [13-1:0] node2286;
	wire [13-1:0] node2287;
	wire [13-1:0] node2290;
	wire [13-1:0] node2293;
	wire [13-1:0] node2294;
	wire [13-1:0] node2296;
	wire [13-1:0] node2297;
	wire [13-1:0] node2301;
	wire [13-1:0] node2303;
	wire [13-1:0] node2304;
	wire [13-1:0] node2308;
	wire [13-1:0] node2309;
	wire [13-1:0] node2310;
	wire [13-1:0] node2311;
	wire [13-1:0] node2312;
	wire [13-1:0] node2313;
	wire [13-1:0] node2314;
	wire [13-1:0] node2315;
	wire [13-1:0] node2318;
	wire [13-1:0] node2321;
	wire [13-1:0] node2323;
	wire [13-1:0] node2326;
	wire [13-1:0] node2327;
	wire [13-1:0] node2328;
	wire [13-1:0] node2332;
	wire [13-1:0] node2335;
	wire [13-1:0] node2336;
	wire [13-1:0] node2337;
	wire [13-1:0] node2338;
	wire [13-1:0] node2342;
	wire [13-1:0] node2343;
	wire [13-1:0] node2347;
	wire [13-1:0] node2349;
	wire [13-1:0] node2350;
	wire [13-1:0] node2353;
	wire [13-1:0] node2356;
	wire [13-1:0] node2357;
	wire [13-1:0] node2358;
	wire [13-1:0] node2359;
	wire [13-1:0] node2363;
	wire [13-1:0] node2365;
	wire [13-1:0] node2366;
	wire [13-1:0] node2370;
	wire [13-1:0] node2371;
	wire [13-1:0] node2372;
	wire [13-1:0] node2373;
	wire [13-1:0] node2377;
	wire [13-1:0] node2378;
	wire [13-1:0] node2382;
	wire [13-1:0] node2384;
	wire [13-1:0] node2387;
	wire [13-1:0] node2388;
	wire [13-1:0] node2389;
	wire [13-1:0] node2390;
	wire [13-1:0] node2391;
	wire [13-1:0] node2392;
	wire [13-1:0] node2395;
	wire [13-1:0] node2398;
	wire [13-1:0] node2400;
	wire [13-1:0] node2403;
	wire [13-1:0] node2404;
	wire [13-1:0] node2405;
	wire [13-1:0] node2408;
	wire [13-1:0] node2411;
	wire [13-1:0] node2413;
	wire [13-1:0] node2416;
	wire [13-1:0] node2417;
	wire [13-1:0] node2418;
	wire [13-1:0] node2421;
	wire [13-1:0] node2423;
	wire [13-1:0] node2426;
	wire [13-1:0] node2427;
	wire [13-1:0] node2428;
	wire [13-1:0] node2431;
	wire [13-1:0] node2434;
	wire [13-1:0] node2436;
	wire [13-1:0] node2439;
	wire [13-1:0] node2440;
	wire [13-1:0] node2441;
	wire [13-1:0] node2442;
	wire [13-1:0] node2444;
	wire [13-1:0] node2447;
	wire [13-1:0] node2449;
	wire [13-1:0] node2452;
	wire [13-1:0] node2453;
	wire [13-1:0] node2454;
	wire [13-1:0] node2457;
	wire [13-1:0] node2461;
	wire [13-1:0] node2462;
	wire [13-1:0] node2463;
	wire [13-1:0] node2464;
	wire [13-1:0] node2468;
	wire [13-1:0] node2469;
	wire [13-1:0] node2473;
	wire [13-1:0] node2474;
	wire [13-1:0] node2477;
	wire [13-1:0] node2479;
	wire [13-1:0] node2482;
	wire [13-1:0] node2483;
	wire [13-1:0] node2484;
	wire [13-1:0] node2485;
	wire [13-1:0] node2486;
	wire [13-1:0] node2487;
	wire [13-1:0] node2488;
	wire [13-1:0] node2491;
	wire [13-1:0] node2495;
	wire [13-1:0] node2497;
	wire [13-1:0] node2500;
	wire [13-1:0] node2501;
	wire [13-1:0] node2502;
	wire [13-1:0] node2505;
	wire [13-1:0] node2506;
	wire [13-1:0] node2509;
	wire [13-1:0] node2512;
	wire [13-1:0] node2514;
	wire [13-1:0] node2515;
	wire [13-1:0] node2518;
	wire [13-1:0] node2521;
	wire [13-1:0] node2522;
	wire [13-1:0] node2523;
	wire [13-1:0] node2524;
	wire [13-1:0] node2525;
	wire [13-1:0] node2528;
	wire [13-1:0] node2531;
	wire [13-1:0] node2532;
	wire [13-1:0] node2535;
	wire [13-1:0] node2538;
	wire [13-1:0] node2539;
	wire [13-1:0] node2541;
	wire [13-1:0] node2544;
	wire [13-1:0] node2545;
	wire [13-1:0] node2548;
	wire [13-1:0] node2551;
	wire [13-1:0] node2552;
	wire [13-1:0] node2553;
	wire [13-1:0] node2554;
	wire [13-1:0] node2558;
	wire [13-1:0] node2559;
	wire [13-1:0] node2563;
	wire [13-1:0] node2564;
	wire [13-1:0] node2565;
	wire [13-1:0] node2568;
	wire [13-1:0] node2571;
	wire [13-1:0] node2572;
	wire [13-1:0] node2575;
	wire [13-1:0] node2578;
	wire [13-1:0] node2579;
	wire [13-1:0] node2580;
	wire [13-1:0] node2581;
	wire [13-1:0] node2582;
	wire [13-1:0] node2583;
	wire [13-1:0] node2587;
	wire [13-1:0] node2589;
	wire [13-1:0] node2592;
	wire [13-1:0] node2593;
	wire [13-1:0] node2594;
	wire [13-1:0] node2597;
	wire [13-1:0] node2600;
	wire [13-1:0] node2601;
	wire [13-1:0] node2604;
	wire [13-1:0] node2607;
	wire [13-1:0] node2608;
	wire [13-1:0] node2609;
	wire [13-1:0] node2610;
	wire [13-1:0] node2614;
	wire [13-1:0] node2615;
	wire [13-1:0] node2619;
	wire [13-1:0] node2620;
	wire [13-1:0] node2623;
	wire [13-1:0] node2624;
	wire [13-1:0] node2627;
	wire [13-1:0] node2630;
	wire [13-1:0] node2631;
	wire [13-1:0] node2632;
	wire [13-1:0] node2634;
	wire [13-1:0] node2635;
	wire [13-1:0] node2639;
	wire [13-1:0] node2640;
	wire [13-1:0] node2641;
	wire [13-1:0] node2644;
	wire [13-1:0] node2647;
	wire [13-1:0] node2649;
	wire [13-1:0] node2652;
	wire [13-1:0] node2653;
	wire [13-1:0] node2654;
	wire [13-1:0] node2656;
	wire [13-1:0] node2660;
	wire [13-1:0] node2661;
	wire [13-1:0] node2662;
	wire [13-1:0] node2665;
	wire [13-1:0] node2668;
	wire [13-1:0] node2669;

	assign outp = (inp[4]) ? node1304 : node1;
		assign node1 = (inp[10]) ? node675 : node2;
			assign node2 = (inp[2]) ? node352 : node3;
				assign node3 = (inp[1]) ? node173 : node4;
					assign node4 = (inp[11]) ? node100 : node5;
						assign node5 = (inp[9]) ? node57 : node6;
							assign node6 = (inp[3]) ? node34 : node7;
								assign node7 = (inp[12]) ? node21 : node8;
									assign node8 = (inp[6]) ? node14 : node9;
										assign node9 = (inp[0]) ? 13'b0011111111111 : node10;
											assign node10 = (inp[8]) ? 13'b0011111111111 : 13'b0111111111111;
										assign node14 = (inp[7]) ? node18 : node15;
											assign node15 = (inp[0]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node18 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node21 = (inp[5]) ? node29 : node22;
										assign node22 = (inp[6]) ? node26 : node23;
											assign node23 = (inp[8]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node26 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node29 = (inp[0]) ? 13'b0000111111111 : node30;
											assign node30 = (inp[6]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node34 = (inp[7]) ? node46 : node35;
									assign node35 = (inp[6]) ? node41 : node36;
										assign node36 = (inp[12]) ? 13'b0001111111111 : node37;
											assign node37 = (inp[0]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node41 = (inp[8]) ? node43 : 13'b0001111111111;
											assign node43 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node46 = (inp[5]) ? node54 : node47;
										assign node47 = (inp[6]) ? node51 : node48;
											assign node48 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node51 = (inp[8]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node54 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node57 = (inp[8]) ? node83 : node58;
								assign node58 = (inp[12]) ? node72 : node59;
									assign node59 = (inp[0]) ? node65 : node60;
										assign node60 = (inp[5]) ? 13'b0001111111111 : node61;
											assign node61 = (inp[6]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node65 = (inp[6]) ? node69 : node66;
											assign node66 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node69 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node72 = (inp[3]) ? node76 : node73;
										assign node73 = (inp[5]) ? 13'b0000111111111 : 13'b0000011111111;
										assign node76 = (inp[0]) ? node80 : node77;
											assign node77 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node80 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node83 = (inp[5]) ? node91 : node84;
									assign node84 = (inp[6]) ? 13'b0000011111111 : node85;
										assign node85 = (inp[0]) ? node87 : 13'b0000111111111;
											assign node87 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node91 = (inp[3]) ? node97 : node92;
										assign node92 = (inp[7]) ? 13'b0000011111111 : node93;
											assign node93 = (inp[0]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node97 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
						assign node100 = (inp[12]) ? node146 : node101;
							assign node101 = (inp[5]) ? node125 : node102;
								assign node102 = (inp[3]) ? node114 : node103;
									assign node103 = (inp[7]) ? node109 : node104;
										assign node104 = (inp[0]) ? node106 : 13'b0001111111111;
											assign node106 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node109 = (inp[0]) ? 13'b0000111111111 : node110;
											assign node110 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node114 = (inp[8]) ? node122 : node115;
										assign node115 = (inp[9]) ? node119 : node116;
											assign node116 = (inp[6]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node119 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node122 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
								assign node125 = (inp[9]) ? node131 : node126;
									assign node126 = (inp[6]) ? node128 : 13'b0000111111111;
										assign node128 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node131 = (inp[0]) ? node139 : node132;
										assign node132 = (inp[8]) ? node136 : node133;
											assign node133 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node136 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node139 = (inp[8]) ? node143 : node140;
											assign node140 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node143 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node146 = (inp[0]) ? node160 : node147;
								assign node147 = (inp[3]) ? node155 : node148;
									assign node148 = (inp[8]) ? 13'b0000011111111 : node149;
										assign node149 = (inp[9]) ? node151 : 13'b0000111111111;
											assign node151 = (inp[6]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node155 = (inp[8]) ? node157 : 13'b0000011111111;
										assign node157 = (inp[9]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node160 = (inp[6]) ? node168 : node161;
									assign node161 = (inp[9]) ? 13'b0000001111111 : node162;
										assign node162 = (inp[7]) ? node164 : 13'b0000011111111;
											assign node164 = (inp[8]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node168 = (inp[3]) ? node170 : 13'b0000001111111;
										assign node170 = (inp[7]) ? 13'b0000000111111 : 13'b0000000011111;
					assign node173 = (inp[8]) ? node269 : node174;
						assign node174 = (inp[6]) ? node224 : node175;
							assign node175 = (inp[12]) ? node205 : node176;
								assign node176 = (inp[5]) ? node192 : node177;
									assign node177 = (inp[3]) ? node185 : node178;
										assign node178 = (inp[0]) ? node182 : node179;
											assign node179 = (inp[9]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node182 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node185 = (inp[7]) ? node189 : node186;
											assign node186 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node189 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node192 = (inp[11]) ? node198 : node193;
										assign node193 = (inp[7]) ? 13'b0000111111111 : node194;
											assign node194 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node198 = (inp[0]) ? node202 : node199;
											assign node199 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node202 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node205 = (inp[7]) ? node211 : node206;
									assign node206 = (inp[11]) ? node208 : 13'b0000111111111;
										assign node208 = (inp[9]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node211 = (inp[0]) ? node219 : node212;
										assign node212 = (inp[9]) ? node216 : node213;
											assign node213 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node216 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node219 = (inp[5]) ? 13'b0000001111111 : node220;
											assign node220 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node224 = (inp[9]) ? node248 : node225;
								assign node225 = (inp[7]) ? node237 : node226;
									assign node226 = (inp[3]) ? node232 : node227;
										assign node227 = (inp[5]) ? 13'b0000111111111 : node228;
											assign node228 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node232 = (inp[12]) ? 13'b0000011111111 : node233;
											assign node233 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node237 = (inp[3]) ? node243 : node238;
										assign node238 = (inp[0]) ? 13'b0000011111111 : node239;
											assign node239 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node243 = (inp[0]) ? node245 : 13'b0000001111111;
											assign node245 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node248 = (inp[12]) ? node258 : node249;
									assign node249 = (inp[3]) ? node251 : 13'b0000011111111;
										assign node251 = (inp[7]) ? node255 : node252;
											assign node252 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node255 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node258 = (inp[11]) ? node264 : node259;
										assign node259 = (inp[0]) ? 13'b0000000111111 : node260;
											assign node260 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node264 = (inp[5]) ? node266 : 13'b0000000111111;
											assign node266 = (inp[0]) ? 13'b0000000001111 : 13'b0000000111111;
						assign node269 = (inp[7]) ? node309 : node270;
							assign node270 = (inp[9]) ? node288 : node271;
								assign node271 = (inp[11]) ? node281 : node272;
									assign node272 = (inp[3]) ? node276 : node273;
										assign node273 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node276 = (inp[12]) ? node278 : 13'b0000111111111;
											assign node278 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node281 = (inp[0]) ? 13'b0000001111111 : node282;
										assign node282 = (inp[6]) ? node284 : 13'b0000111111111;
											assign node284 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node288 = (inp[12]) ? node298 : node289;
									assign node289 = (inp[6]) ? node291 : 13'b0000011111111;
										assign node291 = (inp[5]) ? node295 : node292;
											assign node292 = (inp[11]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node295 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node298 = (inp[0]) ? node304 : node299;
										assign node299 = (inp[11]) ? 13'b0000001111111 : node300;
											assign node300 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node304 = (inp[11]) ? node306 : 13'b0000000111111;
											assign node306 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node309 = (inp[11]) ? node335 : node310;
								assign node310 = (inp[3]) ? node322 : node311;
									assign node311 = (inp[12]) ? node315 : node312;
										assign node312 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node315 = (inp[6]) ? node319 : node316;
											assign node316 = (inp[9]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node319 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node322 = (inp[5]) ? node328 : node323;
										assign node323 = (inp[12]) ? 13'b0000001111111 : node324;
											assign node324 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node328 = (inp[6]) ? node332 : node329;
											assign node329 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node332 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node335 = (inp[0]) ? node347 : node336;
									assign node336 = (inp[12]) ? node342 : node337;
										assign node337 = (inp[3]) ? 13'b0000000111111 : node338;
											assign node338 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node342 = (inp[9]) ? node344 : 13'b0000000111111;
											assign node344 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node347 = (inp[6]) ? 13'b0000000001111 : node348;
										assign node348 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
				assign node352 = (inp[3]) ? node532 : node353;
					assign node353 = (inp[5]) ? node437 : node354;
						assign node354 = (inp[12]) ? node400 : node355;
							assign node355 = (inp[9]) ? node383 : node356;
								assign node356 = (inp[7]) ? node370 : node357;
									assign node357 = (inp[1]) ? node363 : node358;
										assign node358 = (inp[0]) ? 13'b0001111111111 : node359;
											assign node359 = (inp[8]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node363 = (inp[6]) ? node367 : node364;
											assign node364 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node367 = (inp[0]) ? 13'b0000111111111 : 13'b0000011111111;
									assign node370 = (inp[0]) ? node378 : node371;
										assign node371 = (inp[8]) ? node375 : node372;
											assign node372 = (inp[1]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node375 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node378 = (inp[1]) ? 13'b0000001111111 : node379;
											assign node379 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node383 = (inp[8]) ? node391 : node384;
									assign node384 = (inp[11]) ? 13'b0000011111111 : node385;
										assign node385 = (inp[7]) ? 13'b0000111111111 : node386;
											assign node386 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node391 = (inp[0]) ? node395 : node392;
										assign node392 = (inp[6]) ? 13'b0000011111111 : 13'b0001111111111;
										assign node395 = (inp[7]) ? 13'b0000000111111 : node396;
											assign node396 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node400 = (inp[6]) ? node416 : node401;
								assign node401 = (inp[11]) ? node409 : node402;
									assign node402 = (inp[7]) ? node406 : node403;
										assign node403 = (inp[1]) ? 13'b0001111111111 : 13'b0000111111111;
										assign node406 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node409 = (inp[1]) ? 13'b0000001111111 : node410;
										assign node410 = (inp[0]) ? node412 : 13'b0000111111111;
											assign node412 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node416 = (inp[7]) ? node426 : node417;
									assign node417 = (inp[1]) ? node419 : 13'b0000011111111;
										assign node419 = (inp[0]) ? node423 : node420;
											assign node420 = (inp[8]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node423 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node426 = (inp[11]) ? node432 : node427;
										assign node427 = (inp[9]) ? node429 : 13'b0000011111111;
											assign node429 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node432 = (inp[1]) ? node434 : 13'b0000000111111;
											assign node434 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node437 = (inp[7]) ? node479 : node438;
							assign node438 = (inp[0]) ? node458 : node439;
								assign node439 = (inp[8]) ? node451 : node440;
									assign node440 = (inp[12]) ? node444 : node441;
										assign node441 = (inp[6]) ? 13'b0001111111111 : 13'b0000111111111;
										assign node444 = (inp[11]) ? node448 : node445;
											assign node445 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node448 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node451 = (inp[9]) ? 13'b0000001111111 : node452;
										assign node452 = (inp[1]) ? node454 : 13'b0000011111111;
											assign node454 = (inp[11]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node458 = (inp[8]) ? node472 : node459;
									assign node459 = (inp[11]) ? node465 : node460;
										assign node460 = (inp[1]) ? node462 : 13'b0000011111111;
											assign node462 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node465 = (inp[1]) ? node469 : node466;
											assign node466 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node469 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node472 = (inp[1]) ? node474 : 13'b0000001111111;
										assign node474 = (inp[9]) ? 13'b0000000011111 : node475;
											assign node475 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node479 = (inp[11]) ? node509 : node480;
								assign node480 = (inp[1]) ? node496 : node481;
									assign node481 = (inp[8]) ? node489 : node482;
										assign node482 = (inp[6]) ? node486 : node483;
											assign node483 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node486 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node489 = (inp[12]) ? node493 : node490;
											assign node490 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node493 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node496 = (inp[9]) ? node504 : node497;
										assign node497 = (inp[12]) ? node501 : node498;
											assign node498 = (inp[0]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node501 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node504 = (inp[6]) ? 13'b0000000011111 : node505;
											assign node505 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node509 = (inp[1]) ? node521 : node510;
									assign node510 = (inp[6]) ? node518 : node511;
										assign node511 = (inp[8]) ? node515 : node512;
											assign node512 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node515 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node518 = (inp[9]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node521 = (inp[12]) ? node525 : node522;
										assign node522 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node525 = (inp[0]) ? node529 : node526;
											assign node526 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node529 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
					assign node532 = (inp[9]) ? node610 : node533;
						assign node533 = (inp[5]) ? node567 : node534;
							assign node534 = (inp[8]) ? node550 : node535;
								assign node535 = (inp[6]) ? node543 : node536;
									assign node536 = (inp[0]) ? 13'b0000011111111 : node537;
										assign node537 = (inp[7]) ? 13'b0000111111111 : node538;
											assign node538 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node543 = (inp[7]) ? 13'b0000001111111 : node544;
										assign node544 = (inp[0]) ? 13'b0000001111111 : node545;
											assign node545 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node550 = (inp[0]) ? node560 : node551;
									assign node551 = (inp[12]) ? node557 : node552;
										assign node552 = (inp[6]) ? node554 : 13'b0000011111111;
											assign node554 = (inp[7]) ? 13'b0000011111111 : 13'b0000001111111;
										assign node557 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node560 = (inp[1]) ? node562 : 13'b0000001111111;
										assign node562 = (inp[11]) ? 13'b0000000111111 : node563;
											assign node563 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node567 = (inp[11]) ? node589 : node568;
								assign node568 = (inp[6]) ? node582 : node569;
									assign node569 = (inp[7]) ? node575 : node570;
										assign node570 = (inp[1]) ? node572 : 13'b0000111111111;
											assign node572 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node575 = (inp[8]) ? node579 : node576;
											assign node576 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node579 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node582 = (inp[0]) ? 13'b0000000111111 : node583;
										assign node583 = (inp[1]) ? 13'b0000001111111 : node584;
											assign node584 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node589 = (inp[1]) ? node601 : node590;
									assign node590 = (inp[12]) ? node596 : node591;
										assign node591 = (inp[8]) ? 13'b0000001111111 : node592;
											assign node592 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node596 = (inp[0]) ? 13'b0000000111111 : node597;
											assign node597 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node601 = (inp[12]) ? node607 : node602;
										assign node602 = (inp[7]) ? node604 : 13'b0000011111111;
											assign node604 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node607 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node610 = (inp[11]) ? node646 : node611;
							assign node611 = (inp[6]) ? node627 : node612;
								assign node612 = (inp[7]) ? node620 : node613;
									assign node613 = (inp[0]) ? 13'b0000000111111 : node614;
										assign node614 = (inp[12]) ? node616 : 13'b0000011111111;
											assign node616 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node620 = (inp[5]) ? node622 : 13'b0000001111111;
										assign node622 = (inp[8]) ? 13'b0000000111111 : node623;
											assign node623 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node627 = (inp[1]) ? node639 : node628;
									assign node628 = (inp[7]) ? node634 : node629;
										assign node629 = (inp[12]) ? node631 : 13'b0000001111111;
											assign node631 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node634 = (inp[5]) ? 13'b0000000111111 : node635;
											assign node635 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node639 = (inp[12]) ? 13'b0000000011111 : node640;
										assign node640 = (inp[8]) ? 13'b0000000001111 : node641;
											assign node641 = (inp[0]) ? 13'b0000000111111 : 13'b0000000111111;
							assign node646 = (inp[6]) ? node662 : node647;
								assign node647 = (inp[12]) ? node655 : node648;
									assign node648 = (inp[8]) ? node650 : 13'b0000000111111;
										assign node650 = (inp[1]) ? 13'b0000000111111 : node651;
											assign node651 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node655 = (inp[0]) ? node657 : 13'b0000000111111;
										assign node657 = (inp[7]) ? 13'b0000000001111 : node658;
											assign node658 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node662 = (inp[0]) ? node670 : node663;
									assign node663 = (inp[7]) ? node665 : 13'b0000000111111;
										assign node665 = (inp[8]) ? node667 : 13'b0000000011111;
											assign node667 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node670 = (inp[1]) ? node672 : 13'b0000000001111;
										assign node672 = (inp[5]) ? 13'b0000000000011 : 13'b0000000001111;
			assign node675 = (inp[3]) ? node997 : node676;
				assign node676 = (inp[1]) ? node830 : node677;
					assign node677 = (inp[8]) ? node755 : node678;
						assign node678 = (inp[9]) ? node726 : node679;
							assign node679 = (inp[11]) ? node709 : node680;
								assign node680 = (inp[0]) ? node694 : node681;
									assign node681 = (inp[6]) ? node689 : node682;
										assign node682 = (inp[7]) ? node686 : node683;
											assign node683 = (inp[2]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node686 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node689 = (inp[5]) ? 13'b0000111111111 : node690;
											assign node690 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node694 = (inp[7]) ? node702 : node695;
										assign node695 = (inp[5]) ? node699 : node696;
											assign node696 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node699 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node702 = (inp[12]) ? node706 : node703;
											assign node703 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node706 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node709 = (inp[12]) ? node723 : node710;
									assign node710 = (inp[5]) ? node718 : node711;
										assign node711 = (inp[7]) ? node715 : node712;
											assign node712 = (inp[0]) ? 13'b0000111111111 : 13'b0011111111111;
											assign node715 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node718 = (inp[7]) ? 13'b0000011111111 : node719;
											assign node719 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node723 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node726 = (inp[5]) ? node746 : node727;
								assign node727 = (inp[12]) ? node737 : node728;
									assign node728 = (inp[2]) ? node734 : node729;
										assign node729 = (inp[6]) ? 13'b0000111111111 : node730;
											assign node730 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node734 = (inp[7]) ? 13'b0000111111111 : 13'b0000011111111;
									assign node737 = (inp[0]) ? node741 : node738;
										assign node738 = (inp[6]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node741 = (inp[2]) ? node743 : 13'b0000001111111;
											assign node743 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node746 = (inp[2]) ? node752 : node747;
									assign node747 = (inp[12]) ? node749 : 13'b0000011111111;
										assign node749 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node752 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node755 = (inp[0]) ? node789 : node756;
							assign node756 = (inp[11]) ? node776 : node757;
								assign node757 = (inp[9]) ? node767 : node758;
									assign node758 = (inp[7]) ? node764 : node759;
										assign node759 = (inp[2]) ? 13'b0000111111111 : node760;
											assign node760 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node764 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node767 = (inp[12]) ? node771 : node768;
										assign node768 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node771 = (inp[7]) ? 13'b0000001111111 : node772;
											assign node772 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node776 = (inp[2]) ? node784 : node777;
									assign node777 = (inp[9]) ? 13'b0000001111111 : node778;
										assign node778 = (inp[5]) ? node780 : 13'b0001111111111;
											assign node780 = (inp[12]) ? 13'b0000011111111 : 13'b0000011111111;
									assign node784 = (inp[5]) ? node786 : 13'b0000011111111;
										assign node786 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node789 = (inp[5]) ? node811 : node790;
								assign node790 = (inp[11]) ? node798 : node791;
									assign node791 = (inp[6]) ? node793 : 13'b0000011111111;
										assign node793 = (inp[12]) ? 13'b0000001111111 : node794;
											assign node794 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node798 = (inp[2]) ? node806 : node799;
										assign node799 = (inp[9]) ? node803 : node800;
											assign node800 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node803 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node806 = (inp[12]) ? 13'b0000000111111 : node807;
											assign node807 = (inp[7]) ? 13'b0000000111111 : 13'b0000000111111;
								assign node811 = (inp[7]) ? node819 : node812;
									assign node812 = (inp[9]) ? 13'b0000000111111 : node813;
										assign node813 = (inp[12]) ? 13'b0000000111111 : node814;
											assign node814 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node819 = (inp[9]) ? node825 : node820;
										assign node820 = (inp[6]) ? 13'b0000000011111 : node821;
											assign node821 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node825 = (inp[6]) ? node827 : 13'b0000000011111;
											assign node827 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node830 = (inp[5]) ? node904 : node831;
						assign node831 = (inp[6]) ? node871 : node832;
							assign node832 = (inp[8]) ? node856 : node833;
								assign node833 = (inp[9]) ? node841 : node834;
									assign node834 = (inp[11]) ? 13'b0000011111111 : node835;
										assign node835 = (inp[12]) ? 13'b0000011111111 : node836;
											assign node836 = (inp[0]) ? 13'b0000111111111 : 13'b0000111111111;
									assign node841 = (inp[7]) ? node849 : node842;
										assign node842 = (inp[2]) ? node846 : node843;
											assign node843 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node846 = (inp[12]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node849 = (inp[12]) ? node853 : node850;
											assign node850 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node853 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node856 = (inp[2]) ? node866 : node857;
									assign node857 = (inp[7]) ? 13'b0000001111111 : node858;
										assign node858 = (inp[9]) ? node862 : node859;
											assign node859 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node862 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node866 = (inp[7]) ? 13'b0000000111111 : node867;
										assign node867 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node871 = (inp[11]) ? node887 : node872;
								assign node872 = (inp[7]) ? node878 : node873;
									assign node873 = (inp[8]) ? 13'b0000001111111 : node874;
										assign node874 = (inp[12]) ? 13'b0000011111111 : 13'b0000001111111;
									assign node878 = (inp[8]) ? 13'b0000000111111 : node879;
										assign node879 = (inp[0]) ? node883 : node880;
											assign node880 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node883 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node887 = (inp[12]) ? node893 : node888;
									assign node888 = (inp[8]) ? 13'b0000000111111 : node889;
										assign node889 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node893 = (inp[9]) ? node899 : node894;
										assign node894 = (inp[0]) ? node896 : 13'b0000001111111;
											assign node896 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node899 = (inp[7]) ? node901 : 13'b0000000011111;
											assign node901 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node904 = (inp[2]) ? node950 : node905;
							assign node905 = (inp[11]) ? node925 : node906;
								assign node906 = (inp[9]) ? node914 : node907;
									assign node907 = (inp[12]) ? 13'b0000001111111 : node908;
										assign node908 = (inp[8]) ? 13'b0000011111111 : node909;
											assign node909 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node914 = (inp[0]) ? node920 : node915;
										assign node915 = (inp[6]) ? 13'b0000001111111 : node916;
											assign node916 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node920 = (inp[6]) ? node922 : 13'b0000001111111;
											assign node922 = (inp[12]) ? 13'b0000000111111 : 13'b0000000111111;
								assign node925 = (inp[8]) ? node937 : node926;
									assign node926 = (inp[12]) ? node932 : node927;
										assign node927 = (inp[6]) ? 13'b0000000111111 : node928;
											assign node928 = (inp[7]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node932 = (inp[6]) ? 13'b0000000011111 : node933;
											assign node933 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node937 = (inp[7]) ? node943 : node938;
										assign node938 = (inp[9]) ? node940 : 13'b0000001111111;
											assign node940 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node943 = (inp[6]) ? node947 : node944;
											assign node944 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node947 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
							assign node950 = (inp[8]) ? node970 : node951;
								assign node951 = (inp[12]) ? node963 : node952;
									assign node952 = (inp[0]) ? node958 : node953;
										assign node953 = (inp[7]) ? node955 : 13'b0000011111111;
											assign node955 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node958 = (inp[7]) ? 13'b0000000011111 : node959;
											assign node959 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node963 = (inp[9]) ? 13'b0000000011111 : node964;
										assign node964 = (inp[6]) ? node966 : 13'b0000000111111;
											assign node966 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node970 = (inp[12]) ? node986 : node971;
									assign node971 = (inp[6]) ? node979 : node972;
										assign node972 = (inp[11]) ? node976 : node973;
											assign node973 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node976 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node979 = (inp[0]) ? node983 : node980;
											assign node980 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node983 = (inp[11]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node986 = (inp[7]) ? node992 : node987;
										assign node987 = (inp[11]) ? node989 : 13'b0000000011111;
											assign node989 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node992 = (inp[0]) ? 13'b0000000000011 : node993;
											assign node993 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
				assign node997 = (inp[7]) ? node1139 : node998;
					assign node998 = (inp[5]) ? node1070 : node999;
						assign node999 = (inp[9]) ? node1031 : node1000;
							assign node1000 = (inp[12]) ? node1012 : node1001;
								assign node1001 = (inp[11]) ? node1007 : node1002;
									assign node1002 = (inp[0]) ? 13'b0000111111111 : node1003;
										assign node1003 = (inp[2]) ? 13'b0000111111111 : 13'b0011111111111;
									assign node1007 = (inp[8]) ? node1009 : 13'b0000011111111;
										assign node1009 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1012 = (inp[11]) ? node1022 : node1013;
									assign node1013 = (inp[2]) ? node1017 : node1014;
										assign node1014 = (inp[0]) ? 13'b0000111111111 : 13'b0000011111111;
										assign node1017 = (inp[8]) ? 13'b0000000111111 : node1018;
											assign node1018 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1022 = (inp[2]) ? node1028 : node1023;
										assign node1023 = (inp[0]) ? 13'b0000001111111 : node1024;
											assign node1024 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1028 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1031 = (inp[11]) ? node1049 : node1032;
								assign node1032 = (inp[1]) ? node1042 : node1033;
									assign node1033 = (inp[0]) ? node1039 : node1034;
										assign node1034 = (inp[6]) ? 13'b0000011111111 : node1035;
											assign node1035 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1039 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1042 = (inp[8]) ? node1044 : 13'b0000001111111;
										assign node1044 = (inp[12]) ? 13'b0000000001111 : node1045;
											assign node1045 = (inp[0]) ? 13'b0000001111111 : 13'b0000000111111;
								assign node1049 = (inp[12]) ? node1061 : node1050;
									assign node1050 = (inp[6]) ? node1056 : node1051;
										assign node1051 = (inp[0]) ? 13'b0000001111111 : node1052;
											assign node1052 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1056 = (inp[2]) ? 13'b0000000111111 : node1057;
											assign node1057 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1061 = (inp[2]) ? 13'b0000000011111 : node1062;
										assign node1062 = (inp[1]) ? node1066 : node1063;
											assign node1063 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1066 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node1070 = (inp[2]) ? node1104 : node1071;
							assign node1071 = (inp[1]) ? node1087 : node1072;
								assign node1072 = (inp[0]) ? node1080 : node1073;
									assign node1073 = (inp[8]) ? node1075 : 13'b0000111111111;
										assign node1075 = (inp[12]) ? 13'b0000011111111 : node1076;
											assign node1076 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1080 = (inp[8]) ? node1082 : 13'b0000001111111;
										assign node1082 = (inp[9]) ? 13'b0000000111111 : node1083;
											assign node1083 = (inp[6]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node1087 = (inp[9]) ? node1097 : node1088;
									assign node1088 = (inp[12]) ? node1092 : node1089;
										assign node1089 = (inp[8]) ? 13'b0000011111111 : 13'b0000001111111;
										assign node1092 = (inp[0]) ? 13'b0000000111111 : node1093;
											assign node1093 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1097 = (inp[12]) ? 13'b0000000111111 : node1098;
										assign node1098 = (inp[11]) ? node1100 : 13'b0000000111111;
											assign node1100 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1104 = (inp[11]) ? node1120 : node1105;
								assign node1105 = (inp[8]) ? node1113 : node1106;
									assign node1106 = (inp[9]) ? node1108 : 13'b0000001111111;
										assign node1108 = (inp[12]) ? 13'b0000000111111 : node1109;
											assign node1109 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1113 = (inp[9]) ? node1115 : 13'b0000000111111;
										assign node1115 = (inp[0]) ? node1117 : 13'b0000000111111;
											assign node1117 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1120 = (inp[12]) ? node1130 : node1121;
									assign node1121 = (inp[0]) ? node1127 : node1122;
										assign node1122 = (inp[8]) ? 13'b0000000111111 : node1123;
											assign node1123 = (inp[9]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node1127 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1130 = (inp[1]) ? 13'b0000000001111 : node1131;
										assign node1131 = (inp[6]) ? node1135 : node1132;
											assign node1132 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1135 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node1139 = (inp[8]) ? node1223 : node1140;
						assign node1140 = (inp[5]) ? node1182 : node1141;
							assign node1141 = (inp[12]) ? node1157 : node1142;
								assign node1142 = (inp[6]) ? node1152 : node1143;
									assign node1143 = (inp[1]) ? node1149 : node1144;
										assign node1144 = (inp[11]) ? node1146 : 13'b0000111111111;
											assign node1146 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1149 = (inp[2]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node1152 = (inp[0]) ? node1154 : 13'b0000001111111;
										assign node1154 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node1157 = (inp[6]) ? node1171 : node1158;
									assign node1158 = (inp[0]) ? node1166 : node1159;
										assign node1159 = (inp[2]) ? node1163 : node1160;
											assign node1160 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1163 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1166 = (inp[1]) ? 13'b0000000111111 : node1167;
											assign node1167 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1171 = (inp[9]) ? node1177 : node1172;
										assign node1172 = (inp[11]) ? 13'b0000000111111 : node1173;
											assign node1173 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1177 = (inp[1]) ? node1179 : 13'b0000000111111;
											assign node1179 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1182 = (inp[11]) ? node1194 : node1183;
								assign node1183 = (inp[1]) ? node1187 : node1184;
									assign node1184 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1187 = (inp[0]) ? node1189 : 13'b0000000111111;
										assign node1189 = (inp[6]) ? 13'b0000000011111 : node1190;
											assign node1190 = (inp[12]) ? 13'b0000000011111 : 13'b0000000011111;
								assign node1194 = (inp[9]) ? node1208 : node1195;
									assign node1195 = (inp[6]) ? node1201 : node1196;
										assign node1196 = (inp[1]) ? node1198 : 13'b0000000111111;
											assign node1198 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1201 = (inp[1]) ? node1205 : node1202;
											assign node1202 = (inp[2]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1205 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1208 = (inp[0]) ? node1216 : node1209;
										assign node1209 = (inp[2]) ? node1213 : node1210;
											assign node1210 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1213 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1216 = (inp[2]) ? node1220 : node1217;
											assign node1217 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1220 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node1223 = (inp[0]) ? node1261 : node1224;
							assign node1224 = (inp[12]) ? node1244 : node1225;
								assign node1225 = (inp[2]) ? node1231 : node1226;
									assign node1226 = (inp[1]) ? node1228 : 13'b0000001111111;
										assign node1228 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1231 = (inp[1]) ? node1239 : node1232;
										assign node1232 = (inp[6]) ? node1236 : node1233;
											assign node1233 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1236 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1239 = (inp[6]) ? node1241 : 13'b0000000011111;
											assign node1241 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1244 = (inp[2]) ? node1252 : node1245;
									assign node1245 = (inp[9]) ? node1247 : 13'b0000000111111;
										assign node1247 = (inp[6]) ? 13'b0000000011111 : node1248;
											assign node1248 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1252 = (inp[5]) ? 13'b0000000000111 : node1253;
										assign node1253 = (inp[1]) ? node1257 : node1254;
											assign node1254 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1257 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1261 = (inp[6]) ? node1275 : node1262;
								assign node1262 = (inp[12]) ? node1268 : node1263;
									assign node1263 = (inp[9]) ? node1265 : 13'b0000000111111;
										assign node1265 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1268 = (inp[1]) ? node1270 : 13'b0000000011111;
										assign node1270 = (inp[11]) ? node1272 : 13'b0000000011111;
											assign node1272 = (inp[2]) ? 13'b0000000000011 : 13'b0000000000111;
								assign node1275 = (inp[12]) ? node1289 : node1276;
									assign node1276 = (inp[9]) ? node1284 : node1277;
										assign node1277 = (inp[1]) ? node1281 : node1278;
											assign node1278 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node1281 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1284 = (inp[1]) ? node1286 : 13'b0000000001111;
											assign node1286 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node1289 = (inp[11]) ? node1297 : node1290;
										assign node1290 = (inp[1]) ? node1294 : node1291;
											assign node1291 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1294 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node1297 = (inp[1]) ? node1301 : node1298;
											assign node1298 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node1301 = (inp[2]) ? 13'b0000000000011 : 13'b0000000000111;
		assign node1304 = (inp[1]) ? node1970 : node1305;
			assign node1305 = (inp[12]) ? node1613 : node1306;
				assign node1306 = (inp[9]) ? node1454 : node1307;
					assign node1307 = (inp[6]) ? node1385 : node1308;
						assign node1308 = (inp[10]) ? node1350 : node1309;
							assign node1309 = (inp[11]) ? node1335 : node1310;
								assign node1310 = (inp[0]) ? node1324 : node1311;
									assign node1311 = (inp[7]) ? node1319 : node1312;
										assign node1312 = (inp[2]) ? node1316 : node1313;
											assign node1313 = (inp[5]) ? 13'b0011111111111 : 13'b0011111111111;
											assign node1316 = (inp[5]) ? 13'b0001111111111 : 13'b0001111111111;
										assign node1319 = (inp[5]) ? node1321 : 13'b0001111111111;
											assign node1321 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1324 = (inp[3]) ? node1332 : node1325;
										assign node1325 = (inp[8]) ? node1329 : node1326;
											assign node1326 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1329 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1332 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1335 = (inp[7]) ? node1345 : node1336;
									assign node1336 = (inp[5]) ? node1340 : node1337;
										assign node1337 = (inp[0]) ? 13'b0001111111111 : 13'b0000111111111;
										assign node1340 = (inp[2]) ? 13'b0000011111111 : node1341;
											assign node1341 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1345 = (inp[0]) ? 13'b0000001111111 : node1346;
										assign node1346 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node1350 = (inp[2]) ? node1368 : node1351;
								assign node1351 = (inp[11]) ? node1361 : node1352;
									assign node1352 = (inp[8]) ? node1358 : node1353;
										assign node1353 = (inp[0]) ? node1355 : 13'b0001111111111;
											assign node1355 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1358 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1361 = (inp[5]) ? node1363 : 13'b0000011111111;
										assign node1363 = (inp[0]) ? node1365 : 13'b0000111111111;
											assign node1365 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1368 = (inp[0]) ? node1376 : node1369;
									assign node1369 = (inp[3]) ? 13'b0000001111111 : node1370;
										assign node1370 = (inp[5]) ? 13'b0000001111111 : node1371;
											assign node1371 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1376 = (inp[5]) ? 13'b0000000111111 : node1377;
										assign node1377 = (inp[7]) ? node1381 : node1378;
											assign node1378 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1381 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node1385 = (inp[5]) ? node1417 : node1386;
							assign node1386 = (inp[8]) ? node1402 : node1387;
								assign node1387 = (inp[10]) ? node1397 : node1388;
									assign node1388 = (inp[3]) ? node1390 : 13'b0000111111111;
										assign node1390 = (inp[0]) ? node1394 : node1391;
											assign node1391 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1394 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1397 = (inp[2]) ? node1399 : 13'b0000011111111;
										assign node1399 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1402 = (inp[10]) ? node1412 : node1403;
									assign node1403 = (inp[0]) ? node1407 : node1404;
										assign node1404 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1407 = (inp[11]) ? 13'b0000000111111 : node1408;
											assign node1408 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1412 = (inp[3]) ? node1414 : 13'b0000001111111;
										assign node1414 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1417 = (inp[7]) ? node1431 : node1418;
								assign node1418 = (inp[8]) ? node1424 : node1419;
									assign node1419 = (inp[10]) ? node1421 : 13'b0000011111111;
										assign node1421 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1424 = (inp[10]) ? 13'b0000000111111 : node1425;
										assign node1425 = (inp[3]) ? node1427 : 13'b0000001111111;
											assign node1427 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1431 = (inp[0]) ? node1441 : node1432;
									assign node1432 = (inp[11]) ? node1436 : node1433;
										assign node1433 = (inp[3]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node1436 = (inp[10]) ? node1438 : 13'b0000000111111;
											assign node1438 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1441 = (inp[11]) ? node1449 : node1442;
										assign node1442 = (inp[8]) ? node1446 : node1443;
											assign node1443 = (inp[10]) ? 13'b0000001111111 : 13'b0000000111111;
											assign node1446 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1449 = (inp[2]) ? node1451 : 13'b0000000011111;
											assign node1451 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node1454 = (inp[5]) ? node1538 : node1455;
						assign node1455 = (inp[8]) ? node1499 : node1456;
							assign node1456 = (inp[0]) ? node1478 : node1457;
								assign node1457 = (inp[3]) ? node1467 : node1458;
									assign node1458 = (inp[6]) ? node1462 : node1459;
										assign node1459 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1462 = (inp[11]) ? 13'b0000001111111 : node1463;
											assign node1463 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1467 = (inp[10]) ? node1473 : node1468;
										assign node1468 = (inp[2]) ? node1470 : 13'b0000011111111;
											assign node1470 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1473 = (inp[11]) ? node1475 : 13'b0000001111111;
											assign node1475 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1478 = (inp[6]) ? node1488 : node1479;
									assign node1479 = (inp[2]) ? node1483 : node1480;
										assign node1480 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1483 = (inp[11]) ? 13'b0000001111111 : node1484;
											assign node1484 = (inp[10]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node1488 = (inp[3]) ? node1496 : node1489;
										assign node1489 = (inp[10]) ? node1493 : node1490;
											assign node1490 = (inp[11]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1493 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node1496 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1499 = (inp[2]) ? node1517 : node1500;
								assign node1500 = (inp[3]) ? node1506 : node1501;
									assign node1501 = (inp[0]) ? node1503 : 13'b0000011111111;
										assign node1503 = (inp[6]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node1506 = (inp[10]) ? node1512 : node1507;
										assign node1507 = (inp[0]) ? node1509 : 13'b0000011111111;
											assign node1509 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1512 = (inp[11]) ? 13'b0000000111111 : node1513;
											assign node1513 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1517 = (inp[11]) ? node1525 : node1518;
									assign node1518 = (inp[7]) ? node1520 : 13'b0000001111111;
										assign node1520 = (inp[10]) ? 13'b0000000111111 : node1521;
											assign node1521 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1525 = (inp[0]) ? node1531 : node1526;
										assign node1526 = (inp[3]) ? node1528 : 13'b0000001111111;
											assign node1528 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1531 = (inp[3]) ? node1535 : node1532;
											assign node1532 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1535 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node1538 = (inp[11]) ? node1570 : node1539;
							assign node1539 = (inp[8]) ? node1553 : node1540;
								assign node1540 = (inp[7]) ? node1544 : node1541;
									assign node1541 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1544 = (inp[2]) ? node1548 : node1545;
										assign node1545 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1548 = (inp[0]) ? 13'b0000000111111 : node1549;
											assign node1549 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1553 = (inp[2]) ? node1561 : node1554;
									assign node1554 = (inp[7]) ? 13'b0000000111111 : node1555;
										assign node1555 = (inp[3]) ? 13'b0000001111111 : node1556;
											assign node1556 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1561 = (inp[0]) ? node1567 : node1562;
										assign node1562 = (inp[7]) ? node1564 : 13'b0000000111111;
											assign node1564 = (inp[10]) ? 13'b0000000111111 : 13'b0000000011111;
										assign node1567 = (inp[10]) ? 13'b0000000011111 : 13'b0000000001111;
							assign node1570 = (inp[6]) ? node1590 : node1571;
								assign node1571 = (inp[0]) ? node1581 : node1572;
									assign node1572 = (inp[3]) ? node1576 : node1573;
										assign node1573 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1576 = (inp[7]) ? node1578 : 13'b0000000111111;
											assign node1578 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1581 = (inp[8]) ? node1587 : node1582;
										assign node1582 = (inp[7]) ? node1584 : 13'b0000011111111;
											assign node1584 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1587 = (inp[10]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node1590 = (inp[2]) ? node1602 : node1591;
									assign node1591 = (inp[3]) ? node1597 : node1592;
										assign node1592 = (inp[8]) ? node1594 : 13'b0000000111111;
											assign node1594 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1597 = (inp[8]) ? 13'b0000000011111 : node1598;
											assign node1598 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1602 = (inp[8]) ? node1610 : node1603;
										assign node1603 = (inp[10]) ? node1607 : node1604;
											assign node1604 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1607 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1610 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
				assign node1613 = (inp[11]) ? node1799 : node1614;
					assign node1614 = (inp[2]) ? node1696 : node1615;
						assign node1615 = (inp[0]) ? node1655 : node1616;
							assign node1616 = (inp[3]) ? node1632 : node1617;
								assign node1617 = (inp[6]) ? node1623 : node1618;
									assign node1618 = (inp[7]) ? node1620 : 13'b0000111111111;
										assign node1620 = (inp[8]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node1623 = (inp[7]) ? 13'b0000001111111 : node1624;
										assign node1624 = (inp[8]) ? node1628 : node1625;
											assign node1625 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1628 = (inp[5]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node1632 = (inp[8]) ? node1644 : node1633;
									assign node1633 = (inp[5]) ? node1639 : node1634;
										assign node1634 = (inp[9]) ? 13'b0000011111111 : node1635;
											assign node1635 = (inp[10]) ? 13'b0000011111111 : 13'b0001111111111;
										assign node1639 = (inp[9]) ? 13'b0000000111111 : node1640;
											assign node1640 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1644 = (inp[9]) ? node1650 : node1645;
										assign node1645 = (inp[5]) ? 13'b0000001111111 : node1646;
											assign node1646 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1650 = (inp[5]) ? 13'b0000000111111 : node1651;
											assign node1651 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1655 = (inp[3]) ? node1677 : node1656;
								assign node1656 = (inp[10]) ? node1672 : node1657;
									assign node1657 = (inp[7]) ? node1665 : node1658;
										assign node1658 = (inp[9]) ? node1662 : node1659;
											assign node1659 = (inp[8]) ? 13'b0000011111111 : 13'b0001111111111;
											assign node1662 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1665 = (inp[9]) ? node1669 : node1666;
											assign node1666 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1669 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1672 = (inp[7]) ? node1674 : 13'b0000001111111;
										assign node1674 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1677 = (inp[9]) ? node1687 : node1678;
									assign node1678 = (inp[7]) ? 13'b0000000111111 : node1679;
										assign node1679 = (inp[8]) ? node1683 : node1680;
											assign node1680 = (inp[10]) ? 13'b0000011111111 : 13'b0000001111111;
											assign node1683 = (inp[5]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1687 = (inp[10]) ? node1689 : 13'b0000000111111;
										assign node1689 = (inp[8]) ? node1693 : node1690;
											assign node1690 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1693 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1696 = (inp[7]) ? node1748 : node1697;
							assign node1697 = (inp[3]) ? node1725 : node1698;
								assign node1698 = (inp[5]) ? node1714 : node1699;
									assign node1699 = (inp[9]) ? node1707 : node1700;
										assign node1700 = (inp[6]) ? node1704 : node1701;
											assign node1701 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1704 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1707 = (inp[0]) ? node1711 : node1708;
											assign node1708 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1711 = (inp[10]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node1714 = (inp[0]) ? node1720 : node1715;
										assign node1715 = (inp[10]) ? 13'b0000000111111 : node1716;
											assign node1716 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1720 = (inp[10]) ? node1722 : 13'b0000000111111;
											assign node1722 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1725 = (inp[10]) ? node1739 : node1726;
									assign node1726 = (inp[8]) ? node1734 : node1727;
										assign node1727 = (inp[6]) ? node1731 : node1728;
											assign node1728 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1731 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1734 = (inp[9]) ? node1736 : 13'b0000000111111;
											assign node1736 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1739 = (inp[5]) ? node1743 : node1740;
										assign node1740 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1743 = (inp[6]) ? node1745 : 13'b0000000011111;
											assign node1745 = (inp[8]) ? 13'b0000000001111 : 13'b0000000001111;
							assign node1748 = (inp[6]) ? node1776 : node1749;
								assign node1749 = (inp[9]) ? node1763 : node1750;
									assign node1750 = (inp[10]) ? node1756 : node1751;
										assign node1751 = (inp[5]) ? node1753 : 13'b0000001111111;
											assign node1753 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1756 = (inp[3]) ? node1760 : node1757;
											assign node1757 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1760 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1763 = (inp[10]) ? node1769 : node1764;
										assign node1764 = (inp[0]) ? node1766 : 13'b0000000111111;
											assign node1766 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1769 = (inp[0]) ? node1773 : node1770;
											assign node1770 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1773 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1776 = (inp[5]) ? node1792 : node1777;
									assign node1777 = (inp[10]) ? node1785 : node1778;
										assign node1778 = (inp[8]) ? node1782 : node1779;
											assign node1779 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1782 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1785 = (inp[9]) ? node1789 : node1786;
											assign node1786 = (inp[0]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1789 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1792 = (inp[8]) ? 13'b0000000001111 : node1793;
										assign node1793 = (inp[3]) ? node1795 : 13'b0000000011111;
											assign node1795 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node1799 = (inp[8]) ? node1885 : node1800;
						assign node1800 = (inp[10]) ? node1834 : node1801;
							assign node1801 = (inp[0]) ? node1813 : node1802;
								assign node1802 = (inp[5]) ? node1804 : 13'b0000011111111;
									assign node1804 = (inp[7]) ? node1810 : node1805;
										assign node1805 = (inp[9]) ? 13'b0000000111111 : node1806;
											assign node1806 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1810 = (inp[9]) ? 13'b0000000111111 : 13'b0000000011111;
								assign node1813 = (inp[2]) ? node1825 : node1814;
									assign node1814 = (inp[3]) ? node1820 : node1815;
										assign node1815 = (inp[5]) ? 13'b0000001111111 : node1816;
											assign node1816 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1820 = (inp[5]) ? 13'b0000000111111 : node1821;
											assign node1821 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1825 = (inp[6]) ? 13'b0000000011111 : node1826;
										assign node1826 = (inp[7]) ? node1830 : node1827;
											assign node1827 = (inp[3]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1830 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1834 = (inp[5]) ? node1862 : node1835;
								assign node1835 = (inp[7]) ? node1851 : node1836;
									assign node1836 = (inp[2]) ? node1844 : node1837;
										assign node1837 = (inp[9]) ? node1841 : node1838;
											assign node1838 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1841 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1844 = (inp[3]) ? node1848 : node1845;
											assign node1845 = (inp[9]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1848 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1851 = (inp[6]) ? node1857 : node1852;
										assign node1852 = (inp[0]) ? 13'b0000000011111 : node1853;
											assign node1853 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1857 = (inp[9]) ? 13'b0000000000111 : node1858;
											assign node1858 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1862 = (inp[2]) ? node1876 : node1863;
									assign node1863 = (inp[0]) ? node1869 : node1864;
										assign node1864 = (inp[7]) ? node1866 : 13'b0000000111111;
											assign node1866 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1869 = (inp[6]) ? node1873 : node1870;
											assign node1870 = (inp[7]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1873 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1876 = (inp[0]) ? node1880 : node1877;
										assign node1877 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1880 = (inp[3]) ? 13'b0000000001111 : node1881;
											assign node1881 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1885 = (inp[7]) ? node1931 : node1886;
							assign node1886 = (inp[2]) ? node1912 : node1887;
								assign node1887 = (inp[5]) ? node1901 : node1888;
									assign node1888 = (inp[6]) ? node1894 : node1889;
										assign node1889 = (inp[9]) ? node1891 : 13'b0000001111111;
											assign node1891 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1894 = (inp[10]) ? node1898 : node1895;
											assign node1895 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1898 = (inp[9]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1901 = (inp[0]) ? node1909 : node1902;
										assign node1902 = (inp[3]) ? node1906 : node1903;
											assign node1903 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1906 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1909 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1912 = (inp[6]) ? node1922 : node1913;
									assign node1913 = (inp[3]) ? 13'b0000000011111 : node1914;
										assign node1914 = (inp[0]) ? node1918 : node1915;
											assign node1915 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1918 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1922 = (inp[9]) ? node1924 : 13'b0000000011111;
										assign node1924 = (inp[3]) ? node1928 : node1925;
											assign node1925 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1928 = (inp[0]) ? 13'b0000000000011 : 13'b0000000000111;
							assign node1931 = (inp[3]) ? node1951 : node1932;
								assign node1932 = (inp[10]) ? node1944 : node1933;
									assign node1933 = (inp[6]) ? node1937 : node1934;
										assign node1934 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1937 = (inp[2]) ? node1941 : node1938;
											assign node1938 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1941 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1944 = (inp[0]) ? 13'b0000000001111 : node1945;
										assign node1945 = (inp[2]) ? node1947 : 13'b0000000011111;
											assign node1947 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1951 = (inp[2]) ? node1959 : node1952;
									assign node1952 = (inp[5]) ? 13'b0000000001111 : node1953;
										assign node1953 = (inp[0]) ? 13'b0000000001111 : node1954;
											assign node1954 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1959 = (inp[0]) ? node1965 : node1960;
										assign node1960 = (inp[6]) ? node1962 : 13'b0000000001111;
											assign node1962 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node1965 = (inp[5]) ? node1967 : 13'b0000000000111;
											assign node1967 = (inp[9]) ? 13'b0000000000001 : 13'b0000000000011;
			assign node1970 = (inp[12]) ? node2308 : node1971;
				assign node1971 = (inp[10]) ? node2145 : node1972;
					assign node1972 = (inp[2]) ? node2056 : node1973;
						assign node1973 = (inp[8]) ? node2011 : node1974;
							assign node1974 = (inp[7]) ? node1992 : node1975;
								assign node1975 = (inp[11]) ? node1983 : node1976;
									assign node1976 = (inp[5]) ? node1978 : 13'b0000111111111;
										assign node1978 = (inp[0]) ? 13'b0000011111111 : node1979;
											assign node1979 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node1983 = (inp[3]) ? 13'b0000001111111 : node1984;
										assign node1984 = (inp[9]) ? node1988 : node1985;
											assign node1985 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1988 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1992 = (inp[11]) ? node2002 : node1993;
									assign node1993 = (inp[5]) ? node1997 : node1994;
										assign node1994 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1997 = (inp[3]) ? node1999 : 13'b0000011111111;
											assign node1999 = (inp[6]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node2002 = (inp[5]) ? node2008 : node2003;
										assign node2003 = (inp[9]) ? node2005 : 13'b0000011111111;
											assign node2005 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2008 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node2011 = (inp[0]) ? node2037 : node2012;
								assign node2012 = (inp[6]) ? node2028 : node2013;
									assign node2013 = (inp[11]) ? node2021 : node2014;
										assign node2014 = (inp[7]) ? node2018 : node2015;
											assign node2015 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2018 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2021 = (inp[7]) ? node2025 : node2022;
											assign node2022 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2025 = (inp[9]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node2028 = (inp[3]) ? 13'b0000000111111 : node2029;
										assign node2029 = (inp[7]) ? node2033 : node2030;
											assign node2030 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2033 = (inp[9]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node2037 = (inp[7]) ? node2049 : node2038;
									assign node2038 = (inp[9]) ? node2044 : node2039;
										assign node2039 = (inp[5]) ? 13'b0000000111111 : node2040;
											assign node2040 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2044 = (inp[6]) ? 13'b0000000111111 : node2045;
											assign node2045 = (inp[5]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node2049 = (inp[5]) ? node2051 : 13'b0000000111111;
										assign node2051 = (inp[6]) ? node2053 : 13'b0000000011111;
											assign node2053 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node2056 = (inp[11]) ? node2100 : node2057;
							assign node2057 = (inp[0]) ? node2075 : node2058;
								assign node2058 = (inp[7]) ? node2070 : node2059;
									assign node2059 = (inp[9]) ? node2065 : node2060;
										assign node2060 = (inp[5]) ? node2062 : 13'b0000111111111;
											assign node2062 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2065 = (inp[6]) ? 13'b0000000111111 : node2066;
											assign node2066 = (inp[5]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node2070 = (inp[5]) ? node2072 : 13'b0000001111111;
										assign node2072 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2075 = (inp[6]) ? node2089 : node2076;
									assign node2076 = (inp[5]) ? node2084 : node2077;
										assign node2077 = (inp[8]) ? node2081 : node2078;
											assign node2078 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2081 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2084 = (inp[9]) ? node2086 : 13'b0000001111111;
											assign node2086 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2089 = (inp[3]) ? node2095 : node2090;
										assign node2090 = (inp[7]) ? 13'b0000000111111 : node2091;
											assign node2091 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2095 = (inp[7]) ? node2097 : 13'b0000000111111;
											assign node2097 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2100 = (inp[8]) ? node2128 : node2101;
								assign node2101 = (inp[9]) ? node2113 : node2102;
									assign node2102 = (inp[0]) ? node2108 : node2103;
										assign node2103 = (inp[3]) ? node2105 : 13'b0000001111111;
											assign node2105 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2108 = (inp[7]) ? node2110 : 13'b0000000111111;
											assign node2110 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2113 = (inp[5]) ? node2121 : node2114;
										assign node2114 = (inp[7]) ? node2118 : node2115;
											assign node2115 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2118 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2121 = (inp[0]) ? node2125 : node2122;
											assign node2122 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2125 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node2128 = (inp[5]) ? node2138 : node2129;
									assign node2129 = (inp[3]) ? node2135 : node2130;
										assign node2130 = (inp[7]) ? node2132 : 13'b0000000111111;
											assign node2132 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2135 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2138 = (inp[0]) ? node2142 : node2139;
										assign node2139 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2142 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node2145 = (inp[9]) ? node2223 : node2146;
						assign node2146 = (inp[0]) ? node2182 : node2147;
							assign node2147 = (inp[11]) ? node2165 : node2148;
								assign node2148 = (inp[6]) ? node2158 : node2149;
									assign node2149 = (inp[7]) ? 13'b0000001111111 : node2150;
										assign node2150 = (inp[8]) ? node2154 : node2151;
											assign node2151 = (inp[2]) ? 13'b0000011111111 : 13'b0001111111111;
											assign node2154 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2158 = (inp[2]) ? node2160 : 13'b0000001111111;
										assign node2160 = (inp[8]) ? 13'b0000000111111 : node2161;
											assign node2161 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2165 = (inp[5]) ? node2175 : node2166;
									assign node2166 = (inp[6]) ? node2172 : node2167;
										assign node2167 = (inp[3]) ? node2169 : 13'b0000001111111;
											assign node2169 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2172 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2175 = (inp[2]) ? node2177 : 13'b0000000111111;
										assign node2177 = (inp[6]) ? 13'b0000000111111 : node2178;
											assign node2178 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2182 = (inp[3]) ? node2200 : node2183;
								assign node2183 = (inp[2]) ? node2195 : node2184;
									assign node2184 = (inp[8]) ? node2190 : node2185;
										assign node2185 = (inp[6]) ? node2187 : 13'b0000001111111;
											assign node2187 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2190 = (inp[7]) ? 13'b0000000111111 : node2191;
											assign node2191 = (inp[5]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node2195 = (inp[6]) ? node2197 : 13'b0000000111111;
										assign node2197 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2200 = (inp[8]) ? node2216 : node2201;
									assign node2201 = (inp[11]) ? node2209 : node2202;
										assign node2202 = (inp[5]) ? node2206 : node2203;
											assign node2203 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2206 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2209 = (inp[5]) ? node2213 : node2210;
											assign node2210 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2213 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2216 = (inp[6]) ? node2218 : 13'b0000000011111;
										assign node2218 = (inp[11]) ? node2220 : 13'b0000000001111;
											assign node2220 = (inp[2]) ? 13'b0000000000011 : 13'b0000000001111;
						assign node2223 = (inp[8]) ? node2271 : node2224;
							assign node2224 = (inp[2]) ? node2250 : node2225;
								assign node2225 = (inp[6]) ? node2239 : node2226;
									assign node2226 = (inp[0]) ? node2232 : node2227;
										assign node2227 = (inp[7]) ? node2229 : 13'b0000001111111;
											assign node2229 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2232 = (inp[3]) ? node2236 : node2233;
											assign node2233 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node2236 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2239 = (inp[11]) ? node2245 : node2240;
										assign node2240 = (inp[0]) ? node2242 : 13'b0000000111111;
											assign node2242 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2245 = (inp[7]) ? node2247 : 13'b0000000011111;
											assign node2247 = (inp[5]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node2250 = (inp[3]) ? node2262 : node2251;
									assign node2251 = (inp[5]) ? node2255 : node2252;
										assign node2252 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2255 = (inp[0]) ? node2259 : node2256;
											assign node2256 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2259 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2262 = (inp[7]) ? node2266 : node2263;
										assign node2263 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2266 = (inp[6]) ? 13'b0000000001111 : node2267;
											assign node2267 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2271 = (inp[6]) ? node2293 : node2272;
								assign node2272 = (inp[3]) ? node2282 : node2273;
									assign node2273 = (inp[0]) ? node2279 : node2274;
										assign node2274 = (inp[5]) ? 13'b0000000011111 : node2275;
											assign node2275 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node2279 = (inp[7]) ? 13'b0000000011111 : 13'b0000000001111;
									assign node2282 = (inp[11]) ? node2286 : node2283;
										assign node2283 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2286 = (inp[5]) ? node2290 : node2287;
											assign node2287 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2290 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node2293 = (inp[2]) ? node2301 : node2294;
									assign node2294 = (inp[5]) ? node2296 : 13'b0000000011111;
										assign node2296 = (inp[11]) ? 13'b0000000001111 : node2297;
											assign node2297 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2301 = (inp[11]) ? node2303 : 13'b0000000001111;
										assign node2303 = (inp[7]) ? 13'b0000000000001 : node2304;
											assign node2304 = (inp[0]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node2308 = (inp[8]) ? node2482 : node2309;
					assign node2309 = (inp[5]) ? node2387 : node2310;
						assign node2310 = (inp[0]) ? node2356 : node2311;
							assign node2311 = (inp[11]) ? node2335 : node2312;
								assign node2312 = (inp[2]) ? node2326 : node2313;
									assign node2313 = (inp[6]) ? node2321 : node2314;
										assign node2314 = (inp[3]) ? node2318 : node2315;
											assign node2315 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2318 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2321 = (inp[7]) ? node2323 : 13'b0000011111111;
											assign node2323 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2326 = (inp[9]) ? node2332 : node2327;
										assign node2327 = (inp[6]) ? 13'b0000001111111 : node2328;
											assign node2328 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2332 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2335 = (inp[3]) ? node2347 : node2336;
									assign node2336 = (inp[7]) ? node2342 : node2337;
										assign node2337 = (inp[9]) ? 13'b0000001111111 : node2338;
											assign node2338 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2342 = (inp[6]) ? 13'b0000000011111 : node2343;
											assign node2343 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2347 = (inp[7]) ? node2349 : 13'b0000000111111;
										assign node2349 = (inp[2]) ? node2353 : node2350;
											assign node2350 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2353 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2356 = (inp[9]) ? node2370 : node2357;
								assign node2357 = (inp[11]) ? node2363 : node2358;
									assign node2358 = (inp[7]) ? 13'b0000000111111 : node2359;
										assign node2359 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2363 = (inp[2]) ? node2365 : 13'b0000000111111;
										assign node2365 = (inp[6]) ? 13'b0000000001111 : node2366;
											assign node2366 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2370 = (inp[3]) ? node2382 : node2371;
									assign node2371 = (inp[7]) ? node2377 : node2372;
										assign node2372 = (inp[10]) ? 13'b0000000111111 : node2373;
											assign node2373 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2377 = (inp[10]) ? 13'b0000000001111 : node2378;
											assign node2378 = (inp[6]) ? 13'b0000000111111 : 13'b0000000011111;
									assign node2382 = (inp[2]) ? node2384 : 13'b0000000011111;
										assign node2384 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node2387 = (inp[11]) ? node2439 : node2388;
							assign node2388 = (inp[7]) ? node2416 : node2389;
								assign node2389 = (inp[9]) ? node2403 : node2390;
									assign node2390 = (inp[0]) ? node2398 : node2391;
										assign node2391 = (inp[3]) ? node2395 : node2392;
											assign node2392 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2395 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2398 = (inp[3]) ? node2400 : 13'b0000000111111;
											assign node2400 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2403 = (inp[10]) ? node2411 : node2404;
										assign node2404 = (inp[2]) ? node2408 : node2405;
											assign node2405 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2408 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node2411 = (inp[2]) ? node2413 : 13'b0000000011111;
											assign node2413 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2416 = (inp[9]) ? node2426 : node2417;
									assign node2417 = (inp[0]) ? node2421 : node2418;
										assign node2418 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2421 = (inp[6]) ? node2423 : 13'b0000000111111;
											assign node2423 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2426 = (inp[2]) ? node2434 : node2427;
										assign node2427 = (inp[0]) ? node2431 : node2428;
											assign node2428 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2431 = (inp[3]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node2434 = (inp[6]) ? node2436 : 13'b0000000001111;
											assign node2436 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node2439 = (inp[0]) ? node2461 : node2440;
								assign node2440 = (inp[2]) ? node2452 : node2441;
									assign node2441 = (inp[10]) ? node2447 : node2442;
										assign node2442 = (inp[7]) ? node2444 : 13'b0000000111111;
											assign node2444 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2447 = (inp[9]) ? node2449 : 13'b0000000011111;
											assign node2449 = (inp[3]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node2452 = (inp[10]) ? 13'b0000000001111 : node2453;
										assign node2453 = (inp[7]) ? node2457 : node2454;
											assign node2454 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2457 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2461 = (inp[3]) ? node2473 : node2462;
									assign node2462 = (inp[6]) ? node2468 : node2463;
										assign node2463 = (inp[2]) ? 13'b0000000011111 : node2464;
											assign node2464 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2468 = (inp[2]) ? 13'b0000000000111 : node2469;
											assign node2469 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2473 = (inp[2]) ? node2477 : node2474;
										assign node2474 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2477 = (inp[9]) ? node2479 : 13'b0000000000111;
											assign node2479 = (inp[6]) ? 13'b0000000000001 : 13'b0000000000111;
					assign node2482 = (inp[11]) ? node2578 : node2483;
						assign node2483 = (inp[10]) ? node2521 : node2484;
							assign node2484 = (inp[0]) ? node2500 : node2485;
								assign node2485 = (inp[9]) ? node2495 : node2486;
									assign node2486 = (inp[2]) ? 13'b0000000111111 : node2487;
										assign node2487 = (inp[6]) ? node2491 : node2488;
											assign node2488 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2491 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2495 = (inp[6]) ? node2497 : 13'b0000000111111;
										assign node2497 = (inp[7]) ? 13'b0000000011111 : 13'b0000000001111;
								assign node2500 = (inp[6]) ? node2512 : node2501;
									assign node2501 = (inp[2]) ? node2505 : node2502;
										assign node2502 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2505 = (inp[9]) ? node2509 : node2506;
											assign node2506 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2509 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2512 = (inp[5]) ? node2514 : 13'b0000000011111;
										assign node2514 = (inp[9]) ? node2518 : node2515;
											assign node2515 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2518 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node2521 = (inp[3]) ? node2551 : node2522;
								assign node2522 = (inp[9]) ? node2538 : node2523;
									assign node2523 = (inp[2]) ? node2531 : node2524;
										assign node2524 = (inp[6]) ? node2528 : node2525;
											assign node2525 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2528 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2531 = (inp[0]) ? node2535 : node2532;
											assign node2532 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2535 = (inp[5]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node2538 = (inp[6]) ? node2544 : node2539;
										assign node2539 = (inp[0]) ? node2541 : 13'b0000000011111;
											assign node2541 = (inp[2]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node2544 = (inp[2]) ? node2548 : node2545;
											assign node2545 = (inp[5]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2548 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node2551 = (inp[0]) ? node2563 : node2552;
									assign node2552 = (inp[5]) ? node2558 : node2553;
										assign node2553 = (inp[2]) ? 13'b0000000001111 : node2554;
											assign node2554 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node2558 = (inp[9]) ? 13'b0000000001111 : node2559;
											assign node2559 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node2563 = (inp[5]) ? node2571 : node2564;
										assign node2564 = (inp[6]) ? node2568 : node2565;
											assign node2565 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2568 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2571 = (inp[9]) ? node2575 : node2572;
											assign node2572 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node2575 = (inp[6]) ? 13'b0000000000001 : 13'b0000000000011;
						assign node2578 = (inp[5]) ? node2630 : node2579;
							assign node2579 = (inp[9]) ? node2607 : node2580;
								assign node2580 = (inp[3]) ? node2592 : node2581;
									assign node2581 = (inp[0]) ? node2587 : node2582;
										assign node2582 = (inp[10]) ? 13'b0000000111111 : node2583;
											assign node2583 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2587 = (inp[7]) ? node2589 : 13'b0000000011111;
											assign node2589 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node2592 = (inp[7]) ? node2600 : node2593;
										assign node2593 = (inp[6]) ? node2597 : node2594;
											assign node2594 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2597 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2600 = (inp[10]) ? node2604 : node2601;
											assign node2601 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2604 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node2607 = (inp[3]) ? node2619 : node2608;
									assign node2608 = (inp[0]) ? node2614 : node2609;
										assign node2609 = (inp[10]) ? 13'b0000000001111 : node2610;
											assign node2610 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2614 = (inp[7]) ? 13'b0000000000111 : node2615;
											assign node2615 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2619 = (inp[6]) ? node2623 : node2620;
										assign node2620 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2623 = (inp[7]) ? node2627 : node2624;
											assign node2624 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node2627 = (inp[2]) ? 13'b0000000000011 : 13'b0000000000111;
							assign node2630 = (inp[9]) ? node2652 : node2631;
								assign node2631 = (inp[7]) ? node2639 : node2632;
									assign node2632 = (inp[10]) ? node2634 : 13'b0000000011111;
										assign node2634 = (inp[2]) ? 13'b0000000000111 : node2635;
											assign node2635 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2639 = (inp[3]) ? node2647 : node2640;
										assign node2640 = (inp[0]) ? node2644 : node2641;
											assign node2641 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2644 = (inp[2]) ? 13'b0000000000011 : 13'b0000000001111;
										assign node2647 = (inp[6]) ? node2649 : 13'b0000000000111;
											assign node2649 = (inp[0]) ? 13'b0000000000011 : 13'b0000000000111;
								assign node2652 = (inp[2]) ? node2660 : node2653;
									assign node2653 = (inp[10]) ? 13'b0000000000111 : node2654;
										assign node2654 = (inp[7]) ? node2656 : 13'b0000000001111;
											assign node2656 = (inp[3]) ? 13'b0000000000111 : 13'b0000000000111;
									assign node2660 = (inp[6]) ? node2668 : node2661;
										assign node2661 = (inp[0]) ? node2665 : node2662;
											assign node2662 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node2665 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000111;
										assign node2668 = (inp[3]) ? 13'b0000000000001 : node2669;
											assign node2669 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;

endmodule