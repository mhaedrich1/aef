module dtc_split5_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node3;
	wire [40-1:0] node4;
	wire [40-1:0] node6;
	wire [40-1:0] node8;
	wire [40-1:0] node10;
	wire [40-1:0] node15;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node50;
	wire [40-1:0] node52;
	wire [40-1:0] node53;
	wire [40-1:0] node55;
	wire [40-1:0] node56;
	wire [40-1:0] node58;
	wire [40-1:0] node61;
	wire [40-1:0] node63;
	wire [40-1:0] node67;
	wire [40-1:0] node68;
	wire [40-1:0] node70;
	wire [40-1:0] node72;
	wire [40-1:0] node73;
	wire [40-1:0] node74;
	wire [40-1:0] node77;
	wire [40-1:0] node80;
	wire [40-1:0] node82;
	wire [40-1:0] node85;
	wire [40-1:0] node86;
	wire [40-1:0] node87;
	wire [40-1:0] node89;
	wire [40-1:0] node90;
	wire [40-1:0] node95;
	wire [40-1:0] node97;
	wire [40-1:0] node99;
	wire [40-1:0] node100;
	wire [40-1:0] node104;
	wire [40-1:0] node105;
	wire [40-1:0] node108;
	wire [40-1:0] node109;
	wire [40-1:0] node111;
	wire [40-1:0] node113;
	wire [40-1:0] node115;
	wire [40-1:0] node117;
	wire [40-1:0] node119;
	wire [40-1:0] node122;
	wire [40-1:0] node123;
	wire [40-1:0] node125;
	wire [40-1:0] node127;
	wire [40-1:0] node128;
	wire [40-1:0] node130;
	wire [40-1:0] node133;
	wire [40-1:0] node134;
	wire [40-1:0] node137;
	wire [40-1:0] node140;
	wire [40-1:0] node141;
	wire [40-1:0] node143;
	wire [40-1:0] node145;
	wire [40-1:0] node147;
	wire [40-1:0] node150;
	wire [40-1:0] node153;
	wire [40-1:0] node154;
	wire [40-1:0] node155;
	wire [40-1:0] node157;
	wire [40-1:0] node159;
	wire [40-1:0] node160;
	wire [40-1:0] node162;
	wire [40-1:0] node164;
	wire [40-1:0] node166;
	wire [40-1:0] node167;
	wire [40-1:0] node170;
	wire [40-1:0] node173;
	wire [40-1:0] node174;
	wire [40-1:0] node176;
	wire [40-1:0] node178;
	wire [40-1:0] node179;
	wire [40-1:0] node183;
	wire [40-1:0] node187;
	wire [40-1:0] node188;
	wire [40-1:0] node190;
	wire [40-1:0] node192;
	wire [40-1:0] node193;
	wire [40-1:0] node195;
	wire [40-1:0] node198;
	wire [40-1:0] node199;
	wire [40-1:0] node202;
	wire [40-1:0] node205;
	wire [40-1:0] node206;
	wire [40-1:0] node209;
	wire [40-1:0] node210;
	wire [40-1:0] node212;
	wire [40-1:0] node214;
	wire [40-1:0] node216;
	wire [40-1:0] node217;
	wire [40-1:0] node219;
	wire [40-1:0] node222;
	wire [40-1:0] node224;
	wire [40-1:0] node227;
	wire [40-1:0] node228;
	wire [40-1:0] node230;
	wire [40-1:0] node232;
	wire [40-1:0] node233;
	wire [40-1:0] node235;
	wire [40-1:0] node238;
	wire [40-1:0] node239;
	wire [40-1:0] node242;
	wire [40-1:0] node245;
	wire [40-1:0] node246;
	wire [40-1:0] node248;
	wire [40-1:0] node250;
	wire [40-1:0] node251;
	wire [40-1:0] node254;
	wire [40-1:0] node257;
	wire [40-1:0] node260;
	wire [40-1:0] node261;
	wire [40-1:0] node262;
	wire [40-1:0] node265;
	wire [40-1:0] node266;
	wire [40-1:0] node267;
	wire [40-1:0] node268;
	wire [40-1:0] node269;
	wire [40-1:0] node272;
	wire [40-1:0] node275;
	wire [40-1:0] node276;
	wire [40-1:0] node279;
	wire [40-1:0] node282;
	wire [40-1:0] node283;
	wire [40-1:0] node284;
	wire [40-1:0] node287;
	wire [40-1:0] node290;
	wire [40-1:0] node291;
	wire [40-1:0] node294;
	wire [40-1:0] node297;
	wire [40-1:0] node298;
	wire [40-1:0] node299;
	wire [40-1:0] node300;
	wire [40-1:0] node303;
	wire [40-1:0] node306;
	wire [40-1:0] node307;
	wire [40-1:0] node310;
	wire [40-1:0] node313;
	wire [40-1:0] node314;
	wire [40-1:0] node315;
	wire [40-1:0] node318;
	wire [40-1:0] node321;
	wire [40-1:0] node322;
	wire [40-1:0] node325;
	wire [40-1:0] node328;
	wire [40-1:0] node329;
	wire [40-1:0] node332;
	wire [40-1:0] node334;
	wire [40-1:0] node335;
	wire [40-1:0] node336;
	wire [40-1:0] node337;
	wire [40-1:0] node338;
	wire [40-1:0] node339;
	wire [40-1:0] node340;
	wire [40-1:0] node341;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node346;
	wire [40-1:0] node349;
	wire [40-1:0] node350;
	wire [40-1:0] node353;
	wire [40-1:0] node356;
	wire [40-1:0] node357;
	wire [40-1:0] node358;
	wire [40-1:0] node361;
	wire [40-1:0] node364;
	wire [40-1:0] node366;
	wire [40-1:0] node369;
	wire [40-1:0] node370;
	wire [40-1:0] node371;
	wire [40-1:0] node372;
	wire [40-1:0] node375;
	wire [40-1:0] node378;
	wire [40-1:0] node379;
	wire [40-1:0] node382;
	wire [40-1:0] node385;
	wire [40-1:0] node386;
	wire [40-1:0] node387;
	wire [40-1:0] node390;
	wire [40-1:0] node393;
	wire [40-1:0] node394;
	wire [40-1:0] node397;
	wire [40-1:0] node400;
	wire [40-1:0] node401;
	wire [40-1:0] node402;
	wire [40-1:0] node403;
	wire [40-1:0] node404;
	wire [40-1:0] node407;
	wire [40-1:0] node410;
	wire [40-1:0] node411;
	wire [40-1:0] node414;
	wire [40-1:0] node417;
	wire [40-1:0] node418;
	wire [40-1:0] node419;
	wire [40-1:0] node422;
	wire [40-1:0] node425;
	wire [40-1:0] node426;
	wire [40-1:0] node429;
	wire [40-1:0] node432;
	wire [40-1:0] node433;
	wire [40-1:0] node434;
	wire [40-1:0] node435;
	wire [40-1:0] node438;
	wire [40-1:0] node441;
	wire [40-1:0] node442;
	wire [40-1:0] node445;
	wire [40-1:0] node448;
	wire [40-1:0] node449;
	wire [40-1:0] node450;
	wire [40-1:0] node453;
	wire [40-1:0] node456;
	wire [40-1:0] node457;
	wire [40-1:0] node460;
	wire [40-1:0] node463;
	wire [40-1:0] node464;
	wire [40-1:0] node465;
	wire [40-1:0] node466;
	wire [40-1:0] node467;
	wire [40-1:0] node468;
	wire [40-1:0] node472;
	wire [40-1:0] node473;
	wire [40-1:0] node476;
	wire [40-1:0] node479;
	wire [40-1:0] node480;
	wire [40-1:0] node481;
	wire [40-1:0] node484;
	wire [40-1:0] node487;
	wire [40-1:0] node488;
	wire [40-1:0] node491;
	wire [40-1:0] node494;
	wire [40-1:0] node495;
	wire [40-1:0] node496;
	wire [40-1:0] node497;
	wire [40-1:0] node500;
	wire [40-1:0] node503;
	wire [40-1:0] node504;
	wire [40-1:0] node507;
	wire [40-1:0] node510;
	wire [40-1:0] node511;
	wire [40-1:0] node512;
	wire [40-1:0] node515;
	wire [40-1:0] node518;
	wire [40-1:0] node519;
	wire [40-1:0] node522;
	wire [40-1:0] node525;
	wire [40-1:0] node526;
	wire [40-1:0] node527;
	wire [40-1:0] node528;
	wire [40-1:0] node529;
	wire [40-1:0] node532;
	wire [40-1:0] node535;
	wire [40-1:0] node536;
	wire [40-1:0] node539;
	wire [40-1:0] node542;
	wire [40-1:0] node543;
	wire [40-1:0] node544;
	wire [40-1:0] node547;
	wire [40-1:0] node550;
	wire [40-1:0] node551;
	wire [40-1:0] node554;
	wire [40-1:0] node557;
	wire [40-1:0] node558;
	wire [40-1:0] node559;
	wire [40-1:0] node561;
	wire [40-1:0] node564;
	wire [40-1:0] node566;
	wire [40-1:0] node569;
	wire [40-1:0] node570;
	wire [40-1:0] node571;
	wire [40-1:0] node574;
	wire [40-1:0] node577;
	wire [40-1:0] node578;
	wire [40-1:0] node581;
	wire [40-1:0] node584;
	wire [40-1:0] node585;
	wire [40-1:0] node586;
	wire [40-1:0] node587;
	wire [40-1:0] node588;
	wire [40-1:0] node589;
	wire [40-1:0] node591;
	wire [40-1:0] node594;
	wire [40-1:0] node600;
	wire [40-1:0] node601;
	wire [40-1:0] node602;
	wire [40-1:0] node603;
	wire [40-1:0] node604;
	wire [40-1:0] node605;
	wire [40-1:0] node608;
	wire [40-1:0] node611;
	wire [40-1:0] node612;
	wire [40-1:0] node615;
	wire [40-1:0] node618;
	wire [40-1:0] node619;
	wire [40-1:0] node620;
	wire [40-1:0] node623;
	wire [40-1:0] node626;
	wire [40-1:0] node627;
	wire [40-1:0] node630;
	wire [40-1:0] node633;
	wire [40-1:0] node634;
	wire [40-1:0] node635;
	wire [40-1:0] node636;
	wire [40-1:0] node639;
	wire [40-1:0] node642;
	wire [40-1:0] node643;
	wire [40-1:0] node646;
	wire [40-1:0] node649;
	wire [40-1:0] node650;
	wire [40-1:0] node651;
	wire [40-1:0] node654;
	wire [40-1:0] node657;
	wire [40-1:0] node658;
	wire [40-1:0] node661;
	wire [40-1:0] node664;
	wire [40-1:0] node665;
	wire [40-1:0] node666;
	wire [40-1:0] node667;
	wire [40-1:0] node668;
	wire [40-1:0] node671;
	wire [40-1:0] node674;
	wire [40-1:0] node675;
	wire [40-1:0] node678;
	wire [40-1:0] node681;
	wire [40-1:0] node682;
	wire [40-1:0] node683;
	wire [40-1:0] node686;
	wire [40-1:0] node689;
	wire [40-1:0] node690;
	wire [40-1:0] node693;
	wire [40-1:0] node696;
	wire [40-1:0] node697;
	wire [40-1:0] node698;
	wire [40-1:0] node699;
	wire [40-1:0] node702;
	wire [40-1:0] node705;
	wire [40-1:0] node706;
	wire [40-1:0] node709;
	wire [40-1:0] node712;
	wire [40-1:0] node713;
	wire [40-1:0] node714;
	wire [40-1:0] node717;
	wire [40-1:0] node720;
	wire [40-1:0] node722;
	wire [40-1:0] node725;
	wire [40-1:0] node726;
	wire [40-1:0] node727;
	wire [40-1:0] node728;
	wire [40-1:0] node729;
	wire [40-1:0] node730;
	wire [40-1:0] node732;
	wire [40-1:0] node733;
	wire [40-1:0] node736;
	wire [40-1:0] node739;
	wire [40-1:0] node740;
	wire [40-1:0] node741;
	wire [40-1:0] node744;
	wire [40-1:0] node748;
	wire [40-1:0] node749;
	wire [40-1:0] node751;
	wire [40-1:0] node752;
	wire [40-1:0] node755;
	wire [40-1:0] node758;
	wire [40-1:0] node759;
	wire [40-1:0] node760;
	wire [40-1:0] node765;
	wire [40-1:0] node766;
	wire [40-1:0] node767;
	wire [40-1:0] node768;
	wire [40-1:0] node770;
	wire [40-1:0] node776;
	wire [40-1:0] node778;
	wire [40-1:0] node780;
	wire [40-1:0] node781;
	wire [40-1:0] node783;
	wire [40-1:0] node784;
	wire [40-1:0] node787;
	wire [40-1:0] node791;
	wire [40-1:0] node793;
	wire [40-1:0] node794;
	wire [40-1:0] node795;
	wire [40-1:0] node796;
	wire [40-1:0] node797;
	wire [40-1:0] node799;
	wire [40-1:0] node802;
	wire [40-1:0] node804;
	wire [40-1:0] node807;
	wire [40-1:0] node808;
	wire [40-1:0] node809;
	wire [40-1:0] node812;
	wire [40-1:0] node815;
	wire [40-1:0] node816;
	wire [40-1:0] node819;
	wire [40-1:0] node822;
	wire [40-1:0] node823;
	wire [40-1:0] node824;
	wire [40-1:0] node825;
	wire [40-1:0] node828;
	wire [40-1:0] node831;
	wire [40-1:0] node832;
	wire [40-1:0] node835;
	wire [40-1:0] node838;
	wire [40-1:0] node839;
	wire [40-1:0] node840;
	wire [40-1:0] node843;
	wire [40-1:0] node846;
	wire [40-1:0] node847;
	wire [40-1:0] node850;
	wire [40-1:0] node853;
	wire [40-1:0] node854;
	wire [40-1:0] node855;
	wire [40-1:0] node856;
	wire [40-1:0] node857;
	wire [40-1:0] node860;
	wire [40-1:0] node863;
	wire [40-1:0] node864;
	wire [40-1:0] node867;
	wire [40-1:0] node870;
	wire [40-1:0] node871;
	wire [40-1:0] node872;
	wire [40-1:0] node875;
	wire [40-1:0] node878;
	wire [40-1:0] node879;
	wire [40-1:0] node882;
	wire [40-1:0] node885;
	wire [40-1:0] node886;
	wire [40-1:0] node887;
	wire [40-1:0] node888;
	wire [40-1:0] node891;
	wire [40-1:0] node894;
	wire [40-1:0] node895;
	wire [40-1:0] node898;
	wire [40-1:0] node901;
	wire [40-1:0] node902;
	wire [40-1:0] node903;
	wire [40-1:0] node906;
	wire [40-1:0] node909;
	wire [40-1:0] node910;
	wire [40-1:0] node913;
	wire [40-1:0] node916;
	wire [40-1:0] node917;
	wire [40-1:0] node918;
	wire [40-1:0] node920;
	wire [40-1:0] node921;
	wire [40-1:0] node922;
	wire [40-1:0] node924;
	wire [40-1:0] node927;
	wire [40-1:0] node928;
	wire [40-1:0] node932;
	wire [40-1:0] node933;
	wire [40-1:0] node935;
	wire [40-1:0] node938;
	wire [40-1:0] node939;
	wire [40-1:0] node943;
	wire [40-1:0] node944;
	wire [40-1:0] node945;
	wire [40-1:0] node947;
	wire [40-1:0] node949;
	wire [40-1:0] node951;
	wire [40-1:0] node953;
	wire [40-1:0] node956;
	wire [40-1:0] node957;
	wire [40-1:0] node959;
	wire [40-1:0] node961;
	wire [40-1:0] node962;
	wire [40-1:0] node965;
	wire [40-1:0] node968;
	wire [40-1:0] node969;
	wire [40-1:0] node971;
	wire [40-1:0] node972;
	wire [40-1:0] node975;
	wire [40-1:0] node978;
	wire [40-1:0] node979;
	wire [40-1:0] node980;
	wire [40-1:0] node983;
	wire [40-1:0] node988;
	wire [40-1:0] node989;
	wire [40-1:0] node991;
	wire [40-1:0] node992;
	wire [40-1:0] node993;
	wire [40-1:0] node994;
	wire [40-1:0] node995;
	wire [40-1:0] node996;
	wire [40-1:0] node999;
	wire [40-1:0] node1002;
	wire [40-1:0] node1003;
	wire [40-1:0] node1006;
	wire [40-1:0] node1009;
	wire [40-1:0] node1010;
	wire [40-1:0] node1011;
	wire [40-1:0] node1014;
	wire [40-1:0] node1017;
	wire [40-1:0] node1018;
	wire [40-1:0] node1021;
	wire [40-1:0] node1024;
	wire [40-1:0] node1025;
	wire [40-1:0] node1026;
	wire [40-1:0] node1027;
	wire [40-1:0] node1030;
	wire [40-1:0] node1033;
	wire [40-1:0] node1034;
	wire [40-1:0] node1037;
	wire [40-1:0] node1040;
	wire [40-1:0] node1041;
	wire [40-1:0] node1042;
	wire [40-1:0] node1045;
	wire [40-1:0] node1048;
	wire [40-1:0] node1049;
	wire [40-1:0] node1052;
	wire [40-1:0] node1055;
	wire [40-1:0] node1056;
	wire [40-1:0] node1057;
	wire [40-1:0] node1058;
	wire [40-1:0] node1059;
	wire [40-1:0] node1062;
	wire [40-1:0] node1065;
	wire [40-1:0] node1066;
	wire [40-1:0] node1069;
	wire [40-1:0] node1072;
	wire [40-1:0] node1073;
	wire [40-1:0] node1074;
	wire [40-1:0] node1077;
	wire [40-1:0] node1080;
	wire [40-1:0] node1081;
	wire [40-1:0] node1084;
	wire [40-1:0] node1087;
	wire [40-1:0] node1088;
	wire [40-1:0] node1089;
	wire [40-1:0] node1090;
	wire [40-1:0] node1093;
	wire [40-1:0] node1096;
	wire [40-1:0] node1097;
	wire [40-1:0] node1100;
	wire [40-1:0] node1103;
	wire [40-1:0] node1104;
	wire [40-1:0] node1105;
	wire [40-1:0] node1108;
	wire [40-1:0] node1111;
	wire [40-1:0] node1112;
	wire [40-1:0] node1115;
	wire [40-1:0] node1118;
	wire [40-1:0] node1119;
	wire [40-1:0] node1120;
	wire [40-1:0] node1121;
	wire [40-1:0] node1122;
	wire [40-1:0] node1123;
	wire [40-1:0] node1124;
	wire [40-1:0] node1127;
	wire [40-1:0] node1130;
	wire [40-1:0] node1131;
	wire [40-1:0] node1134;
	wire [40-1:0] node1137;
	wire [40-1:0] node1138;
	wire [40-1:0] node1139;
	wire [40-1:0] node1142;
	wire [40-1:0] node1145;
	wire [40-1:0] node1146;
	wire [40-1:0] node1149;
	wire [40-1:0] node1152;
	wire [40-1:0] node1153;
	wire [40-1:0] node1154;
	wire [40-1:0] node1155;
	wire [40-1:0] node1158;
	wire [40-1:0] node1161;
	wire [40-1:0] node1162;
	wire [40-1:0] node1165;
	wire [40-1:0] node1168;
	wire [40-1:0] node1169;
	wire [40-1:0] node1170;
	wire [40-1:0] node1173;
	wire [40-1:0] node1176;
	wire [40-1:0] node1177;
	wire [40-1:0] node1180;
	wire [40-1:0] node1183;
	wire [40-1:0] node1184;
	wire [40-1:0] node1185;
	wire [40-1:0] node1186;
	wire [40-1:0] node1187;
	wire [40-1:0] node1190;
	wire [40-1:0] node1193;
	wire [40-1:0] node1194;
	wire [40-1:0] node1197;
	wire [40-1:0] node1200;
	wire [40-1:0] node1201;
	wire [40-1:0] node1202;
	wire [40-1:0] node1205;
	wire [40-1:0] node1208;
	wire [40-1:0] node1209;
	wire [40-1:0] node1212;
	wire [40-1:0] node1215;
	wire [40-1:0] node1216;
	wire [40-1:0] node1217;
	wire [40-1:0] node1218;
	wire [40-1:0] node1221;
	wire [40-1:0] node1224;
	wire [40-1:0] node1225;
	wire [40-1:0] node1228;
	wire [40-1:0] node1231;
	wire [40-1:0] node1232;
	wire [40-1:0] node1233;
	wire [40-1:0] node1236;
	wire [40-1:0] node1239;
	wire [40-1:0] node1240;
	wire [40-1:0] node1243;

	assign outp = (inp[9]) ? node260 : node1;
		assign node1 = (inp[1]) ? node15 : node2;
			assign node2 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node3;
				assign node3 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node4;
					assign node4 = (inp[4]) ? node6 : 40'b0000000000000000000000000000000000000000;
						assign node6 = (inp[8]) ? node8 : 40'b0000000000000000000000000000000000000000;
							assign node8 = (inp[7]) ? node10 : 40'b0000000000000000000000000000000000000000;
								assign node10 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
			assign node15 = (inp[4]) ? node17 : 40'b0000000001000000000000000000000000000000;
				assign node17 = (inp[7]) ? node153 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[11]) ? node24 : node21;
								assign node21 = (inp[3]) ? 40'b0000000000100010000000000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[3]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000000010000001000000000000000000;
							assign node27 = (inp[11]) ? node31 : node28;
								assign node28 = (inp[3]) ? 40'b0000000000100000000000000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[3]) ? node33 : 40'b0000000000000000000001000000000010000000;
									assign node33 = (inp[13]) ? node39 : node34;
										assign node34 = (inp[0]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[10]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[10]) ? node43 : node40;
											assign node40 = (inp[0]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000010000000;
						assign node46 = (inp[14]) ? node104 : node47;
							assign node47 = (inp[0]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[3]) ? node67 : node50;
									assign node50 = (inp[15]) ? node52 : 40'b0000000000000000000000000000000000000000;
										assign node52 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node53;
											assign node53 = (inp[12]) ? node55 : 40'b0000000000000000000000000000000000000000;
												assign node55 = (inp[13]) ? node61 : node56;
													assign node56 = (inp[6]) ? node58 : 40'b0000000000000000000000000000000000000000;
														assign node58 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node61 = (inp[2]) ? node63 : 40'b0000000000000000000000000000000000000000;
														assign node63 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000100000000000000010;
									assign node67 = (inp[10]) ? node85 : node68;
										assign node68 = (inp[15]) ? node70 : 40'b0000000000000000000000000000000000000000;
											assign node70 = (inp[12]) ? node72 : 40'b0000000000000000000000000000000000000000;
												assign node72 = (inp[13]) ? node80 : node73;
													assign node73 = (inp[2]) ? node77 : node74;
														assign node74 = (inp[5]) ? 40'b0000000010000001010000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node77 = (inp[6]) ? 40'b0000000000000001010000000000000000000010 : 40'b0000000000000001010000000000001000000000;
													assign node80 = (inp[5]) ? node82 : 40'b0000000000000000000000000000000000000000;
														assign node82 = (inp[11]) ? 40'b0000000000000010010000100000010000000000 : 40'b0000000000000000000000000000000000000000;
										assign node85 = (inp[11]) ? node95 : node86;
											assign node86 = (inp[13]) ? 40'b0000000000000000000000000000001000000000 : node87;
												assign node87 = (inp[12]) ? node89 : 40'b0000000000000000000000000000000000000000;
													assign node89 = (inp[6]) ? 40'b0000000010000000010000100000000010000000 : node90;
														assign node90 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node95 = (inp[15]) ? node97 : 40'b0000000000000000000000000000000000000000;
												assign node97 = (inp[12]) ? node99 : 40'b0000000000000000000000000000000000000000;
													assign node99 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node100;
														assign node100 = (inp[2]) ? 40'b0000000000000000010000100000011010000000 : 40'b0000000000000000000000000000000000000000;
							assign node104 = (inp[3]) ? node108 : node105;
								assign node105 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node108 = (inp[0]) ? node122 : node109;
									assign node109 = (inp[2]) ? node111 : 40'b0000000000000000000000000000000000000000;
										assign node111 = (inp[6]) ? node113 : 40'b0000000000000000000000000000000000000000;
											assign node113 = (inp[15]) ? node115 : 40'b0000000000000000000000000000000000000000;
												assign node115 = (inp[12]) ? node117 : 40'b0000000000000000000000000000000000000000;
													assign node117 = (inp[5]) ? node119 : 40'b0000000000000000000000000000000000000000;
														assign node119 = (inp[11]) ? 40'b0000000000001000000000000000000001000000 : 40'b0000000000000000000100000000000001000000;
									assign node122 = (inp[13]) ? node140 : node123;
										assign node123 = (inp[12]) ? node125 : 40'b0000000000000000000000000000000000000000;
											assign node125 = (inp[15]) ? node127 : 40'b0000000000000000000000000000000000000000;
												assign node127 = (inp[5]) ? node133 : node128;
													assign node128 = (inp[2]) ? node130 : 40'b0000000000000000000000000000000000000000;
														assign node130 = (inp[6]) ? 40'b0000000000000000010000100000000011000010 : 40'b0000000000000000000000000000000000000000;
													assign node133 = (inp[10]) ? node137 : node134;
														assign node134 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000001001000000;
														assign node137 = (inp[6]) ? 40'b0000000010000000010100100000000011000000 : 40'b0000000000000000010100100000001011000000;
										assign node140 = (inp[10]) ? node150 : node141;
											assign node141 = (inp[12]) ? node143 : 40'b0000000000000000000000000000000000000000;
												assign node143 = (inp[5]) ? node145 : 40'b0000000000000000000000000000000000000000;
													assign node145 = (inp[15]) ? node147 : 40'b0000000000000000000000000000000000000000;
														assign node147 = (inp[6]) ? 40'b0000000010001010010000100000000001000000 : 40'b0000000000000000000000000000000000000000;
											assign node150 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node153 = (inp[14]) ? node187 : node154;
						assign node154 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node155;
							assign node155 = (inp[8]) ? node157 : 40'b0000000000000000000000000000000000000000;
								assign node157 = (inp[0]) ? node159 : 40'b0000000000000000000000000000000000000000;
									assign node159 = (inp[10]) ? node173 : node160;
										assign node160 = (inp[12]) ? node162 : 40'b0000000000000000000000000000000000000000;
											assign node162 = (inp[15]) ? node164 : 40'b0000000000000000000000000000000000000000;
												assign node164 = (inp[13]) ? node166 : 40'b0000000000000000000000000000000000000000;
													assign node166 = (inp[5]) ? node170 : node167;
														assign node167 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node170 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node173 = (inp[13]) ? node183 : node174;
											assign node174 = (inp[12]) ? node176 : 40'b0000000000000000000000000000000000000000;
												assign node176 = (inp[6]) ? node178 : 40'b0000000000000000000000000000000000000000;
													assign node178 = (inp[2]) ? 40'b0000000000000000000000100000000110000010 : node179;
														assign node179 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node183 = (inp[3]) ? 40'b0000000000000000000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
						assign node187 = (inp[8]) ? node205 : node188;
							assign node188 = (inp[11]) ? node190 : 40'b0000000000000000000000000000000000000000;
								assign node190 = (inp[3]) ? node192 : 40'b0000000000000000000000000000000000000000;
									assign node192 = (inp[13]) ? node198 : node193;
										assign node193 = (inp[10]) ? node195 : 40'b0000000000000000000000000000000000000000;
											assign node195 = (inp[0]) ? 40'b0000000000000000000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
										assign node198 = (inp[10]) ? node202 : node199;
											assign node199 = (inp[0]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
											assign node202 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000110000000;
							assign node205 = (inp[3]) ? node209 : node206;
								assign node206 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node209 = (inp[0]) ? node227 : node210;
									assign node210 = (inp[6]) ? node212 : 40'b0000000000000000000000000000000000000000;
										assign node212 = (inp[12]) ? node214 : 40'b0000000000000000000000000000000000000000;
											assign node214 = (inp[13]) ? node216 : 40'b0000000000000000000000000000000000000000;
												assign node216 = (inp[11]) ? node222 : node217;
													assign node217 = (inp[2]) ? node219 : 40'b0000000000000000000000000000000000000000;
														assign node219 = (inp[10]) ? 40'b0100000000000000000000001000010000000000 : 40'b0100000000000000000000001000000000000000;
													assign node222 = (inp[2]) ? node224 : 40'b0000000000000000000000000000000000000000;
														assign node224 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node227 = (inp[13]) ? node245 : node228;
										assign node228 = (inp[12]) ? node230 : 40'b0000000000000000000000000000000000000000;
											assign node230 = (inp[15]) ? node232 : 40'b0000000000000000000000000000000000000000;
												assign node232 = (inp[2]) ? node238 : node233;
													assign node233 = (inp[5]) ? node235 : 40'b0000000000000000000000000000000000000000;
														assign node235 = (inp[11]) ? 40'b0100000010000000000000000000000100000001 : 40'b0000000000000000000000000000000000000000;
													assign node238 = (inp[10]) ? node242 : node239;
														assign node239 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000000000001000000001000000100000000;
														assign node242 = (inp[6]) ? 40'b0100000000000000000000101000000110000010 : 40'b0100000000000000000000101000001110000000;
										assign node245 = (inp[10]) ? node257 : node246;
											assign node246 = (inp[15]) ? node248 : 40'b0000000000000000000000000000000000000000;
												assign node248 = (inp[12]) ? node250 : 40'b0000000000000000000000000000000000000000;
													assign node250 = (inp[5]) ? node254 : node251;
														assign node251 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node254 = (inp[2]) ? 40'b0100000000000010000000100000001100000000 : 40'b0100000010000010000000100000000100000000;
											assign node257 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node260 = (inp[1]) ? node328 : node261;
			assign node261 = (inp[8]) ? node265 : node262;
				assign node262 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node265 = (inp[7]) ? node297 : node266;
					assign node266 = (inp[3]) ? node282 : node267;
						assign node267 = (inp[11]) ? node275 : node268;
							assign node268 = (inp[14]) ? node272 : node269;
								assign node269 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node272 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
							assign node275 = (inp[14]) ? node279 : node276;
								assign node276 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node279 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
						assign node282 = (inp[14]) ? node290 : node283;
							assign node283 = (inp[11]) ? node287 : node284;
								assign node284 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node287 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
							assign node290 = (inp[11]) ? node294 : node291;
								assign node291 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
								assign node294 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node297 = (inp[11]) ? node313 : node298;
						assign node298 = (inp[3]) ? node306 : node299;
							assign node299 = (inp[14]) ? node303 : node300;
								assign node300 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node303 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
							assign node306 = (inp[14]) ? node310 : node307;
								assign node307 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node310 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
						assign node313 = (inp[3]) ? node321 : node314;
							assign node314 = (inp[14]) ? node318 : node315;
								assign node315 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
								assign node318 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
							assign node321 = (inp[14]) ? node325 : node322;
								assign node322 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
								assign node325 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node328 = (inp[8]) ? node332 : node329;
				assign node329 = (inp[4]) ? 40'b0000100000000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node332 = (inp[4]) ? node334 : 40'b0000000001000000000000000000000000000000;
					assign node334 = (inp[7]) ? node916 : node335;
						assign node335 = (inp[3]) ? node725 : node336;
							assign node336 = (inp[14]) ? node584 : node337;
								assign node337 = (inp[11]) ? node463 : node338;
									assign node338 = (inp[0]) ? node400 : node339;
										assign node339 = (inp[15]) ? node369 : node340;
											assign node340 = (inp[10]) ? node356 : node341;
												assign node341 = (inp[13]) ? node349 : node342;
													assign node342 = (inp[2]) ? node346 : node343;
														assign node343 = (inp[5]) ? 40'b1001000000010101010010000001101000010000 : 40'b1001000000010101010010000000101000010000;
														assign node346 = (inp[12]) ? 40'b0001000000010101010010000001101000010000 : 40'b0001000000010101010110000010101000010000;
													assign node349 = (inp[12]) ? node353 : node350;
														assign node350 = (inp[2]) ? 40'b0001000000010101010110000010001000010000 : 40'b1001000000010101010010000000001000010000;
														assign node353 = (inp[2]) ? 40'b0001000000010101010010000001001000010000 : 40'b0001000000011101010010000010001000010000;
												assign node356 = (inp[5]) ? node364 : node357;
													assign node357 = (inp[2]) ? node361 : node358;
														assign node358 = (inp[13]) ? 40'b1001000000011001010010000010001000010000 : 40'b1001000000011001010010000010101000010000;
														assign node361 = (inp[12]) ? 40'b1001000000010001010010000001001000010000 : 40'b1001000000010001010110000010001000010000;
													assign node364 = (inp[6]) ? node366 : 40'b0001000000010001010110000010101000010000;
														assign node366 = (inp[2]) ? 40'b0001000000010001010010000001101000010000 : 40'b1001000000010001010010000001001000010000;
											assign node369 = (inp[10]) ? node385 : node370;
												assign node370 = (inp[5]) ? node378 : node371;
													assign node371 = (inp[13]) ? node375 : node372;
														assign node372 = (inp[6]) ? 40'b0001000000001101010010000010101000010000 : 40'b1001000000000101010110000010101000010000;
														assign node375 = (inp[2]) ? 40'b0001000000000101010110000010001000010000 : 40'b1001000000001101010010000010001000010000;
													assign node378 = (inp[6]) ? node382 : node379;
														assign node379 = (inp[13]) ? 40'b0001000000000101010110000010001000010000 : 40'b0001000000000101010110000011101000010000;
														assign node382 = (inp[2]) ? 40'b0001000000000101010010000001001000010000 : 40'b1001000000000101010010000001001000010000;
												assign node385 = (inp[2]) ? node393 : node386;
													assign node386 = (inp[5]) ? node390 : node387;
														assign node387 = (inp[6]) ? 40'b0001000000001001010010000010101000010000 : 40'b1001000000000001010010000000101000010000;
														assign node390 = (inp[6]) ? 40'b1001000000000001010010000001001000010000 : 40'b1001000000000001010110000010001000010000;
													assign node393 = (inp[12]) ? node397 : node394;
														assign node394 = (inp[13]) ? 40'b0001000000001001010110000010001000010000 : 40'b0001000000000001010110000010101000010000;
														assign node397 = (inp[6]) ? 40'b0001000000001001010010000011001000010000 : 40'b0001000000000001010010000001101000010000;
										assign node400 = (inp[13]) ? node432 : node401;
											assign node401 = (inp[15]) ? node417 : node402;
												assign node402 = (inp[5]) ? node410 : node403;
													assign node403 = (inp[6]) ? node407 : node404;
														assign node404 = (inp[10]) ? 40'b1000000000010001010010000000101000010000 : 40'b1000000000010101010010000000101000010000;
														assign node407 = (inp[2]) ? 40'b0000000000011101010010000010101000010000 : 40'b1000000000011101010010000010101000010000;
													assign node410 = (inp[10]) ? node414 : node411;
														assign node411 = (inp[2]) ? 40'b0000000000010101010110000011101000010000 : 40'b1000000000010101010110000010101000010000;
														assign node414 = (inp[12]) ? 40'b0000000000010001010110000011101000010000 : 40'b0000000000010001010110000010101000010000;
												assign node417 = (inp[10]) ? node425 : node418;
													assign node418 = (inp[2]) ? node422 : node419;
														assign node419 = (inp[12]) ? 40'b0000000000001101010010000010101000010000 : 40'b1000000000000101010010000001101000010000;
														assign node422 = (inp[5]) ? 40'b0000000000000101010110000010101000010000 : 40'b1000000000000101010010000000101000010000;
													assign node425 = (inp[6]) ? node429 : node426;
														assign node426 = (inp[5]) ? 40'b0000000000000001010110000010101000010000 : 40'b1000000000000001010010000000101000010000;
														assign node429 = (inp[12]) ? 40'b0000000000001001010010000011101000010000 : 40'b0000000000000001010110000010101000010000;
											assign node432 = (inp[10]) ? node448 : node433;
												assign node433 = (inp[15]) ? node441 : node434;
													assign node434 = (inp[12]) ? node438 : node435;
														assign node435 = (inp[2]) ? 40'b0000000000010101010110000010001000010000 : 40'b1000000000010101010010000000001000010000;
														assign node438 = (inp[2]) ? 40'b0000000000010101010010000011001000010000 : 40'b0000000000011101010110000010001000010000;
													assign node441 = (inp[12]) ? node445 : node442;
														assign node442 = (inp[5]) ? 40'b1000000000000101010010000001001000010000 : 40'b0000000000000101010110000010001000010000;
														assign node445 = (inp[6]) ? 40'b0000000000001101010010000010001000010000 : 40'b0000000000001101010110000010001000010000;
												assign node448 = (inp[15]) ? node456 : node449;
													assign node449 = (inp[6]) ? node453 : node450;
														assign node450 = (inp[12]) ? 40'b0000000000010001010110000010001000010000 : 40'b1000000000010001010110000010001000010000;
														assign node453 = (inp[5]) ? 40'b0000000000010001010010000001001000010000 : 40'b0000000000011001010010000010001000010000;
													assign node456 = (inp[5]) ? node460 : node457;
														assign node457 = (inp[12]) ? 40'b1000000000000001010010000001001000010000 : 40'b1000000000000001010010000000001000010000;
														assign node460 = (inp[2]) ? 40'b0000000000000001010110000011001000010000 : 40'b0000000000001001010010000010001000010000;
									assign node463 = (inp[10]) ? node525 : node464;
										assign node464 = (inp[0]) ? node494 : node465;
											assign node465 = (inp[15]) ? node479 : node466;
												assign node466 = (inp[2]) ? node472 : node467;
													assign node467 = (inp[13]) ? 40'b1001000000011101010010000010001000000000 : node468;
														assign node468 = (inp[12]) ? 40'b0001000000011101010010000010101000000000 : 40'b1001000000010101010110000010101000000000;
													assign node472 = (inp[6]) ? node476 : node473;
														assign node473 = (inp[5]) ? 40'b0001000000010101010110000010101000000000 : 40'b1001000000010101010010000001101000000000;
														assign node476 = (inp[5]) ? 40'b0001000000010101010010000001001000000000 : 40'b0001000000011101010010000011001000000000;
												assign node479 = (inp[13]) ? node487 : node480;
													assign node480 = (inp[12]) ? node484 : node481;
														assign node481 = (inp[2]) ? 40'b0001000000001101010110000010101000000000 : 40'b1001000000000101010010000000101000000000;
														assign node484 = (inp[2]) ? 40'b0001000000000101010010000001101000000000 : 40'b0001000000001101010010000010101000000000;
													assign node487 = (inp[5]) ? node491 : node488;
														assign node488 = (inp[6]) ? 40'b0001000000001101010010000010001000000000 : 40'b1001000000000101010010000010001000000000;
														assign node491 = (inp[2]) ? 40'b0001000000000101010110000011001000000000 : 40'b1001000000000101010010000001001000000000;
											assign node494 = (inp[15]) ? node510 : node495;
												assign node495 = (inp[13]) ? node503 : node496;
													assign node496 = (inp[2]) ? node500 : node497;
														assign node497 = (inp[12]) ? 40'b0000000000011101010010000010101000000000 : 40'b1000000000010101010010000000101000000000;
														assign node500 = (inp[5]) ? 40'b0000000000010101010110000011101000000000 : 40'b0000000000010101010110000010101000000000;
													assign node503 = (inp[5]) ? node507 : node504;
														assign node504 = (inp[2]) ? 40'b1000000000010101010010000001001000000000 : 40'b1000000000011101010010000010001000000000;
														assign node507 = (inp[6]) ? 40'b0000000000010101010010000001001000000000 : 40'b0000000000010101010110000010001000000000;
												assign node510 = (inp[2]) ? node518 : node511;
													assign node511 = (inp[13]) ? node515 : node512;
														assign node512 = (inp[12]) ? 40'b0000000000001101010010000010101000000000 : 40'b1000000000001101010010000010101000000000;
														assign node515 = (inp[12]) ? 40'b0000000000001101010010000010001000000000 : 40'b1000000000000101010010000000001000000000;
													assign node518 = (inp[13]) ? node522 : node519;
														assign node519 = (inp[6]) ? 40'b0000000000000101010010000011101000000000 : 40'b0000000000000101010110000010101000000000;
														assign node522 = (inp[5]) ? 40'b0000000000000101010110000011001000000000 : 40'b0000000000001101010010000011001000000000;
										assign node525 = (inp[13]) ? node557 : node526;
											assign node526 = (inp[0]) ? node542 : node527;
												assign node527 = (inp[15]) ? node535 : node528;
													assign node528 = (inp[12]) ? node532 : node529;
														assign node529 = (inp[6]) ? 40'b0001000000011001010110000010101000000000 : 40'b0001000000010001010110000010101000000000;
														assign node532 = (inp[2]) ? 40'b0001000000010001010010000001101000000000 : 40'b0001000000011001010010000010101000000000;
													assign node535 = (inp[6]) ? node539 : node536;
														assign node536 = (inp[12]) ? 40'b0001000000001001010110000010101000000000 : 40'b0001000000000001010110000010101000000000;
														assign node539 = (inp[12]) ? 40'b0001000000000001010010000001101000000000 : 40'b0001000000001001010010000010101000000000;
												assign node542 = (inp[15]) ? node550 : node543;
													assign node543 = (inp[5]) ? node547 : node544;
														assign node544 = (inp[6]) ? 40'b0000000000011001010010000010101000000000 : 40'b1000000000010001010010000001101000000000;
														assign node547 = (inp[2]) ? 40'b0000000000010001010110000011101000000000 : 40'b0000000000010001010110000010101000000000;
													assign node550 = (inp[6]) ? node554 : node551;
														assign node551 = (inp[12]) ? 40'b0000000000000001010110000011101000000000 : 40'b1000000000000001010110000010101000000000;
														assign node554 = (inp[5]) ? 40'b0000000000000001010010000001101000000000 : 40'b0000000000001001010010000010101000000000;
											assign node557 = (inp[0]) ? node569 : node558;
												assign node558 = (inp[5]) ? node564 : node559;
													assign node559 = (inp[6]) ? node561 : 40'b1001000000000001010110000010001000000000;
														assign node561 = (inp[15]) ? 40'b0001000000001001010010000010001000000000 : 40'b0001000000011001010010000010001000000000;
													assign node564 = (inp[6]) ? node566 : 40'b0001000000001001010110000010001000000000;
														assign node566 = (inp[2]) ? 40'b0001000000000001010110000011001000000000 : 40'b1001000000010001010010000001001000000000;
												assign node569 = (inp[15]) ? node577 : node570;
													assign node570 = (inp[2]) ? node574 : node571;
														assign node571 = (inp[12]) ? 40'b0000000000011001010010000010001000000000 : 40'b1000000000010001010010000010001000000000;
														assign node574 = (inp[12]) ? 40'b0000000000010001010010000001001000000000 : 40'b0000000000010001010110000010001000000000;
													assign node577 = (inp[6]) ? node581 : node578;
														assign node578 = (inp[5]) ? 40'b0000000000000001010110000010001000000000 : 40'b1000000000000001010010000000001000000000;
														assign node581 = (inp[5]) ? 40'b0000000000000001010010000001001000000000 : 40'b0000000000001001010010000010001000000000;
								assign node584 = (inp[11]) ? node600 : node585;
									assign node585 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node586;
										assign node586 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node587;
											assign node587 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node588;
												assign node588 = (inp[10]) ? node594 : node589;
													assign node589 = (inp[2]) ? node591 : 40'b0000000000000000000000000000000000000000;
														assign node591 = (inp[0]) ? 40'b0000000000000100001100000010000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node594 = (inp[13]) ? 40'b1001000000010000001000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node600 = (inp[0]) ? node664 : node601;
										assign node601 = (inp[10]) ? node633 : node602;
											assign node602 = (inp[13]) ? node618 : node603;
												assign node603 = (inp[15]) ? node611 : node604;
													assign node604 = (inp[6]) ? node608 : node605;
														assign node605 = (inp[12]) ? 40'b1001010000010100000000000001100000000000 : 40'b1001010000010100000000000000100000000000;
														assign node608 = (inp[5]) ? 40'b0001010000010100000000000001100000000000 : 40'b0001010000011100000000000011100000000000;
													assign node611 = (inp[12]) ? node615 : node612;
														assign node612 = (inp[2]) ? 40'b0001010000000100000100000010100000000000 : 40'b1001010000000100000000000010100000000000;
														assign node615 = (inp[2]) ? 40'b0001010000000100000000000001100000000000 : 40'b0001010000001100000000000010100000000000;
												assign node618 = (inp[12]) ? node626 : node619;
													assign node619 = (inp[15]) ? node623 : node620;
														assign node620 = (inp[6]) ? 40'b1001010000010100000000000000000000000000 : 40'b1001010000010100000100000010000000000000;
														assign node623 = (inp[2]) ? 40'b0001010000000100000100000011000000000000 : 40'b1001010000000100000000000000000000000000;
													assign node626 = (inp[15]) ? node630 : node627;
														assign node627 = (inp[6]) ? 40'b0001010000011100000000000011000000000000 : 40'b0001010000010100000100000010000000000000;
														assign node630 = (inp[6]) ? 40'b0001010000001100000000000011000000000000 : 40'b0001010000000100000100000011000000000000;
											assign node633 = (inp[15]) ? node649 : node634;
												assign node634 = (inp[13]) ? node642 : node635;
													assign node635 = (inp[5]) ? node639 : node636;
														assign node636 = (inp[12]) ? 40'b0001010000011000000000000010100000000000 : 40'b0001010000011000000000000010100000000000;
														assign node639 = (inp[12]) ? 40'b0001010000011000000100000010100000000000 : 40'b0001010000010000000100000010100000000000;
													assign node642 = (inp[2]) ? node646 : node643;
														assign node643 = (inp[5]) ? 40'b1001010000010000000100000010000000000000 : 40'b1001010000011000000000000010000000000000;
														assign node646 = (inp[12]) ? 40'b0001010000010000000000000011000000000000 : 40'b0001010000010000000100000010000000000000;
												assign node649 = (inp[13]) ? node657 : node650;
													assign node650 = (inp[2]) ? node654 : node651;
														assign node651 = (inp[12]) ? 40'b0001010000001000000000000010100000000000 : 40'b1001010000000000000000000000100000000000;
														assign node654 = (inp[12]) ? 40'b0001010000000000000000000011100000000000 : 40'b0001010000000000000100000010100000000000;
													assign node657 = (inp[5]) ? node661 : node658;
														assign node658 = (inp[6]) ? 40'b0001010000001000000000000010000000000000 : 40'b1001010000000000000000000000000000000000;
														assign node661 = (inp[2]) ? 40'b0001010000000000000100000010000000000000 : 40'b0001010000001000000100000010000000000000;
										assign node664 = (inp[13]) ? node696 : node665;
											assign node665 = (inp[15]) ? node681 : node666;
												assign node666 = (inp[10]) ? node674 : node667;
													assign node667 = (inp[5]) ? node671 : node668;
														assign node668 = (inp[6]) ? 40'b0000010000011100000000000010100000000000 : 40'b1000010000010100000000000000100000000000;
														assign node671 = (inp[6]) ? 40'b0000010000010100000000000001100000000000 : 40'b0000010000010100000100000010100000000000;
													assign node674 = (inp[2]) ? node678 : node675;
														assign node675 = (inp[5]) ? 40'b1000010000010000000000000001100000000000 : 40'b1000010000010000000000000000100000000000;
														assign node678 = (inp[6]) ? 40'b0000010000010000000000000011100000000000 : 40'b1000010000010000000000000001100000000000;
												assign node681 = (inp[10]) ? node689 : node682;
													assign node682 = (inp[2]) ? node686 : node683;
														assign node683 = (inp[12]) ? 40'b0000010000001100000000000010100000000000 : 40'b1000010000000100000000000000100000000000;
														assign node686 = (inp[12]) ? 40'b0000010000000100000000000011100000000000 : 40'b0000010000001100000100000010100000000000;
													assign node689 = (inp[2]) ? node693 : node690;
														assign node690 = (inp[12]) ? 40'b0000010000001000000000000010100000000000 : 40'b1000010000000000000000000000100000000000;
														assign node693 = (inp[12]) ? 40'b0000010000000000000000000001100000000000 : 40'b0000010000000000000100000010100000000000;
											assign node696 = (inp[10]) ? node712 : node697;
												assign node697 = (inp[5]) ? node705 : node698;
													assign node698 = (inp[12]) ? node702 : node699;
														assign node699 = (inp[6]) ? 40'b1000010000001100000000000010000000000000 : 40'b1000010000010100000000000000000000000000;
														assign node702 = (inp[15]) ? 40'b0000010000001100000000000010000000000000 : 40'b0000010000011100000000000010000000000000;
													assign node705 = (inp[2]) ? node709 : node706;
														assign node706 = (inp[15]) ? 40'b1000010000000100000000000001000000000000 : 40'b1000010000010100000000000001000000000000;
														assign node709 = (inp[12]) ? 40'b0000010000000100000000000001000000000000 : 40'b0000010000010100000100000011000000000000;
												assign node712 = (inp[12]) ? node720 : node713;
													assign node713 = (inp[15]) ? node717 : node714;
														assign node714 = (inp[6]) ? 40'b0000010000011000000100000010000000000000 : 40'b1000010000010000000100000010000000000000;
														assign node717 = (inp[5]) ? 40'b0000010000000000000100000010000000000000 : 40'b0000010000001000000100000010000000000000;
													assign node720 = (inp[6]) ? node722 : 40'b1000010000011000000000000010000000000000;
														assign node722 = (inp[15]) ? 40'b0000010000001000000000000011000000000000 : 40'b0000010000011000000000000011000000000000;
							assign node725 = (inp[14]) ? node791 : node726;
								assign node726 = (inp[11]) ? node776 : node727;
									assign node727 = (inp[12]) ? node765 : node728;
										assign node728 = (inp[6]) ? node748 : node729;
											assign node729 = (inp[13]) ? node739 : node730;
												assign node730 = (inp[15]) ? node732 : 40'b0000000000000000000000000000000000000000;
													assign node732 = (inp[2]) ? node736 : node733;
														assign node733 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node736 = (inp[10]) ? 40'b0001000000000000000100000010100000100000 : 40'b0000000000000100000100000010100000100000;
												assign node739 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node740;
													assign node740 = (inp[5]) ? node744 : node741;
														assign node741 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b1001000000010000000000000000000000100000;
														assign node744 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node748 = (inp[0]) ? node758 : node749;
												assign node749 = (inp[10]) ? node751 : 40'b0000000000000000000000000000000000000000;
													assign node751 = (inp[13]) ? node755 : node752;
														assign node752 = (inp[2]) ? 40'b0001000000000000000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
														assign node755 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node758 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node759;
													assign node759 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node760;
														assign node760 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000011100000000000010000000100000;
										assign node765 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node766;
											assign node766 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node767;
												assign node767 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node768;
													assign node768 = (inp[5]) ? node770 : 40'b0000000000000000000000000000000000000000;
														assign node770 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0001000000001000000100000010100000100000;
									assign node776 = (inp[2]) ? node778 : 40'b0000000000000000000000000000000000000000;
										assign node778 = (inp[12]) ? node780 : 40'b0000000000000000000000000000000000000000;
											assign node780 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node781;
												assign node781 = (inp[5]) ? node783 : 40'b0000000000000000000000000000000000000000;
													assign node783 = (inp[15]) ? node787 : node784;
														assign node784 = (inp[0]) ? 40'b1000000000010100001000000000100000010000 : 40'b0000000000000000000000000000000000000000;
														assign node787 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
								assign node791 = (inp[11]) ? node793 : 40'b0000000000000000000000000000000000000000;
									assign node793 = (inp[15]) ? node853 : node794;
										assign node794 = (inp[13]) ? node822 : node795;
											assign node795 = (inp[10]) ? node807 : node796;
												assign node796 = (inp[6]) ? node802 : node797;
													assign node797 = (inp[0]) ? node799 : 40'b1011000000010100000000000001100000000000;
														assign node799 = (inp[2]) ? 40'b0010000000010100000100000010100000000000 : 40'b0010000000011100000000000010100000000000;
													assign node802 = (inp[12]) ? node804 : 40'b1010000000010100000000000001100000000000;
														assign node804 = (inp[2]) ? 40'b0010000000010100000000000001100000000000 : 40'b0010000000011100000000000011100000000000;
												assign node807 = (inp[5]) ? node815 : node808;
													assign node808 = (inp[2]) ? node812 : node809;
														assign node809 = (inp[0]) ? 40'b1010000000011000000000000010100000000000 : 40'b1011000000011000000000000010100000000000;
														assign node812 = (inp[12]) ? 40'b1010000000010000000000000001100000000000 : 40'b0010000000010000000100000010100000000000;
													assign node815 = (inp[0]) ? node819 : node816;
														assign node816 = (inp[2]) ? 40'b0011000000010000000100000011100000000000 : 40'b0011000000011000000000000011100000000000;
														assign node819 = (inp[2]) ? 40'b0010000000010000000100000011100000000000 : 40'b1010000000010000000000000001100000000000;
											assign node822 = (inp[0]) ? node838 : node823;
												assign node823 = (inp[10]) ? node831 : node824;
													assign node824 = (inp[6]) ? node828 : node825;
														assign node825 = (inp[12]) ? 40'b0011000000011100000100000010000000000000 : 40'b1011000000010100000100000010000000000000;
														assign node828 = (inp[5]) ? 40'b1011000000010100000000000001000000000000 : 40'b0011000000011100000000000010000000000000;
													assign node831 = (inp[5]) ? node835 : node832;
														assign node832 = (inp[6]) ? 40'b0011000000011000000000000010000000000000 : 40'b1011000000010000000000000001000000000000;
														assign node835 = (inp[2]) ? 40'b0011000000010000000100000011000000000000 : 40'b0011000000010000000100000010000000000000;
												assign node838 = (inp[12]) ? node846 : node839;
													assign node839 = (inp[10]) ? node843 : node840;
														assign node840 = (inp[2]) ? 40'b0010000000010100000100000010000000000000 : 40'b1010000000010100000000000010000000000000;
														assign node843 = (inp[2]) ? 40'b0010000000010000000100000010000000000000 : 40'b1010000000010000000100000010000000000000;
													assign node846 = (inp[10]) ? node850 : node847;
														assign node847 = (inp[6]) ? 40'b0010000000011100000000000011000000000000 : 40'b0010000000011100000100000010000000000000;
														assign node850 = (inp[2]) ? 40'b0010000000010000000000000001000000000000 : 40'b0010000000011000000000000010000000000000;
										assign node853 = (inp[0]) ? node885 : node854;
											assign node854 = (inp[13]) ? node870 : node855;
												assign node855 = (inp[2]) ? node863 : node856;
													assign node856 = (inp[12]) ? node860 : node857;
														assign node857 = (inp[10]) ? 40'b1011000000000000000000000000100000000000 : 40'b1011000000001100000000000010100000000000;
														assign node860 = (inp[6]) ? 40'b0011000000001000000000000010100000000000 : 40'b0011000000001000000100000010100000000000;
													assign node863 = (inp[10]) ? node867 : node864;
														assign node864 = (inp[5]) ? 40'b0011000000000100000000000001100000000000 : 40'b1011000000000100000000000001100000000000;
														assign node867 = (inp[5]) ? 40'b0011000000000000000100000011100000000000 : 40'b0011000000001000000000000011100000000000;
												assign node870 = (inp[10]) ? node878 : node871;
													assign node871 = (inp[6]) ? node875 : node872;
														assign node872 = (inp[5]) ? 40'b1011000000000100000100000010000000000000 : 40'b1011000000000100000000000000000000000000;
														assign node875 = (inp[12]) ? 40'b0011000000001100000000000011000000000000 : 40'b0011000000000100000100000010000000000000;
													assign node878 = (inp[6]) ? node882 : node879;
														assign node879 = (inp[12]) ? 40'b0011000000000000000100000011000000000000 : 40'b0011000000000000000100000010000000000000;
														assign node882 = (inp[2]) ? 40'b0011000000000000000000000001000000000000 : 40'b0011000000000000000000000001000000000000;
											assign node885 = (inp[10]) ? node901 : node886;
												assign node886 = (inp[13]) ? node894 : node887;
													assign node887 = (inp[6]) ? node891 : node888;
														assign node888 = (inp[5]) ? 40'b0010000000000100000100000010100000000000 : 40'b1010000000000100000000000000100000000000;
														assign node891 = (inp[5]) ? 40'b0010000000000100000000000001100000000000 : 40'b0010000000001100000000000010100000000000;
													assign node894 = (inp[2]) ? node898 : node895;
														assign node895 = (inp[6]) ? 40'b1010000000001100000000000010000000000000 : 40'b1010000000000100000000000000000000000000;
														assign node898 = (inp[12]) ? 40'b0010000000000100000000000001000000000000 : 40'b0010000000000100000100000010000000000000;
												assign node901 = (inp[13]) ? node909 : node902;
													assign node902 = (inp[12]) ? node906 : node903;
														assign node903 = (inp[5]) ? 40'b1010000000000000000000000001100000000000 : 40'b1010000000000000000000000000100000000000;
														assign node906 = (inp[6]) ? 40'b0010000000001000000000000011100000000000 : 40'b0010000000001000000000000010100000000000;
													assign node909 = (inp[12]) ? node913 : node910;
														assign node910 = (inp[2]) ? 40'b0010000000000000000100000010000000000000 : 40'b1010000000000000000000000000000000000000;
														assign node913 = (inp[2]) ? 40'b0010000000000000000000000001000000000000 : 40'b0010000000001000000000000010000000000000;
						assign node916 = (inp[3]) ? node988 : node917;
							assign node917 = (inp[14]) ? node943 : node918;
								assign node918 = (inp[11]) ? node920 : 40'b0000000000000000000000000000000000000000;
									assign node920 = (inp[15]) ? node932 : node921;
										assign node921 = (inp[0]) ? node927 : node922;
											assign node922 = (inp[10]) ? node924 : 40'b0000000000000000000000000000000000000000;
												assign node924 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
											assign node927 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node928;
												assign node928 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
										assign node932 = (inp[0]) ? node938 : node933;
											assign node933 = (inp[10]) ? node935 : 40'b0000000000000000000000000000000000000000;
												assign node935 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
											assign node938 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node939;
												assign node939 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
								assign node943 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node944;
									assign node944 = (inp[13]) ? node956 : node945;
										assign node945 = (inp[10]) ? node947 : 40'b0000000000000000000000000000000000000000;
											assign node947 = (inp[15]) ? node949 : 40'b0000000000000000000000000000000000000000;
												assign node949 = (inp[0]) ? node951 : 40'b0000000000000000000000000000000000000000;
													assign node951 = (inp[12]) ? node953 : 40'b1000001100000000000100000010100000000000;
														assign node953 = (inp[2]) ? 40'b0000001100000000000000000001100000000000 : 40'b0000001100001000000000000010100000000000;
										assign node956 = (inp[15]) ? node968 : node957;
											assign node957 = (inp[0]) ? node959 : 40'b0000000000000000000000000000000000000000;
												assign node959 = (inp[10]) ? node961 : 40'b0000000000000000000000000000000000000000;
													assign node961 = (inp[2]) ? node965 : node962;
														assign node962 = (inp[5]) ? 40'b1000001100010000000000000001000000000000 : 40'b1000001100011000000000000010000000000000;
														assign node965 = (inp[5]) ? 40'b0000001100010000000100000011000000000000 : 40'b1000001100010000000100000010000000000000;
											assign node968 = (inp[10]) ? node978 : node969;
												assign node969 = (inp[0]) ? node971 : 40'b0000000000000000000000000000000000000000;
													assign node971 = (inp[6]) ? node975 : node972;
														assign node972 = (inp[12]) ? 40'b0000001100000100000000000001000000000000 : 40'b0000001100000100000100000010000000000000;
														assign node975 = (inp[5]) ? 40'b0000001100000100000000000001000000000000 : 40'b0000001100001100000000000010000000000000;
												assign node978 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node979;
													assign node979 = (inp[12]) ? node983 : node980;
														assign node980 = (inp[2]) ? 40'b0001001100000000000100000010000000000000 : 40'b1001001100000000000000000000000000000000;
														assign node983 = (inp[6]) ? 40'b0001001100001000000000000011000000000000 : 40'b0001001100001000000000000010000000000000;
							assign node988 = (inp[11]) ? node1118 : node989;
								assign node989 = (inp[14]) ? node991 : 40'b0000000000000000000000000000000000000000;
									assign node991 = (inp[13]) ? node1055 : node992;
										assign node992 = (inp[10]) ? node1024 : node993;
											assign node993 = (inp[0]) ? node1009 : node994;
												assign node994 = (inp[2]) ? node1002 : node995;
													assign node995 = (inp[6]) ? node999 : node996;
														assign node996 = (inp[12]) ? 40'b1001001000001100000000000010100000000000 : 40'b1001001000010100000000000000100000000000;
														assign node999 = (inp[12]) ? 40'b0001001000011100000000000011100000000000 : 40'b1001001000001100000000000010100000000000;
													assign node1002 = (inp[5]) ? node1006 : node1003;
														assign node1003 = (inp[12]) ? 40'b0001001000011100000000000011100000000000 : 40'b0001001000001100000100000010100000000000;
														assign node1006 = (inp[15]) ? 40'b0001001000000100000100000011100000000000 : 40'b0001001000010100000100000011100000000000;
												assign node1009 = (inp[12]) ? node1017 : node1010;
													assign node1010 = (inp[2]) ? node1014 : node1011;
														assign node1011 = (inp[15]) ? 40'b1000001000000100000000000000100000000000 : 40'b1000001000010100000000000010100000000000;
														assign node1014 = (inp[15]) ? 40'b0000001000000100000100000010100000000000 : 40'b0000001000010100000100000010100000000000;
													assign node1017 = (inp[15]) ? node1021 : node1018;
														assign node1018 = (inp[6]) ? 40'b0000001000011100000000000011100000000000 : 40'b0000001000011100000000000010100000000000;
														assign node1021 = (inp[6]) ? 40'b0000001000001100000000000010100000000000 : 40'b0000001000001100000100000010100000000000;
											assign node1024 = (inp[15]) ? node1040 : node1025;
												assign node1025 = (inp[0]) ? node1033 : node1026;
													assign node1026 = (inp[6]) ? node1030 : node1027;
														assign node1027 = (inp[5]) ? 40'b0001001000010000000100000010100000000000 : 40'b1001001000010000000000000000100000000000;
														assign node1030 = (inp[5]) ? 40'b0001001000010000000000000001100000000000 : 40'b0001001000011000000000000010100000000000;
													assign node1033 = (inp[5]) ? node1037 : node1034;
														assign node1034 = (inp[6]) ? 40'b0000001000011000000100000010100000000000 : 40'b1000001000010000000100000010100000000000;
														assign node1037 = (inp[12]) ? 40'b0000001000010000000000000001100000000000 : 40'b0000001000010000000100000011100000000000;
												assign node1040 = (inp[5]) ? node1048 : node1041;
													assign node1041 = (inp[6]) ? node1045 : node1042;
														assign node1042 = (inp[0]) ? 40'b1000001000000000000000000000100000000000 : 40'b1001001000000000000000000000100000000000;
														assign node1045 = (inp[12]) ? 40'b0000001000001000000000000011100000000000 : 40'b1000001000001000000000000010100000000000;
													assign node1048 = (inp[2]) ? node1052 : node1049;
														assign node1049 = (inp[12]) ? 40'b0000001000001000000100000010100000000000 : 40'b1001001000000000000100000010100000000000;
														assign node1052 = (inp[0]) ? 40'b0000001000000000000100000011100000000000 : 40'b0001001000000000000100000011100000000000;
										assign node1055 = (inp[15]) ? node1087 : node1056;
											assign node1056 = (inp[0]) ? node1072 : node1057;
												assign node1057 = (inp[10]) ? node1065 : node1058;
													assign node1058 = (inp[5]) ? node1062 : node1059;
														assign node1059 = (inp[6]) ? 40'b0001001000011100000000000010000000000000 : 40'b1001001000010100000000000000000000000000;
														assign node1062 = (inp[6]) ? 40'b0001001000010100000000000001000000000000 : 40'b0001001000010100000100000011000000000000;
													assign node1065 = (inp[12]) ? node1069 : node1066;
														assign node1066 = (inp[2]) ? 40'b0001001000010000000100000010000000000000 : 40'b1001001000010000000000000000000000000000;
														assign node1069 = (inp[6]) ? 40'b0001001000011000000000000011000000000000 : 40'b0001001000011000000000000010000000000000;
												assign node1072 = (inp[10]) ? node1080 : node1073;
													assign node1073 = (inp[2]) ? node1077 : node1074;
														assign node1074 = (inp[12]) ? 40'b0000001000011100000100000010000000000000 : 40'b1000001000010100000000000000000000000000;
														assign node1077 = (inp[5]) ? 40'b0000001000010100000100000011000000000000 : 40'b0000001000011100000000000011000000000000;
													assign node1080 = (inp[5]) ? node1084 : node1081;
														assign node1081 = (inp[6]) ? 40'b0000001000011000000000000010000000000000 : 40'b1000001000010000000000000000000000000000;
														assign node1084 = (inp[2]) ? 40'b0000001000010000000100000011000000000000 : 40'b0000001000011000000000000011000000000000;
											assign node1087 = (inp[10]) ? node1103 : node1088;
												assign node1088 = (inp[0]) ? node1096 : node1089;
													assign node1089 = (inp[6]) ? node1093 : node1090;
														assign node1090 = (inp[12]) ? 40'b0001001000001100000000000010000000000000 : 40'b1001001000000100000100000010000000000000;
														assign node1093 = (inp[12]) ? 40'b0001001000001100000000000011000000000000 : 40'b0001001000000100000100000010000000000000;
													assign node1096 = (inp[2]) ? node1100 : node1097;
														assign node1097 = (inp[6]) ? 40'b0000001000001100000000000010000000000000 : 40'b0000001000001100000000000010000000000000;
														assign node1100 = (inp[12]) ? 40'b0000001000000100000000000001000000000000 : 40'b0000001000000100000100000010000000000000;
												assign node1103 = (inp[0]) ? node1111 : node1104;
													assign node1104 = (inp[5]) ? node1108 : node1105;
														assign node1105 = (inp[2]) ? 40'b0001001000000000000000000001000000000000 : 40'b1001001000001000000000000010000000000000;
														assign node1108 = (inp[2]) ? 40'b0001001000000000000000000001000000000000 : 40'b1001001000000000000000000001000000000000;
													assign node1111 = (inp[5]) ? node1115 : node1112;
														assign node1112 = (inp[6]) ? 40'b0000001000001000000000000010000000000000 : 40'b1000001000001000000000000010000000000000;
														assign node1115 = (inp[6]) ? 40'b0000001000000000000000000001000000000000 : 40'b0000001000000000000100000010000000000000;
								assign node1118 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node1119;
									assign node1119 = (inp[0]) ? node1183 : node1120;
										assign node1120 = (inp[15]) ? node1152 : node1121;
											assign node1121 = (inp[10]) ? node1137 : node1122;
												assign node1122 = (inp[13]) ? node1130 : node1123;
													assign node1123 = (inp[12]) ? node1127 : node1124;
														assign node1124 = (inp[6]) ? 40'b1001001000011100000000000010100000001000 : 40'b1001001000010100000100000010100000001000;
														assign node1127 = (inp[6]) ? 40'b0001001000011100000000000011100000001000 : 40'b0001001000010100000000000010100000001000;
													assign node1130 = (inp[5]) ? node1134 : node1131;
														assign node1131 = (inp[6]) ? 40'b0001001000011100000100000010000000001000 : 40'b1001001000010100000000000000000000001000;
														assign node1134 = (inp[6]) ? 40'b0001001000011100000000000011000000001000 : 40'b0001001000010100000100000010000000001000;
												assign node1137 = (inp[13]) ? node1145 : node1138;
													assign node1138 = (inp[2]) ? node1142 : node1139;
														assign node1139 = (inp[12]) ? 40'b0001001000011000000100000010100000001000 : 40'b1001001000010000000000000000100000001000;
														assign node1142 = (inp[5]) ? 40'b0001001000010000000100000010100000001000 : 40'b0001001000011000000100000010100000001000;
													assign node1145 = (inp[2]) ? node1149 : node1146;
														assign node1146 = (inp[5]) ? 40'b0001001000010000000100000010000000001000 : 40'b1001001000011000000000000010000000001000;
														assign node1149 = (inp[12]) ? 40'b0001001000010000000000000001000000001000 : 40'b0001001000010000000100000010000000001000;
											assign node1152 = (inp[6]) ? node1168 : node1153;
												assign node1153 = (inp[10]) ? node1161 : node1154;
													assign node1154 = (inp[13]) ? node1158 : node1155;
														assign node1155 = (inp[12]) ? 40'b1001001000000100000000000000100000001000 : 40'b1001001000000100000100000010100000001000;
														assign node1158 = (inp[12]) ? 40'b1001001000000100000000000001000000001000 : 40'b1001001000000100000100000010000000001000;
													assign node1161 = (inp[5]) ? node1165 : node1162;
														assign node1162 = (inp[13]) ? 40'b1001001000000000000000000000000000001000 : 40'b1001001000000000000100000010100000001000;
														assign node1165 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000001000000100000010100000001000;
												assign node1168 = (inp[13]) ? node1176 : node1169;
													assign node1169 = (inp[10]) ? node1173 : node1170;
														assign node1170 = (inp[2]) ? 40'b0001001000000100000000000001100000001000 : 40'b0001001000001100000000000011100000001000;
														assign node1173 = (inp[2]) ? 40'b0001001000000000000000000001100000001000 : 40'b0001001000000000000000000001100000001000;
													assign node1176 = (inp[10]) ? node1180 : node1177;
														assign node1177 = (inp[2]) ? 40'b0001001000000100000000000011000000001000 : 40'b1001001000000100000000000001000000001000;
														assign node1180 = (inp[12]) ? 40'b0001001000001000000000000011000000001000 : 40'b1001001000000000000000000001000000001000;
										assign node1183 = (inp[15]) ? node1215 : node1184;
											assign node1184 = (inp[10]) ? node1200 : node1185;
												assign node1185 = (inp[13]) ? node1193 : node1186;
													assign node1186 = (inp[5]) ? node1190 : node1187;
														assign node1187 = (inp[2]) ? 40'b0000001000010100000000000000100000001000 : 40'b1000001000011100000000000010100000001000;
														assign node1190 = (inp[12]) ? 40'b0000001000011100000000000011100000001000 : 40'b1000001000010100000000000001100000001000;
													assign node1193 = (inp[12]) ? node1197 : node1194;
														assign node1194 = (inp[6]) ? 40'b0000001000010100000000000001000000001000 : 40'b1000001000010100000100000010000000001000;
														assign node1197 = (inp[2]) ? 40'b0000001000010100000100000011000000001000 : 40'b0000001000011100000000000010000000001000;
												assign node1200 = (inp[13]) ? node1208 : node1201;
													assign node1201 = (inp[12]) ? node1205 : node1202;
														assign node1202 = (inp[6]) ? 40'b0000001000010000000100000010100000001000 : 40'b1000001000010000000100000010100000001000;
														assign node1205 = (inp[5]) ? 40'b0000001000010000000000000001100000001000 : 40'b1000001000010000000000000001100000001000;
													assign node1208 = (inp[2]) ? node1212 : node1209;
														assign node1209 = (inp[5]) ? 40'b1000001000010000000000000001000000001000 : 40'b1000001000011000000000000010000000001000;
														assign node1212 = (inp[12]) ? 40'b0000001000010000000000000011000000001000 : 40'b0000001000010000000100000010000000001000;
											assign node1215 = (inp[10]) ? node1231 : node1216;
												assign node1216 = (inp[13]) ? node1224 : node1217;
													assign node1217 = (inp[12]) ? node1221 : node1218;
														assign node1218 = (inp[2]) ? 40'b0000001000000100000100000010100000001000 : 40'b1000001000000100000000000000100000001000;
														assign node1221 = (inp[6]) ? 40'b0000001000001100000000000011100000001000 : 40'b0000001000001100000000000010100000001000;
													assign node1224 = (inp[12]) ? node1228 : node1225;
														assign node1225 = (inp[2]) ? 40'b0000001000000100000100000010000000001000 : 40'b1000001000000100000000000000000000001000;
														assign node1228 = (inp[2]) ? 40'b0000001000000100000000000011000000001000 : 40'b0000001000001100000000000010000000001000;
												assign node1231 = (inp[13]) ? node1239 : node1232;
													assign node1232 = (inp[2]) ? node1236 : node1233;
														assign node1233 = (inp[12]) ? 40'b0000001000001000000000000010100000001000 : 40'b1000001000000000000000000001100000001000;
														assign node1236 = (inp[12]) ? 40'b1000001000000000000000000001100000001000 : 40'b0000001000000000000100000010100000001000;
													assign node1239 = (inp[12]) ? node1243 : node1240;
														assign node1240 = (inp[2]) ? 40'b0000001000000000000100000010000000001000 : 40'b1000001000000000000000000000000000001000;
														assign node1243 = (inp[6]) ? 40'b0000001000001000000000000011000000001000 : 40'b0000001000000000000100000010000000001000;

endmodule