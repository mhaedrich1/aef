module dtc_split75_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node359;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node384;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node453;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node754;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node788;

	assign outp = (inp[9]) ? node516 : node1;
		assign node1 = (inp[6]) ? node235 : node2;
			assign node2 = (inp[10]) ? node98 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? node13 : 3'b111;
										assign node13 = (inp[5]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node53 : node18;
						assign node18 = (inp[8]) ? node34 : node19;
							assign node19 = (inp[3]) ? node21 : 3'b111;
								assign node21 = (inp[4]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? node29 : node24;
										assign node24 = (inp[1]) ? node26 : 3'b111;
											assign node26 = (inp[0]) ? 3'b011 : 3'b111;
										assign node29 = (inp[1]) ? 3'b011 : node30;
											assign node30 = (inp[0]) ? 3'b011 : 3'b111;
							assign node34 = (inp[3]) ? 3'b011 : node35;
								assign node35 = (inp[4]) ? node37 : 3'b111;
									assign node37 = (inp[5]) ? node45 : node38;
										assign node38 = (inp[0]) ? node40 : 3'b111;
											assign node40 = (inp[2]) ? 3'b011 : node41;
												assign node41 = (inp[1]) ? 3'b011 : 3'b111;
										assign node45 = (inp[0]) ? 3'b011 : node46;
											assign node46 = (inp[1]) ? 3'b011 : node47;
												assign node47 = (inp[2]) ? 3'b011 : 3'b111;
						assign node53 = (inp[8]) ? node79 : node54;
							assign node54 = (inp[4]) ? node72 : node55;
								assign node55 = (inp[3]) ? 3'b011 : node56;
									assign node56 = (inp[0]) ? node64 : node57;
										assign node57 = (inp[5]) ? node59 : 3'b111;
											assign node59 = (inp[1]) ? node61 : 3'b111;
												assign node61 = (inp[2]) ? 3'b011 : 3'b111;
										assign node64 = (inp[5]) ? 3'b011 : node65;
											assign node65 = (inp[2]) ? node67 : 3'b111;
												assign node67 = (inp[1]) ? 3'b011 : 3'b111;
								assign node72 = (inp[3]) ? node74 : 3'b011;
									assign node74 = (inp[0]) ? 3'b101 : node75;
										assign node75 = (inp[5]) ? 3'b101 : 3'b011;
							assign node79 = (inp[3]) ? node87 : node80;
								assign node80 = (inp[4]) ? node82 : 3'b011;
									assign node82 = (inp[5]) ? 3'b101 : node83;
										assign node83 = (inp[0]) ? 3'b101 : 3'b011;
								assign node87 = (inp[2]) ? node89 : 3'b101;
									assign node89 = (inp[5]) ? node91 : 3'b101;
										assign node91 = (inp[0]) ? node93 : 3'b101;
											assign node93 = (inp[1]) ? node95 : 3'b101;
												assign node95 = (inp[4]) ? 3'b001 : 3'b101;
				assign node98 = (inp[7]) ? node158 : node99;
					assign node99 = (inp[11]) ? node137 : node100;
						assign node100 = (inp[8]) ? node122 : node101;
							assign node101 = (inp[3]) ? node111 : node102;
								assign node102 = (inp[4]) ? node104 : 3'b111;
									assign node104 = (inp[1]) ? node106 : 3'b111;
										assign node106 = (inp[5]) ? node108 : 3'b111;
											assign node108 = (inp[0]) ? 3'b011 : 3'b111;
								assign node111 = (inp[2]) ? 3'b011 : node112;
									assign node112 = (inp[0]) ? 3'b011 : node113;
										assign node113 = (inp[5]) ? 3'b011 : node114;
											assign node114 = (inp[1]) ? 3'b011 : node115;
												assign node115 = (inp[4]) ? 3'b011 : 3'b111;
							assign node122 = (inp[3]) ? node124 : 3'b011;
								assign node124 = (inp[4]) ? 3'b101 : node125;
									assign node125 = (inp[0]) ? node131 : node126;
										assign node126 = (inp[5]) ? node128 : 3'b011;
											assign node128 = (inp[1]) ? 3'b101 : 3'b011;
										assign node131 = (inp[5]) ? 3'b101 : node132;
											assign node132 = (inp[2]) ? 3'b101 : 3'b011;
						assign node137 = (inp[3]) ? node147 : node138;
							assign node138 = (inp[8]) ? 3'b101 : node139;
								assign node139 = (inp[0]) ? node141 : 3'b011;
									assign node141 = (inp[4]) ? node143 : 3'b011;
										assign node143 = (inp[5]) ? 3'b101 : 3'b011;
							assign node147 = (inp[8]) ? node149 : 3'b101;
								assign node149 = (inp[4]) ? 3'b001 : node150;
									assign node150 = (inp[5]) ? 3'b001 : node151;
										assign node151 = (inp[1]) ? node153 : 3'b101;
											assign node153 = (inp[0]) ? 3'b001 : 3'b101;
					assign node158 = (inp[11]) ? node198 : node159;
						assign node159 = (inp[8]) ? node177 : node160;
							assign node160 = (inp[3]) ? node170 : node161;
								assign node161 = (inp[4]) ? 3'b101 : node162;
									assign node162 = (inp[5]) ? 3'b101 : node163;
										assign node163 = (inp[1]) ? node165 : 3'b011;
											assign node165 = (inp[0]) ? 3'b101 : 3'b011;
								assign node170 = (inp[4]) ? node172 : 3'b101;
									assign node172 = (inp[5]) ? 3'b001 : node173;
										assign node173 = (inp[0]) ? 3'b001 : 3'b101;
							assign node177 = (inp[3]) ? node189 : node178;
								assign node178 = (inp[4]) ? node184 : node179;
									assign node179 = (inp[1]) ? node181 : 3'b101;
										assign node181 = (inp[2]) ? 3'b001 : 3'b101;
									assign node184 = (inp[0]) ? 3'b001 : node185;
										assign node185 = (inp[5]) ? 3'b001 : 3'b101;
								assign node189 = (inp[5]) ? node191 : 3'b001;
									assign node191 = (inp[4]) ? node193 : 3'b001;
										assign node193 = (inp[1]) ? node195 : 3'b001;
											assign node195 = (inp[0]) ? 3'b110 : 3'b001;
						assign node198 = (inp[8]) ? node220 : node199;
							assign node199 = (inp[3]) ? node207 : node200;
								assign node200 = (inp[4]) ? 3'b001 : node201;
									assign node201 = (inp[0]) ? 3'b001 : node202;
										assign node202 = (inp[5]) ? 3'b001 : 3'b101;
								assign node207 = (inp[4]) ? node215 : node208;
									assign node208 = (inp[5]) ? node210 : 3'b001;
										assign node210 = (inp[0]) ? node212 : 3'b001;
											assign node212 = (inp[1]) ? 3'b110 : 3'b001;
									assign node215 = (inp[0]) ? 3'b110 : node216;
										assign node216 = (inp[5]) ? 3'b110 : 3'b001;
							assign node220 = (inp[3]) ? node228 : node221;
								assign node221 = (inp[4]) ? 3'b110 : node222;
									assign node222 = (inp[1]) ? node224 : 3'b001;
										assign node224 = (inp[0]) ? 3'b110 : 3'b001;
								assign node228 = (inp[5]) ? node230 : 3'b110;
									assign node230 = (inp[4]) ? node232 : 3'b110;
										assign node232 = (inp[0]) ? 3'b010 : 3'b110;
			assign node235 = (inp[10]) ? node393 : node236;
				assign node236 = (inp[7]) ? node300 : node237;
					assign node237 = (inp[11]) ? node267 : node238;
						assign node238 = (inp[8]) ? node248 : node239;
							assign node239 = (inp[3]) ? node241 : 3'b011;
								assign node241 = (inp[4]) ? 3'b101 : node242;
									assign node242 = (inp[0]) ? 3'b101 : node243;
										assign node243 = (inp[5]) ? 3'b101 : 3'b011;
							assign node248 = (inp[3]) ? node260 : node249;
								assign node249 = (inp[2]) ? 3'b101 : node250;
									assign node250 = (inp[1]) ? 3'b101 : node251;
										assign node251 = (inp[5]) ? 3'b101 : node252;
											assign node252 = (inp[0]) ? 3'b101 : node253;
												assign node253 = (inp[4]) ? 3'b101 : 3'b011;
								assign node260 = (inp[4]) ? 3'b001 : node261;
									assign node261 = (inp[0]) ? node263 : 3'b101;
										assign node263 = (inp[5]) ? 3'b001 : 3'b101;
						assign node267 = (inp[8]) ? node289 : node268;
							assign node268 = (inp[3]) ? node280 : node269;
								assign node269 = (inp[4]) ? node271 : 3'b101;
									assign node271 = (inp[0]) ? node273 : 3'b101;
										assign node273 = (inp[5]) ? node275 : 3'b101;
											assign node275 = (inp[1]) ? 3'b001 : node276;
												assign node276 = (inp[2]) ? 3'b001 : 3'b101;
								assign node280 = (inp[5]) ? 3'b001 : node281;
									assign node281 = (inp[0]) ? 3'b001 : node282;
										assign node282 = (inp[2]) ? 3'b001 : node283;
											assign node283 = (inp[4]) ? 3'b001 : 3'b101;
							assign node289 = (inp[3]) ? node291 : 3'b001;
								assign node291 = (inp[5]) ? 3'b110 : node292;
									assign node292 = (inp[4]) ? 3'b110 : node293;
										assign node293 = (inp[0]) ? node295 : 3'b001;
											assign node295 = (inp[2]) ? 3'b110 : 3'b001;
					assign node300 = (inp[11]) ? node340 : node301;
						assign node301 = (inp[8]) ? node323 : node302;
							assign node302 = (inp[4]) ? node316 : node303;
								assign node303 = (inp[3]) ? 3'b001 : node304;
									assign node304 = (inp[5]) ? node310 : node305;
										assign node305 = (inp[0]) ? node307 : 3'b101;
											assign node307 = (inp[2]) ? 3'b001 : 3'b101;
										assign node310 = (inp[0]) ? 3'b001 : node311;
											assign node311 = (inp[1]) ? 3'b001 : 3'b101;
								assign node316 = (inp[3]) ? node318 : 3'b001;
									assign node318 = (inp[5]) ? 3'b110 : node319;
										assign node319 = (inp[0]) ? 3'b110 : 3'b001;
							assign node323 = (inp[3]) ? node331 : node324;
								assign node324 = (inp[4]) ? node326 : 3'b001;
									assign node326 = (inp[0]) ? 3'b110 : node327;
										assign node327 = (inp[5]) ? 3'b110 : 3'b001;
								assign node331 = (inp[4]) ? node333 : 3'b110;
									assign node333 = (inp[5]) ? node335 : 3'b110;
										assign node335 = (inp[1]) ? node337 : 3'b110;
											assign node337 = (inp[0]) ? 3'b010 : 3'b110;
						assign node340 = (inp[8]) ? node366 : node341;
							assign node341 = (inp[3]) ? node359 : node342;
								assign node342 = (inp[4]) ? 3'b110 : node343;
									assign node343 = (inp[5]) ? node351 : node344;
										assign node344 = (inp[0]) ? node346 : 3'b001;
											assign node346 = (inp[1]) ? 3'b110 : node347;
												assign node347 = (inp[2]) ? 3'b110 : 3'b001;
										assign node351 = (inp[0]) ? 3'b110 : node352;
											assign node352 = (inp[2]) ? 3'b110 : node353;
												assign node353 = (inp[1]) ? 3'b110 : 3'b001;
								assign node359 = (inp[4]) ? node361 : 3'b110;
									assign node361 = (inp[0]) ? 3'b010 : node362;
										assign node362 = (inp[5]) ? 3'b010 : 3'b110;
							assign node366 = (inp[3]) ? node384 : node367;
								assign node367 = (inp[4]) ? node377 : node368;
									assign node368 = (inp[5]) ? node370 : 3'b110;
										assign node370 = (inp[2]) ? node372 : 3'b110;
											assign node372 = (inp[1]) ? node374 : 3'b110;
												assign node374 = (inp[0]) ? 3'b010 : 3'b110;
									assign node377 = (inp[1]) ? 3'b010 : node378;
										assign node378 = (inp[0]) ? 3'b010 : node379;
											assign node379 = (inp[5]) ? 3'b010 : 3'b110;
								assign node384 = (inp[4]) ? node386 : 3'b010;
									assign node386 = (inp[0]) ? node388 : 3'b010;
										assign node388 = (inp[1]) ? 3'b100 : node389;
											assign node389 = (inp[2]) ? 3'b100 : 3'b010;
				assign node393 = (inp[7]) ? node443 : node394;
					assign node394 = (inp[11]) ? node420 : node395;
						assign node395 = (inp[3]) ? node405 : node396;
							assign node396 = (inp[8]) ? 3'b110 : node397;
								assign node397 = (inp[4]) ? node399 : 3'b001;
									assign node399 = (inp[0]) ? node401 : 3'b001;
										assign node401 = (inp[5]) ? 3'b110 : 3'b001;
							assign node405 = (inp[8]) ? node407 : 3'b110;
								assign node407 = (inp[4]) ? 3'b010 : node408;
									assign node408 = (inp[1]) ? node414 : node409;
										assign node409 = (inp[2]) ? node411 : 3'b110;
											assign node411 = (inp[0]) ? 3'b010 : 3'b110;
										assign node414 = (inp[5]) ? 3'b010 : node415;
											assign node415 = (inp[0]) ? 3'b010 : 3'b110;
						assign node420 = (inp[3]) ? node434 : node421;
							assign node421 = (inp[8]) ? 3'b010 : node422;
								assign node422 = (inp[0]) ? node424 : 3'b110;
									assign node424 = (inp[4]) ? node426 : 3'b110;
										assign node426 = (inp[5]) ? 3'b010 : node427;
											assign node427 = (inp[1]) ? node429 : 3'b110;
												assign node429 = (inp[2]) ? 3'b010 : 3'b110;
							assign node434 = (inp[8]) ? node436 : 3'b010;
								assign node436 = (inp[4]) ? 3'b100 : node437;
									assign node437 = (inp[5]) ? 3'b100 : node438;
										assign node438 = (inp[0]) ? 3'b100 : 3'b010;
					assign node443 = (inp[11]) ? node481 : node444;
						assign node444 = (inp[8]) ? node464 : node445;
							assign node445 = (inp[4]) ? node453 : node446;
								assign node446 = (inp[5]) ? 3'b010 : node447;
									assign node447 = (inp[3]) ? 3'b010 : node448;
										assign node448 = (inp[0]) ? 3'b010 : 3'b110;
								assign node453 = (inp[3]) ? node455 : 3'b010;
									assign node455 = (inp[5]) ? 3'b100 : node456;
										assign node456 = (inp[0]) ? 3'b100 : node457;
											assign node457 = (inp[1]) ? node459 : 3'b010;
												assign node459 = (inp[2]) ? 3'b100 : 3'b010;
							assign node464 = (inp[3]) ? node474 : node465;
								assign node465 = (inp[4]) ? 3'b100 : node466;
									assign node466 = (inp[5]) ? node468 : 3'b010;
										assign node468 = (inp[0]) ? node470 : 3'b010;
											assign node470 = (inp[2]) ? 3'b100 : 3'b010;
								assign node474 = (inp[0]) ? node476 : 3'b100;
									assign node476 = (inp[4]) ? node478 : 3'b100;
										assign node478 = (inp[5]) ? 3'b000 : 3'b100;
						assign node481 = (inp[8]) ? node507 : node482;
							assign node482 = (inp[3]) ? node494 : node483;
								assign node483 = (inp[0]) ? 3'b100 : node484;
									assign node484 = (inp[4]) ? 3'b100 : node485;
										assign node485 = (inp[5]) ? 3'b100 : node486;
											assign node486 = (inp[1]) ? node488 : 3'b010;
												assign node488 = (inp[2]) ? 3'b100 : 3'b010;
								assign node494 = (inp[4]) ? node500 : node495;
									assign node495 = (inp[5]) ? node497 : 3'b100;
										assign node497 = (inp[0]) ? 3'b000 : 3'b100;
									assign node500 = (inp[1]) ? 3'b000 : node501;
										assign node501 = (inp[2]) ? 3'b000 : node502;
											assign node502 = (inp[5]) ? 3'b000 : 3'b100;
							assign node507 = (inp[4]) ? 3'b000 : node508;
								assign node508 = (inp[3]) ? 3'b000 : node509;
									assign node509 = (inp[0]) ? node511 : 3'b100;
										assign node511 = (inp[5]) ? 3'b000 : 3'b100;
		assign node516 = (inp[6]) ? node744 : node517;
			assign node517 = (inp[10]) ? node647 : node518;
				assign node518 = (inp[7]) ? node562 : node519;
					assign node519 = (inp[11]) ? node539 : node520;
						assign node520 = (inp[3]) ? node530 : node521;
							assign node521 = (inp[8]) ? 3'b001 : node522;
								assign node522 = (inp[4]) ? node524 : 3'b101;
									assign node524 = (inp[5]) ? node526 : 3'b101;
										assign node526 = (inp[0]) ? 3'b001 : 3'b101;
							assign node530 = (inp[8]) ? node532 : 3'b001;
								assign node532 = (inp[5]) ? 3'b110 : node533;
									assign node533 = (inp[4]) ? 3'b110 : node534;
										assign node534 = (inp[1]) ? 3'b110 : 3'b001;
						assign node539 = (inp[3]) ? node551 : node540;
							assign node540 = (inp[8]) ? 3'b110 : node541;
								assign node541 = (inp[4]) ? node543 : 3'b001;
									assign node543 = (inp[1]) ? 3'b110 : node544;
										assign node544 = (inp[5]) ? node546 : 3'b001;
											assign node546 = (inp[0]) ? 3'b110 : 3'b001;
							assign node551 = (inp[8]) ? node553 : 3'b110;
								assign node553 = (inp[0]) ? 3'b010 : node554;
									assign node554 = (inp[4]) ? 3'b010 : node555;
										assign node555 = (inp[5]) ? 3'b010 : node556;
											assign node556 = (inp[1]) ? 3'b010 : 3'b110;
					assign node562 = (inp[11]) ? node610 : node563;
						assign node563 = (inp[8]) ? node591 : node564;
							assign node564 = (inp[3]) ? node576 : node565;
								assign node565 = (inp[4]) ? 3'b110 : node566;
									assign node566 = (inp[0]) ? 3'b110 : node567;
										assign node567 = (inp[5]) ? 3'b110 : node568;
											assign node568 = (inp[2]) ? node570 : 3'b001;
												assign node570 = (inp[1]) ? 3'b110 : 3'b001;
								assign node576 = (inp[4]) ? node584 : node577;
									assign node577 = (inp[1]) ? node579 : 3'b110;
										assign node579 = (inp[0]) ? node581 : 3'b110;
											assign node581 = (inp[5]) ? 3'b010 : 3'b110;
									assign node584 = (inp[5]) ? 3'b010 : node585;
										assign node585 = (inp[0]) ? 3'b010 : node586;
											assign node586 = (inp[1]) ? 3'b010 : 3'b110;
							assign node591 = (inp[3]) ? node599 : node592;
								assign node592 = (inp[4]) ? 3'b010 : node593;
									assign node593 = (inp[5]) ? node595 : 3'b110;
										assign node595 = (inp[0]) ? 3'b010 : 3'b110;
								assign node599 = (inp[4]) ? node601 : 3'b010;
									assign node601 = (inp[5]) ? node603 : 3'b010;
										assign node603 = (inp[0]) ? 3'b100 : node604;
											assign node604 = (inp[1]) ? node606 : 3'b010;
												assign node606 = (inp[2]) ? 3'b100 : 3'b010;
						assign node610 = (inp[8]) ? node622 : node611;
							assign node611 = (inp[3]) ? node613 : 3'b010;
								assign node613 = (inp[4]) ? 3'b100 : node614;
									assign node614 = (inp[5]) ? node616 : 3'b010;
										assign node616 = (inp[0]) ? node618 : 3'b010;
											assign node618 = (inp[1]) ? 3'b100 : 3'b010;
							assign node622 = (inp[4]) ? node634 : node623;
								assign node623 = (inp[3]) ? 3'b100 : node624;
									assign node624 = (inp[5]) ? node626 : 3'b010;
										assign node626 = (inp[0]) ? 3'b100 : node627;
											assign node627 = (inp[1]) ? node629 : 3'b010;
												assign node629 = (inp[2]) ? 3'b100 : 3'b010;
								assign node634 = (inp[3]) ? node636 : 3'b100;
									assign node636 = (inp[0]) ? node642 : node637;
										assign node637 = (inp[5]) ? node639 : 3'b100;
											assign node639 = (inp[1]) ? 3'b000 : 3'b100;
										assign node642 = (inp[1]) ? 3'b000 : node643;
											assign node643 = (inp[5]) ? 3'b000 : 3'b100;
				assign node647 = (inp[7]) ? node715 : node648;
					assign node648 = (inp[11]) ? node686 : node649;
						assign node649 = (inp[8]) ? node667 : node650;
							assign node650 = (inp[3]) ? 3'b010 : node651;
								assign node651 = (inp[4]) ? node653 : 3'b110;
									assign node653 = (inp[0]) ? node659 : node654;
										assign node654 = (inp[1]) ? node656 : 3'b110;
											assign node656 = (inp[5]) ? 3'b010 : 3'b110;
										assign node659 = (inp[5]) ? 3'b010 : node660;
											assign node660 = (inp[2]) ? 3'b010 : node661;
												assign node661 = (inp[1]) ? 3'b010 : 3'b110;
							assign node667 = (inp[3]) ? node677 : node668;
								assign node668 = (inp[0]) ? node670 : 3'b010;
									assign node670 = (inp[1]) ? node672 : 3'b010;
										assign node672 = (inp[4]) ? node674 : 3'b010;
											assign node674 = (inp[5]) ? 3'b100 : 3'b010;
								assign node677 = (inp[4]) ? 3'b100 : node678;
									assign node678 = (inp[5]) ? 3'b100 : node679;
										assign node679 = (inp[1]) ? 3'b100 : node680;
											assign node680 = (inp[0]) ? 3'b100 : 3'b010;
						assign node686 = (inp[8]) ? node696 : node687;
							assign node687 = (inp[3]) ? 3'b100 : node688;
								assign node688 = (inp[4]) ? node690 : 3'b010;
									assign node690 = (inp[5]) ? 3'b100 : node691;
										assign node691 = (inp[0]) ? 3'b100 : 3'b010;
							assign node696 = (inp[3]) ? node704 : node697;
								assign node697 = (inp[0]) ? node699 : 3'b100;
									assign node699 = (inp[5]) ? node701 : 3'b100;
										assign node701 = (inp[4]) ? 3'b000 : 3'b100;
								assign node704 = (inp[2]) ? 3'b000 : node705;
									assign node705 = (inp[0]) ? 3'b000 : node706;
										assign node706 = (inp[1]) ? 3'b000 : node707;
											assign node707 = (inp[5]) ? 3'b000 : node708;
												assign node708 = (inp[4]) ? 3'b000 : 3'b100;
					assign node715 = (inp[11]) ? 3'b000 : node716;
						assign node716 = (inp[8]) ? node728 : node717;
							assign node717 = (inp[3]) ? node719 : 3'b100;
								assign node719 = (inp[4]) ? 3'b000 : node720;
									assign node720 = (inp[5]) ? node722 : 3'b100;
										assign node722 = (inp[0]) ? 3'b000 : node723;
											assign node723 = (inp[1]) ? 3'b000 : 3'b100;
							assign node728 = (inp[3]) ? 3'b000 : node729;
								assign node729 = (inp[4]) ? 3'b000 : node730;
									assign node730 = (inp[0]) ? node736 : node731;
										assign node731 = (inp[5]) ? node733 : 3'b100;
											assign node733 = (inp[2]) ? 3'b000 : 3'b100;
										assign node736 = (inp[1]) ? 3'b000 : node737;
											assign node737 = (inp[5]) ? 3'b000 : 3'b100;
			assign node744 = (inp[7]) ? 3'b000 : node745;
				assign node745 = (inp[10]) ? 3'b000 : node746;
					assign node746 = (inp[11]) ? node780 : node747;
						assign node747 = (inp[8]) ? node763 : node748;
							assign node748 = (inp[3]) ? 3'b100 : node749;
								assign node749 = (inp[4]) ? node751 : 3'b010;
									assign node751 = (inp[5]) ? node757 : node752;
										assign node752 = (inp[1]) ? node754 : 3'b010;
											assign node754 = (inp[0]) ? 3'b100 : 3'b010;
										assign node757 = (inp[0]) ? 3'b100 : node758;
											assign node758 = (inp[1]) ? 3'b100 : 3'b010;
							assign node763 = (inp[3]) ? node773 : node764;
								assign node764 = (inp[5]) ? node766 : 3'b100;
									assign node766 = (inp[4]) ? node768 : 3'b100;
										assign node768 = (inp[2]) ? node770 : 3'b100;
											assign node770 = (inp[1]) ? 3'b000 : 3'b100;
								assign node773 = (inp[0]) ? 3'b000 : node774;
									assign node774 = (inp[5]) ? 3'b000 : node775;
										assign node775 = (inp[4]) ? 3'b000 : 3'b100;
						assign node780 = (inp[8]) ? 3'b000 : node781;
							assign node781 = (inp[3]) ? 3'b000 : node782;
								assign node782 = (inp[4]) ? node784 : 3'b100;
									assign node784 = (inp[5]) ? 3'b000 : node785;
										assign node785 = (inp[0]) ? node787 : 3'b100;
											assign node787 = (inp[1]) ? 3'b000 : node788;
												assign node788 = (inp[2]) ? 3'b000 : 3'b100;

endmodule