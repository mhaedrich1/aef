module dtc_split66_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node414;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node693;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;

	assign outp = (inp[9]) ? node456 : node1;
		assign node1 = (inp[6]) ? node195 : node2;
			assign node2 = (inp[10]) ? node80 : node3;
				assign node3 = (inp[7]) ? node15 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? 3'b011 : 3'b111;
					assign node15 = (inp[11]) ? node43 : node16;
						assign node16 = (inp[8]) ? node28 : node17;
							assign node17 = (inp[4]) ? node19 : 3'b111;
								assign node19 = (inp[3]) ? node21 : 3'b111;
									assign node21 = (inp[5]) ? node23 : 3'b111;
										assign node23 = (inp[0]) ? 3'b011 : node24;
											assign node24 = (inp[1]) ? 3'b011 : 3'b111;
							assign node28 = (inp[3]) ? 3'b011 : node29;
								assign node29 = (inp[4]) ? node31 : 3'b111;
									assign node31 = (inp[0]) ? node37 : node32;
										assign node32 = (inp[1]) ? node34 : 3'b111;
											assign node34 = (inp[5]) ? 3'b011 : 3'b111;
										assign node37 = (inp[2]) ? 3'b011 : node38;
											assign node38 = (inp[5]) ? 3'b011 : 3'b111;
						assign node43 = (inp[3]) ? node61 : node44;
							assign node44 = (inp[4]) ? node54 : node45;
								assign node45 = (inp[8]) ? 3'b011 : node46;
									assign node46 = (inp[0]) ? node48 : 3'b111;
										assign node48 = (inp[5]) ? 3'b011 : node49;
											assign node49 = (inp[1]) ? 3'b011 : 3'b111;
								assign node54 = (inp[8]) ? node56 : 3'b011;
									assign node56 = (inp[0]) ? 3'b101 : node57;
										assign node57 = (inp[5]) ? 3'b101 : 3'b011;
							assign node61 = (inp[8]) ? node69 : node62;
								assign node62 = (inp[4]) ? node64 : 3'b011;
									assign node64 = (inp[5]) ? 3'b101 : node65;
										assign node65 = (inp[0]) ? 3'b101 : 3'b011;
								assign node69 = (inp[2]) ? node71 : 3'b101;
									assign node71 = (inp[1]) ? node73 : 3'b101;
										assign node73 = (inp[5]) ? node75 : 3'b101;
											assign node75 = (inp[0]) ? node77 : 3'b101;
												assign node77 = (inp[4]) ? 3'b001 : 3'b101;
				assign node80 = (inp[7]) ? node118 : node81;
					assign node81 = (inp[11]) ? node97 : node82;
						assign node82 = (inp[3]) ? node86 : node83;
							assign node83 = (inp[8]) ? 3'b011 : 3'b111;
							assign node86 = (inp[8]) ? node88 : 3'b011;
								assign node88 = (inp[4]) ? 3'b101 : node89;
									assign node89 = (inp[0]) ? node91 : 3'b011;
										assign node91 = (inp[5]) ? 3'b101 : node92;
											assign node92 = (inp[2]) ? 3'b101 : 3'b011;
						assign node97 = (inp[3]) ? node107 : node98;
							assign node98 = (inp[8]) ? 3'b101 : node99;
								assign node99 = (inp[0]) ? node101 : 3'b011;
									assign node101 = (inp[4]) ? node103 : 3'b011;
										assign node103 = (inp[5]) ? 3'b101 : 3'b011;
							assign node107 = (inp[8]) ? node109 : 3'b101;
								assign node109 = (inp[4]) ? 3'b001 : node110;
									assign node110 = (inp[5]) ? 3'b001 : node111;
										assign node111 = (inp[0]) ? node113 : 3'b101;
											assign node113 = (inp[1]) ? 3'b001 : 3'b101;
					assign node118 = (inp[11]) ? node160 : node119;
						assign node119 = (inp[3]) ? node145 : node120;
							assign node120 = (inp[8]) ? node130 : node121;
								assign node121 = (inp[4]) ? 3'b101 : node122;
									assign node122 = (inp[0]) ? node124 : 3'b011;
										assign node124 = (inp[1]) ? 3'b101 : node125;
											assign node125 = (inp[5]) ? 3'b101 : 3'b011;
								assign node130 = (inp[4]) ? node138 : node131;
									assign node131 = (inp[5]) ? node133 : 3'b101;
										assign node133 = (inp[2]) ? node135 : 3'b101;
											assign node135 = (inp[1]) ? 3'b001 : 3'b101;
									assign node138 = (inp[5]) ? 3'b001 : node139;
										assign node139 = (inp[2]) ? 3'b001 : node140;
											assign node140 = (inp[0]) ? 3'b001 : 3'b101;
							assign node145 = (inp[8]) ? node149 : node146;
								assign node146 = (inp[4]) ? 3'b001 : 3'b101;
								assign node149 = (inp[5]) ? node151 : 3'b001;
									assign node151 = (inp[2]) ? node153 : 3'b001;
										assign node153 = (inp[1]) ? node155 : 3'b001;
											assign node155 = (inp[0]) ? node157 : 3'b001;
												assign node157 = (inp[4]) ? 3'b110 : 3'b001;
						assign node160 = (inp[8]) ? node178 : node161;
							assign node161 = (inp[3]) ? node169 : node162;
								assign node162 = (inp[5]) ? 3'b001 : node163;
									assign node163 = (inp[0]) ? 3'b001 : node164;
										assign node164 = (inp[4]) ? 3'b001 : 3'b101;
								assign node169 = (inp[4]) ? node171 : 3'b001;
									assign node171 = (inp[0]) ? 3'b110 : node172;
										assign node172 = (inp[2]) ? 3'b110 : node173;
											assign node173 = (inp[5]) ? 3'b110 : 3'b001;
							assign node178 = (inp[3]) ? node188 : node179;
								assign node179 = (inp[4]) ? 3'b110 : node180;
									assign node180 = (inp[0]) ? node182 : 3'b001;
										assign node182 = (inp[5]) ? node184 : 3'b001;
											assign node184 = (inp[1]) ? 3'b110 : 3'b001;
								assign node188 = (inp[4]) ? node190 : 3'b110;
									assign node190 = (inp[5]) ? node192 : 3'b110;
										assign node192 = (inp[0]) ? 3'b010 : 3'b110;
			assign node195 = (inp[10]) ? node335 : node196;
				assign node196 = (inp[7]) ? node252 : node197;
					assign node197 = (inp[11]) ? node219 : node198;
						assign node198 = (inp[8]) ? node210 : node199;
							assign node199 = (inp[3]) ? node201 : 3'b011;
								assign node201 = (inp[0]) ? 3'b101 : node202;
									assign node202 = (inp[1]) ? 3'b101 : node203;
										assign node203 = (inp[5]) ? 3'b101 : node204;
											assign node204 = (inp[4]) ? 3'b101 : 3'b011;
							assign node210 = (inp[3]) ? node212 : 3'b101;
								assign node212 = (inp[4]) ? 3'b001 : node213;
									assign node213 = (inp[5]) ? node215 : 3'b101;
										assign node215 = (inp[0]) ? 3'b001 : 3'b101;
						assign node219 = (inp[8]) ? node241 : node220;
							assign node220 = (inp[3]) ? node230 : node221;
								assign node221 = (inp[4]) ? node223 : 3'b101;
									assign node223 = (inp[0]) ? node225 : 3'b101;
										assign node225 = (inp[5]) ? node227 : 3'b101;
											assign node227 = (inp[1]) ? 3'b001 : 3'b101;
								assign node230 = (inp[2]) ? 3'b001 : node231;
									assign node231 = (inp[4]) ? 3'b001 : node232;
										assign node232 = (inp[1]) ? 3'b001 : node233;
											assign node233 = (inp[5]) ? 3'b001 : node234;
												assign node234 = (inp[0]) ? 3'b001 : 3'b101;
							assign node241 = (inp[3]) ? node243 : 3'b001;
								assign node243 = (inp[4]) ? 3'b110 : node244;
									assign node244 = (inp[5]) ? node246 : 3'b001;
										assign node246 = (inp[0]) ? 3'b110 : node247;
											assign node247 = (inp[1]) ? 3'b110 : 3'b001;
					assign node252 = (inp[11]) ? node296 : node253;
						assign node253 = (inp[8]) ? node279 : node254;
							assign node254 = (inp[3]) ? node264 : node255;
								assign node255 = (inp[4]) ? 3'b001 : node256;
									assign node256 = (inp[5]) ? node258 : 3'b101;
										assign node258 = (inp[1]) ? 3'b001 : node259;
											assign node259 = (inp[0]) ? 3'b001 : 3'b101;
								assign node264 = (inp[4]) ? node266 : 3'b001;
									assign node266 = (inp[0]) ? node272 : node267;
										assign node267 = (inp[5]) ? node269 : 3'b001;
											assign node269 = (inp[2]) ? 3'b110 : 3'b001;
										assign node272 = (inp[5]) ? 3'b110 : node273;
											assign node273 = (inp[2]) ? 3'b110 : node274;
												assign node274 = (inp[1]) ? 3'b110 : 3'b001;
							assign node279 = (inp[3]) ? node287 : node280;
								assign node280 = (inp[4]) ? node282 : 3'b001;
									assign node282 = (inp[5]) ? 3'b110 : node283;
										assign node283 = (inp[0]) ? 3'b110 : 3'b001;
								assign node287 = (inp[5]) ? node289 : 3'b110;
									assign node289 = (inp[0]) ? node291 : 3'b110;
										assign node291 = (inp[1]) ? node293 : 3'b110;
											assign node293 = (inp[4]) ? 3'b010 : 3'b110;
						assign node296 = (inp[8]) ? node316 : node297;
							assign node297 = (inp[0]) ? node311 : node298;
								assign node298 = (inp[4]) ? node306 : node299;
									assign node299 = (inp[3]) ? 3'b110 : node300;
										assign node300 = (inp[5]) ? node302 : 3'b001;
											assign node302 = (inp[1]) ? 3'b110 : 3'b001;
									assign node306 = (inp[5]) ? node308 : 3'b110;
										assign node308 = (inp[3]) ? 3'b010 : 3'b110;
								assign node311 = (inp[3]) ? node313 : 3'b110;
									assign node313 = (inp[4]) ? 3'b010 : 3'b110;
							assign node316 = (inp[4]) ? node320 : node317;
								assign node317 = (inp[3]) ? 3'b010 : 3'b110;
								assign node320 = (inp[2]) ? node322 : 3'b010;
									assign node322 = (inp[5]) ? node330 : node323;
										assign node323 = (inp[3]) ? 3'b010 : node324;
											assign node324 = (inp[1]) ? 3'b010 : node325;
												assign node325 = (inp[0]) ? 3'b010 : 3'b110;
										assign node330 = (inp[0]) ? node332 : 3'b010;
											assign node332 = (inp[3]) ? 3'b100 : 3'b010;
				assign node335 = (inp[7]) ? node379 : node336;
					assign node336 = (inp[11]) ? node360 : node337;
						assign node337 = (inp[3]) ? node347 : node338;
							assign node338 = (inp[8]) ? 3'b110 : node339;
								assign node339 = (inp[4]) ? node341 : 3'b001;
									assign node341 = (inp[5]) ? node343 : 3'b001;
										assign node343 = (inp[0]) ? 3'b110 : 3'b001;
							assign node347 = (inp[8]) ? node349 : 3'b110;
								assign node349 = (inp[4]) ? 3'b010 : node350;
									assign node350 = (inp[1]) ? node354 : node351;
										assign node351 = (inp[2]) ? 3'b010 : 3'b110;
										assign node354 = (inp[0]) ? 3'b010 : node355;
											assign node355 = (inp[2]) ? 3'b110 : 3'b010;
						assign node360 = (inp[3]) ? node370 : node361;
							assign node361 = (inp[8]) ? 3'b010 : node362;
								assign node362 = (inp[0]) ? node364 : 3'b110;
									assign node364 = (inp[4]) ? node366 : 3'b110;
										assign node366 = (inp[5]) ? 3'b010 : 3'b110;
							assign node370 = (inp[8]) ? node372 : 3'b010;
								assign node372 = (inp[4]) ? 3'b100 : node373;
									assign node373 = (inp[0]) ? 3'b100 : node374;
										assign node374 = (inp[5]) ? 3'b100 : 3'b010;
					assign node379 = (inp[11]) ? node421 : node380;
						assign node380 = (inp[8]) ? node400 : node381;
							assign node381 = (inp[3]) ? node389 : node382;
								assign node382 = (inp[0]) ? 3'b010 : node383;
									assign node383 = (inp[4]) ? 3'b010 : node384;
										assign node384 = (inp[5]) ? 3'b010 : 3'b110;
								assign node389 = (inp[4]) ? node391 : 3'b010;
									assign node391 = (inp[0]) ? 3'b100 : node392;
										assign node392 = (inp[5]) ? 3'b100 : node393;
											assign node393 = (inp[2]) ? node395 : 3'b010;
												assign node395 = (inp[1]) ? 3'b100 : 3'b010;
							assign node400 = (inp[3]) ? node414 : node401;
								assign node401 = (inp[4]) ? node407 : node402;
									assign node402 = (inp[5]) ? node404 : 3'b010;
										assign node404 = (inp[0]) ? 3'b100 : 3'b010;
									assign node407 = (inp[2]) ? 3'b100 : node408;
										assign node408 = (inp[5]) ? 3'b100 : node409;
											assign node409 = (inp[0]) ? 3'b100 : 3'b010;
								assign node414 = (inp[4]) ? node416 : 3'b100;
									assign node416 = (inp[5]) ? node418 : 3'b100;
										assign node418 = (inp[0]) ? 3'b000 : 3'b100;
						assign node421 = (inp[8]) ? node447 : node422;
							assign node422 = (inp[3]) ? node432 : node423;
								assign node423 = (inp[4]) ? 3'b100 : node424;
									assign node424 = (inp[0]) ? 3'b100 : node425;
										assign node425 = (inp[5]) ? 3'b100 : node426;
											assign node426 = (inp[2]) ? 3'b100 : 3'b010;
								assign node432 = (inp[4]) ? node440 : node433;
									assign node433 = (inp[0]) ? node435 : 3'b100;
										assign node435 = (inp[5]) ? node437 : 3'b100;
											assign node437 = (inp[2]) ? 3'b100 : 3'b000;
									assign node440 = (inp[1]) ? 3'b000 : node441;
										assign node441 = (inp[5]) ? 3'b000 : node442;
											assign node442 = (inp[2]) ? 3'b000 : 3'b100;
							assign node447 = (inp[3]) ? 3'b000 : node448;
								assign node448 = (inp[4]) ? 3'b000 : node449;
									assign node449 = (inp[5]) ? node451 : 3'b100;
										assign node451 = (inp[0]) ? 3'b000 : 3'b100;
		assign node456 = (inp[6]) ? node674 : node457;
			assign node457 = (inp[10]) ? node577 : node458;
				assign node458 = (inp[7]) ? node502 : node459;
					assign node459 = (inp[11]) ? node481 : node460;
						assign node460 = (inp[3]) ? node472 : node461;
							assign node461 = (inp[8]) ? 3'b001 : node462;
								assign node462 = (inp[5]) ? node464 : 3'b101;
									assign node464 = (inp[4]) ? node466 : 3'b101;
										assign node466 = (inp[0]) ? 3'b001 : node467;
											assign node467 = (inp[1]) ? 3'b001 : 3'b101;
							assign node472 = (inp[8]) ? node474 : 3'b001;
								assign node474 = (inp[4]) ? 3'b110 : node475;
									assign node475 = (inp[2]) ? 3'b110 : node476;
										assign node476 = (inp[5]) ? 3'b110 : 3'b001;
						assign node481 = (inp[8]) ? node493 : node482;
							assign node482 = (inp[3]) ? 3'b110 : node483;
								assign node483 = (inp[1]) ? node485 : 3'b001;
									assign node485 = (inp[4]) ? node487 : 3'b001;
										assign node487 = (inp[0]) ? 3'b110 : node488;
											assign node488 = (inp[5]) ? 3'b110 : 3'b001;
							assign node493 = (inp[3]) ? node495 : 3'b110;
								assign node495 = (inp[4]) ? 3'b010 : node496;
									assign node496 = (inp[0]) ? 3'b010 : node497;
										assign node497 = (inp[5]) ? 3'b010 : 3'b110;
					assign node502 = (inp[11]) ? node540 : node503;
						assign node503 = (inp[8]) ? node521 : node504;
							assign node504 = (inp[3]) ? node514 : node505;
								assign node505 = (inp[0]) ? 3'b110 : node506;
									assign node506 = (inp[4]) ? 3'b110 : node507;
										assign node507 = (inp[2]) ? node509 : 3'b001;
											assign node509 = (inp[1]) ? 3'b110 : 3'b001;
								assign node514 = (inp[4]) ? node516 : 3'b110;
									assign node516 = (inp[1]) ? 3'b010 : node517;
										assign node517 = (inp[0]) ? 3'b010 : 3'b110;
							assign node521 = (inp[4]) ? node531 : node522;
								assign node522 = (inp[3]) ? 3'b010 : node523;
									assign node523 = (inp[5]) ? node525 : 3'b110;
										assign node525 = (inp[0]) ? node527 : 3'b110;
											assign node527 = (inp[1]) ? 3'b010 : 3'b110;
								assign node531 = (inp[3]) ? node533 : 3'b010;
									assign node533 = (inp[5]) ? node535 : 3'b010;
										assign node535 = (inp[0]) ? 3'b100 : node536;
											assign node536 = (inp[2]) ? 3'b100 : 3'b010;
						assign node540 = (inp[8]) ? node560 : node541;
							assign node541 = (inp[3]) ? node549 : node542;
								assign node542 = (inp[4]) ? 3'b010 : node543;
									assign node543 = (inp[5]) ? 3'b010 : node544;
										assign node544 = (inp[0]) ? 3'b010 : 3'b110;
								assign node549 = (inp[4]) ? 3'b100 : node550;
									assign node550 = (inp[5]) ? node552 : 3'b010;
										assign node552 = (inp[0]) ? node554 : 3'b010;
											assign node554 = (inp[2]) ? 3'b100 : node555;
												assign node555 = (inp[1]) ? 3'b100 : 3'b010;
							assign node560 = (inp[4]) ? node572 : node561;
								assign node561 = (inp[3]) ? 3'b100 : node562;
									assign node562 = (inp[5]) ? node564 : 3'b010;
										assign node564 = (inp[0]) ? 3'b100 : node565;
											assign node565 = (inp[1]) ? node567 : 3'b010;
												assign node567 = (inp[2]) ? 3'b100 : 3'b010;
								assign node572 = (inp[3]) ? node574 : 3'b100;
									assign node574 = (inp[1]) ? 3'b000 : 3'b100;
				assign node577 = (inp[7]) ? node643 : node578;
					assign node578 = (inp[11]) ? node606 : node579;
						assign node579 = (inp[8]) ? node589 : node580;
							assign node580 = (inp[3]) ? 3'b010 : node581;
								assign node581 = (inp[4]) ? node583 : 3'b110;
									assign node583 = (inp[5]) ? 3'b010 : node584;
										assign node584 = (inp[0]) ? 3'b010 : 3'b110;
							assign node589 = (inp[3]) ? node599 : node590;
								assign node590 = (inp[4]) ? node592 : 3'b010;
									assign node592 = (inp[5]) ? node594 : 3'b010;
										assign node594 = (inp[0]) ? node596 : 3'b010;
											assign node596 = (inp[1]) ? 3'b100 : 3'b010;
								assign node599 = (inp[5]) ? 3'b100 : node600;
									assign node600 = (inp[4]) ? 3'b100 : node601;
										assign node601 = (inp[1]) ? 3'b100 : 3'b010;
						assign node606 = (inp[8]) ? node626 : node607;
							assign node607 = (inp[3]) ? node615 : node608;
								assign node608 = (inp[4]) ? node610 : 3'b010;
									assign node610 = (inp[0]) ? 3'b100 : node611;
										assign node611 = (inp[5]) ? 3'b100 : 3'b010;
								assign node615 = (inp[0]) ? node617 : 3'b100;
									assign node617 = (inp[2]) ? node619 : 3'b100;
										assign node619 = (inp[5]) ? node621 : 3'b100;
											assign node621 = (inp[4]) ? node623 : 3'b100;
												assign node623 = (inp[1]) ? 3'b000 : 3'b100;
							assign node626 = (inp[3]) ? node634 : node627;
								assign node627 = (inp[4]) ? node629 : 3'b100;
									assign node629 = (inp[5]) ? node631 : 3'b100;
										assign node631 = (inp[0]) ? 3'b000 : 3'b100;
								assign node634 = (inp[2]) ? 3'b000 : node635;
									assign node635 = (inp[4]) ? 3'b000 : node636;
										assign node636 = (inp[0]) ? 3'b000 : node637;
											assign node637 = (inp[5]) ? 3'b000 : 3'b100;
					assign node643 = (inp[11]) ? 3'b000 : node644;
						assign node644 = (inp[8]) ? node658 : node645;
							assign node645 = (inp[3]) ? node655 : node646;
								assign node646 = (inp[4]) ? 3'b100 : node647;
									assign node647 = (inp[1]) ? 3'b100 : node648;
										assign node648 = (inp[0]) ? 3'b100 : node649;
											assign node649 = (inp[2]) ? 3'b100 : 3'b010;
								assign node655 = (inp[4]) ? 3'b000 : 3'b100;
							assign node658 = (inp[4]) ? 3'b000 : node659;
								assign node659 = (inp[3]) ? 3'b000 : node660;
									assign node660 = (inp[1]) ? node666 : node661;
										assign node661 = (inp[5]) ? node663 : 3'b100;
											assign node663 = (inp[0]) ? 3'b000 : 3'b100;
										assign node666 = (inp[0]) ? 3'b000 : node667;
											assign node667 = (inp[5]) ? 3'b000 : 3'b100;
			assign node674 = (inp[10]) ? 3'b000 : node675;
				assign node675 = (inp[7]) ? 3'b000 : node676;
					assign node676 = (inp[11]) ? node704 : node677;
						assign node677 = (inp[8]) ? node693 : node678;
							assign node678 = (inp[3]) ? 3'b100 : node679;
								assign node679 = (inp[4]) ? node681 : 3'b010;
									assign node681 = (inp[0]) ? node687 : node682;
										assign node682 = (inp[5]) ? node684 : 3'b010;
											assign node684 = (inp[2]) ? 3'b010 : 3'b100;
										assign node687 = (inp[1]) ? 3'b100 : node688;
											assign node688 = (inp[5]) ? 3'b100 : 3'b010;
							assign node693 = (inp[3]) ? node695 : 3'b100;
								assign node695 = (inp[0]) ? 3'b000 : node696;
									assign node696 = (inp[4]) ? 3'b000 : node697;
										assign node697 = (inp[2]) ? node699 : 3'b100;
											assign node699 = (inp[1]) ? 3'b000 : 3'b100;
						assign node704 = (inp[3]) ? 3'b000 : node705;
							assign node705 = (inp[8]) ? 3'b000 : node706;
								assign node706 = (inp[4]) ? node708 : 3'b100;
									assign node708 = (inp[5]) ? 3'b000 : node709;
										assign node709 = (inp[1]) ? 3'b000 : node710;
											assign node710 = (inp[2]) ? 3'b000 : 3'b100;

endmodule