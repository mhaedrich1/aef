module dtc_split75_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1080;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1142;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1169;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1190;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1204;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1224;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1234;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1270;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1293;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1371;
	wire [3-1:0] node1372;
	wire [3-1:0] node1374;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1384;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1391;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1400;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1441;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1448;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1456;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1470;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1481;
	wire [3-1:0] node1482;
	wire [3-1:0] node1484;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1493;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1513;
	wire [3-1:0] node1516;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;

	assign outp = (inp[3]) ? node872 : node1;
		assign node1 = (inp[4]) ? node385 : node2;
			assign node2 = (inp[9]) ? node158 : node3;
				assign node3 = (inp[7]) ? node103 : node4;
					assign node4 = (inp[0]) ? node66 : node5;
						assign node5 = (inp[6]) ? node35 : node6;
							assign node6 = (inp[1]) ? node22 : node7;
								assign node7 = (inp[11]) ? node15 : node8;
									assign node8 = (inp[8]) ? node12 : node9;
										assign node9 = (inp[10]) ? 3'b001 : 3'b101;
										assign node12 = (inp[5]) ? 3'b101 : 3'b001;
									assign node15 = (inp[10]) ? node19 : node16;
										assign node16 = (inp[5]) ? 3'b001 : 3'b001;
										assign node19 = (inp[5]) ? 3'b110 : 3'b001;
								assign node22 = (inp[5]) ? node30 : node23;
									assign node23 = (inp[11]) ? node27 : node24;
										assign node24 = (inp[2]) ? 3'b011 : 3'b001;
										assign node27 = (inp[10]) ? 3'b101 : 3'b111;
									assign node30 = (inp[8]) ? node32 : 3'b001;
										assign node32 = (inp[11]) ? 3'b001 : 3'b111;
							assign node35 = (inp[5]) ? node51 : node36;
								assign node36 = (inp[10]) ? node44 : node37;
									assign node37 = (inp[8]) ? node41 : node38;
										assign node38 = (inp[1]) ? 3'b101 : 3'b111;
										assign node41 = (inp[1]) ? 3'b101 : 3'b001;
									assign node44 = (inp[11]) ? node48 : node45;
										assign node45 = (inp[1]) ? 3'b011 : 3'b011;
										assign node48 = (inp[1]) ? 3'b111 : 3'b011;
								assign node51 = (inp[8]) ? node59 : node52;
									assign node52 = (inp[10]) ? node56 : node53;
										assign node53 = (inp[2]) ? 3'b011 : 3'b011;
										assign node56 = (inp[2]) ? 3'b011 : 3'b001;
									assign node59 = (inp[11]) ? node63 : node60;
										assign node60 = (inp[10]) ? 3'b111 : 3'b111;
										assign node63 = (inp[1]) ? 3'b011 : 3'b101;
						assign node66 = (inp[5]) ? node86 : node67;
							assign node67 = (inp[1]) ? node77 : node68;
								assign node68 = (inp[8]) ? node72 : node69;
									assign node69 = (inp[2]) ? 3'b111 : 3'b011;
									assign node72 = (inp[2]) ? node74 : 3'b111;
										assign node74 = (inp[11]) ? 3'b111 : 3'b011;
								assign node77 = (inp[6]) ? 3'b111 : node78;
									assign node78 = (inp[11]) ? node82 : node79;
										assign node79 = (inp[8]) ? 3'b111 : 3'b111;
										assign node82 = (inp[8]) ? 3'b111 : 3'b011;
							assign node86 = (inp[1]) ? node96 : node87;
								assign node87 = (inp[2]) ? node91 : node88;
									assign node88 = (inp[8]) ? 3'b101 : 3'b001;
									assign node91 = (inp[11]) ? 3'b101 : node92;
										assign node92 = (inp[8]) ? 3'b001 : 3'b101;
								assign node96 = (inp[6]) ? 3'b111 : node97;
									assign node97 = (inp[10]) ? 3'b011 : node98;
										assign node98 = (inp[2]) ? 3'b011 : 3'b011;
					assign node103 = (inp[5]) ? node125 : node104;
						assign node104 = (inp[0]) ? node114 : node105;
							assign node105 = (inp[11]) ? 3'b111 : node106;
								assign node106 = (inp[8]) ? node108 : 3'b111;
									assign node108 = (inp[2]) ? node110 : 3'b111;
										assign node110 = (inp[6]) ? 3'b101 : 3'b101;
							assign node114 = (inp[6]) ? 3'b111 : node115;
								assign node115 = (inp[1]) ? node117 : 3'b111;
									assign node117 = (inp[2]) ? node121 : node118;
										assign node118 = (inp[11]) ? 3'b111 : 3'b111;
										assign node121 = (inp[11]) ? 3'b111 : 3'b011;
						assign node125 = (inp[0]) ? node147 : node126;
							assign node126 = (inp[1]) ? node134 : node127;
								assign node127 = (inp[2]) ? 3'b111 : node128;
									assign node128 = (inp[8]) ? 3'b111 : node129;
										assign node129 = (inp[11]) ? 3'b101 : 3'b111;
								assign node134 = (inp[6]) ? node142 : node135;
									assign node135 = (inp[8]) ? node139 : node136;
										assign node136 = (inp[11]) ? 3'b101 : 3'b011;
										assign node139 = (inp[11]) ? 3'b011 : 3'b011;
									assign node142 = (inp[2]) ? 3'b111 : node143;
										assign node143 = (inp[11]) ? 3'b101 : 3'b111;
							assign node147 = (inp[1]) ? node149 : 3'b011;
								assign node149 = (inp[6]) ? 3'b111 : node150;
									assign node150 = (inp[2]) ? node154 : node151;
										assign node151 = (inp[8]) ? 3'b011 : 3'b011;
										assign node154 = (inp[11]) ? 3'b011 : 3'b111;
				assign node158 = (inp[6]) ? node278 : node159;
					assign node159 = (inp[0]) ? node219 : node160;
						assign node160 = (inp[10]) ? node190 : node161;
							assign node161 = (inp[7]) ? node177 : node162;
								assign node162 = (inp[5]) ? node170 : node163;
									assign node163 = (inp[1]) ? node167 : node164;
										assign node164 = (inp[8]) ? 3'b001 : 3'b110;
										assign node167 = (inp[8]) ? 3'b101 : 3'b001;
									assign node170 = (inp[11]) ? node174 : node171;
										assign node171 = (inp[1]) ? 3'b001 : 3'b110;
										assign node174 = (inp[1]) ? 3'b110 : 3'b010;
								assign node177 = (inp[5]) ? node185 : node178;
									assign node178 = (inp[11]) ? node182 : node179;
										assign node179 = (inp[1]) ? 3'b101 : 3'b101;
										assign node182 = (inp[1]) ? 3'b101 : 3'b001;
									assign node185 = (inp[8]) ? 3'b001 : node186;
										assign node186 = (inp[2]) ? 3'b001 : 3'b110;
							assign node190 = (inp[5]) ? node206 : node191;
								assign node191 = (inp[1]) ? node199 : node192;
									assign node192 = (inp[7]) ? node196 : node193;
										assign node193 = (inp[8]) ? 3'b110 : 3'b010;
										assign node196 = (inp[8]) ? 3'b000 : 3'b110;
									assign node199 = (inp[11]) ? node203 : node200;
										assign node200 = (inp[2]) ? 3'b001 : 3'b001;
										assign node203 = (inp[7]) ? 3'b000 : 3'b110;
								assign node206 = (inp[7]) ? node212 : node207;
									assign node207 = (inp[1]) ? 3'b010 : node208;
										assign node208 = (inp[2]) ? 3'b010 : 3'b100;
									assign node212 = (inp[11]) ? node216 : node213;
										assign node213 = (inp[1]) ? 3'b110 : 3'b110;
										assign node216 = (inp[1]) ? 3'b110 : 3'b010;
						assign node219 = (inp[1]) ? node249 : node220;
							assign node220 = (inp[10]) ? node234 : node221;
								assign node221 = (inp[11]) ? node229 : node222;
									assign node222 = (inp[5]) ? node226 : node223;
										assign node223 = (inp[7]) ? 3'b011 : 3'b000;
										assign node226 = (inp[7]) ? 3'b101 : 3'b001;
									assign node229 = (inp[5]) ? node231 : 3'b101;
										assign node231 = (inp[7]) ? 3'b101 : 3'b001;
								assign node234 = (inp[5]) ? node242 : node235;
									assign node235 = (inp[7]) ? node239 : node236;
										assign node236 = (inp[2]) ? 3'b001 : 3'b001;
										assign node239 = (inp[8]) ? 3'b101 : 3'b101;
									assign node242 = (inp[7]) ? node246 : node243;
										assign node243 = (inp[11]) ? 3'b110 : 3'b110;
										assign node246 = (inp[8]) ? 3'b001 : 3'b110;
							assign node249 = (inp[10]) ? node263 : node250;
								assign node250 = (inp[5]) ? node258 : node251;
									assign node251 = (inp[7]) ? node255 : node252;
										assign node252 = (inp[8]) ? 3'b011 : 3'b001;
										assign node255 = (inp[11]) ? 3'b011 : 3'b111;
									assign node258 = (inp[11]) ? 3'b101 : node259;
										assign node259 = (inp[7]) ? 3'b011 : 3'b101;
								assign node263 = (inp[5]) ? node271 : node264;
									assign node264 = (inp[2]) ? node268 : node265;
										assign node265 = (inp[11]) ? 3'b101 : 3'b101;
										assign node268 = (inp[7]) ? 3'b011 : 3'b101;
									assign node271 = (inp[7]) ? node275 : node272;
										assign node272 = (inp[11]) ? 3'b110 : 3'b001;
										assign node275 = (inp[11]) ? 3'b001 : 3'b101;
					assign node278 = (inp[0]) ? node334 : node279;
						assign node279 = (inp[7]) ? node305 : node280;
							assign node280 = (inp[5]) ? node294 : node281;
								assign node281 = (inp[10]) ? node287 : node282;
									assign node282 = (inp[1]) ? node284 : 3'b101;
										assign node284 = (inp[8]) ? 3'b011 : 3'b001;
									assign node287 = (inp[1]) ? node291 : node288;
										assign node288 = (inp[2]) ? 3'b001 : 3'b001;
										assign node291 = (inp[2]) ? 3'b101 : 3'b101;
								assign node294 = (inp[1]) ? node298 : node295;
									assign node295 = (inp[10]) ? 3'b110 : 3'b001;
									assign node298 = (inp[10]) ? node302 : node299;
										assign node299 = (inp[11]) ? 3'b101 : 3'b001;
										assign node302 = (inp[8]) ? 3'b001 : 3'b001;
							assign node305 = (inp[5]) ? node319 : node306;
								assign node306 = (inp[1]) ? node312 : node307;
									assign node307 = (inp[10]) ? 3'b101 : node308;
										assign node308 = (inp[11]) ? 3'b011 : 3'b011;
									assign node312 = (inp[10]) ? node316 : node313;
										assign node313 = (inp[8]) ? 3'b111 : 3'b111;
										assign node316 = (inp[8]) ? 3'b011 : 3'b011;
								assign node319 = (inp[10]) ? node327 : node320;
									assign node320 = (inp[1]) ? node324 : node321;
										assign node321 = (inp[11]) ? 3'b101 : 3'b101;
										assign node324 = (inp[11]) ? 3'b011 : 3'b011;
									assign node327 = (inp[1]) ? node331 : node328;
										assign node328 = (inp[2]) ? 3'b001 : 3'b001;
										assign node331 = (inp[11]) ? 3'b001 : 3'b101;
						assign node334 = (inp[7]) ? node364 : node335;
							assign node335 = (inp[5]) ? node349 : node336;
								assign node336 = (inp[11]) ? node344 : node337;
									assign node337 = (inp[1]) ? node341 : node338;
										assign node338 = (inp[10]) ? 3'b011 : 3'b111;
										assign node341 = (inp[2]) ? 3'b111 : 3'b111;
									assign node344 = (inp[8]) ? node346 : 3'b011;
										assign node346 = (inp[2]) ? 3'b111 : 3'b011;
								assign node349 = (inp[1]) ? node357 : node350;
									assign node350 = (inp[10]) ? node354 : node351;
										assign node351 = (inp[11]) ? 3'b101 : 3'b011;
										assign node354 = (inp[8]) ? 3'b101 : 3'b001;
									assign node357 = (inp[10]) ? node361 : node358;
										assign node358 = (inp[8]) ? 3'b111 : 3'b011;
										assign node361 = (inp[11]) ? 3'b101 : 3'b011;
							assign node364 = (inp[5]) ? node372 : node365;
								assign node365 = (inp[1]) ? 3'b111 : node366;
									assign node366 = (inp[10]) ? node368 : 3'b111;
										assign node368 = (inp[2]) ? 3'b111 : 3'b011;
								assign node372 = (inp[10]) ? node378 : node373;
									assign node373 = (inp[1]) ? 3'b111 : node374;
										assign node374 = (inp[8]) ? 3'b111 : 3'b011;
									assign node378 = (inp[1]) ? node382 : node379;
										assign node379 = (inp[2]) ? 3'b011 : 3'b001;
										assign node382 = (inp[8]) ? 3'b011 : 3'b011;
			assign node385 = (inp[0]) ? node625 : node386;
				assign node386 = (inp[9]) ? node512 : node387;
					assign node387 = (inp[11]) ? node451 : node388;
						assign node388 = (inp[1]) ? node420 : node389;
							assign node389 = (inp[7]) ? node405 : node390;
								assign node390 = (inp[6]) ? node398 : node391;
									assign node391 = (inp[10]) ? node395 : node392;
										assign node392 = (inp[5]) ? 3'b110 : 3'b001;
										assign node395 = (inp[5]) ? 3'b010 : 3'b110;
									assign node398 = (inp[10]) ? node402 : node399;
										assign node399 = (inp[8]) ? 3'b001 : 3'b101;
										assign node402 = (inp[5]) ? 3'b000 : 3'b101;
								assign node405 = (inp[5]) ? node413 : node406;
									assign node406 = (inp[2]) ? node410 : node407;
										assign node407 = (inp[10]) ? 3'b101 : 3'b001;
										assign node410 = (inp[8]) ? 3'b101 : 3'b001;
									assign node413 = (inp[2]) ? node417 : node414;
										assign node414 = (inp[8]) ? 3'b001 : 3'b101;
										assign node417 = (inp[8]) ? 3'b001 : 3'b001;
							assign node420 = (inp[8]) ? node436 : node421;
								assign node421 = (inp[5]) ? node429 : node422;
									assign node422 = (inp[7]) ? node426 : node423;
										assign node423 = (inp[10]) ? 3'b001 : 3'b001;
										assign node426 = (inp[6]) ? 3'b011 : 3'b000;
									assign node429 = (inp[10]) ? node433 : node430;
										assign node430 = (inp[7]) ? 3'b001 : 3'b010;
										assign node433 = (inp[6]) ? 3'b101 : 3'b110;
								assign node436 = (inp[6]) ? node444 : node437;
									assign node437 = (inp[5]) ? node441 : node438;
										assign node438 = (inp[7]) ? 3'b110 : 3'b101;
										assign node441 = (inp[10]) ? 3'b110 : 3'b011;
									assign node444 = (inp[7]) ? node448 : node445;
										assign node445 = (inp[10]) ? 3'b110 : 3'b010;
										assign node448 = (inp[2]) ? 3'b110 : 3'b111;
						assign node451 = (inp[6]) ? node481 : node452;
							assign node452 = (inp[1]) ? node466 : node453;
								assign node453 = (inp[7]) ? node461 : node454;
									assign node454 = (inp[10]) ? node458 : node455;
										assign node455 = (inp[5]) ? 3'b010 : 3'b010;
										assign node458 = (inp[5]) ? 3'b100 : 3'b010;
									assign node461 = (inp[5]) ? 3'b110 : node462;
										assign node462 = (inp[10]) ? 3'b110 : 3'b010;
								assign node466 = (inp[7]) ? node474 : node467;
									assign node467 = (inp[5]) ? node471 : node468;
										assign node468 = (inp[10]) ? 3'b110 : 3'b010;
										assign node471 = (inp[10]) ? 3'b010 : 3'b110;
									assign node474 = (inp[10]) ? node478 : node475;
										assign node475 = (inp[5]) ? 3'b000 : 3'b101;
										assign node478 = (inp[5]) ? 3'b110 : 3'b000;
							assign node481 = (inp[8]) ? node497 : node482;
								assign node482 = (inp[7]) ? node490 : node483;
									assign node483 = (inp[1]) ? node487 : node484;
										assign node484 = (inp[10]) ? 3'b000 : 3'b001;
										assign node487 = (inp[10]) ? 3'b110 : 3'b010;
									assign node490 = (inp[1]) ? node494 : node491;
										assign node491 = (inp[5]) ? 3'b010 : 3'b010;
										assign node494 = (inp[2]) ? 3'b001 : 3'b000;
								assign node497 = (inp[1]) ? node505 : node498;
									assign node498 = (inp[7]) ? node502 : node499;
										assign node499 = (inp[10]) ? 3'b010 : 3'b001;
										assign node502 = (inp[2]) ? 3'b010 : 3'b010;
									assign node505 = (inp[7]) ? node509 : node506;
										assign node506 = (inp[5]) ? 3'b010 : 3'b110;
										assign node509 = (inp[10]) ? 3'b001 : 3'b111;
					assign node512 = (inp[6]) ? node564 : node513;
						assign node513 = (inp[10]) ? node543 : node514;
							assign node514 = (inp[5]) ? node528 : node515;
								assign node515 = (inp[1]) ? node523 : node516;
									assign node516 = (inp[8]) ? node520 : node517;
										assign node517 = (inp[11]) ? 3'b100 : 3'b100;
										assign node520 = (inp[2]) ? 3'b010 : 3'b000;
									assign node523 = (inp[7]) ? node525 : 3'b010;
										assign node525 = (inp[8]) ? 3'b110 : 3'b010;
								assign node528 = (inp[7]) ? node536 : node529;
									assign node529 = (inp[1]) ? node533 : node530;
										assign node530 = (inp[2]) ? 3'b100 : 3'b000;
										assign node533 = (inp[11]) ? 3'b100 : 3'b100;
									assign node536 = (inp[2]) ? node540 : node537;
										assign node537 = (inp[1]) ? 3'b010 : 3'b100;
										assign node540 = (inp[1]) ? 3'b000 : 3'b010;
							assign node543 = (inp[5]) ? node557 : node544;
								assign node544 = (inp[7]) ? node550 : node545;
									assign node545 = (inp[8]) ? 3'b100 : node546;
										assign node546 = (inp[2]) ? 3'b100 : 3'b000;
									assign node550 = (inp[11]) ? node554 : node551;
										assign node551 = (inp[8]) ? 3'b010 : 3'b000;
										assign node554 = (inp[2]) ? 3'b000 : 3'b100;
								assign node557 = (inp[7]) ? node559 : 3'b000;
									assign node559 = (inp[1]) ? node561 : 3'b000;
										assign node561 = (inp[8]) ? 3'b100 : 3'b000;
						assign node564 = (inp[5]) ? node594 : node565;
							assign node565 = (inp[7]) ? node579 : node566;
								assign node566 = (inp[1]) ? node574 : node567;
									assign node567 = (inp[10]) ? node571 : node568;
										assign node568 = (inp[8]) ? 3'b110 : 3'b110;
										assign node571 = (inp[8]) ? 3'b010 : 3'b010;
									assign node574 = (inp[10]) ? 3'b110 : node575;
										assign node575 = (inp[8]) ? 3'b001 : 3'b111;
								assign node579 = (inp[10]) ? node587 : node580;
									assign node580 = (inp[8]) ? node584 : node581;
										assign node581 = (inp[1]) ? 3'b010 : 3'b001;
										assign node584 = (inp[1]) ? 3'b101 : 3'b001;
									assign node587 = (inp[1]) ? node591 : node588;
										assign node588 = (inp[2]) ? 3'b110 : 3'b110;
										assign node591 = (inp[11]) ? 3'b110 : 3'b001;
							assign node594 = (inp[11]) ? node610 : node595;
								assign node595 = (inp[8]) ? node603 : node596;
									assign node596 = (inp[2]) ? node600 : node597;
										assign node597 = (inp[10]) ? 3'b010 : 3'b110;
										assign node600 = (inp[7]) ? 3'b000 : 3'b010;
									assign node603 = (inp[10]) ? node607 : node604;
										assign node604 = (inp[7]) ? 3'b001 : 3'b000;
										assign node607 = (inp[7]) ? 3'b010 : 3'b010;
								assign node610 = (inp[7]) ? node618 : node611;
									assign node611 = (inp[10]) ? node615 : node612;
										assign node612 = (inp[8]) ? 3'b000 : 3'b110;
										assign node615 = (inp[1]) ? 3'b100 : 3'b100;
									assign node618 = (inp[10]) ? node622 : node619;
										assign node619 = (inp[1]) ? 3'b110 : 3'b110;
										assign node622 = (inp[1]) ? 3'b010 : 3'b000;
				assign node625 = (inp[9]) ? node751 : node626;
					assign node626 = (inp[7]) ? node688 : node627;
						assign node627 = (inp[1]) ? node659 : node628;
							assign node628 = (inp[5]) ? node644 : node629;
								assign node629 = (inp[8]) ? node637 : node630;
									assign node630 = (inp[11]) ? node634 : node631;
										assign node631 = (inp[6]) ? 3'b000 : 3'b001;
										assign node634 = (inp[2]) ? 3'b101 : 3'b111;
									assign node637 = (inp[2]) ? node641 : node638;
										assign node638 = (inp[11]) ? 3'b101 : 3'b100;
										assign node641 = (inp[10]) ? 3'b000 : 3'b100;
								assign node644 = (inp[10]) ? node652 : node645;
									assign node645 = (inp[6]) ? node649 : node646;
										assign node646 = (inp[8]) ? 3'b011 : 3'b011;
										assign node649 = (inp[11]) ? 3'b101 : 3'b011;
									assign node652 = (inp[6]) ? node656 : node653;
										assign node653 = (inp[2]) ? 3'b110 : 3'b110;
										assign node656 = (inp[11]) ? 3'b011 : 3'b111;
							assign node659 = (inp[6]) ? node675 : node660;
								assign node660 = (inp[5]) ? node668 : node661;
									assign node661 = (inp[11]) ? node665 : node662;
										assign node662 = (inp[10]) ? 3'b101 : 3'b101;
										assign node665 = (inp[8]) ? 3'b101 : 3'b001;
									assign node668 = (inp[11]) ? node672 : node669;
										assign node669 = (inp[2]) ? 3'b001 : 3'b000;
										assign node672 = (inp[10]) ? 3'b110 : 3'b100;
								assign node675 = (inp[5]) ? node683 : node676;
									assign node676 = (inp[8]) ? node680 : node677;
										assign node677 = (inp[2]) ? 3'b011 : 3'b101;
										assign node680 = (inp[2]) ? 3'b101 : 3'b011;
									assign node683 = (inp[2]) ? node685 : 3'b101;
										assign node685 = (inp[11]) ? 3'b101 : 3'b011;
						assign node688 = (inp[5]) ? node720 : node689;
							assign node689 = (inp[2]) ? node705 : node690;
								assign node690 = (inp[11]) ? node698 : node691;
									assign node691 = (inp[10]) ? node695 : node692;
										assign node692 = (inp[1]) ? 3'b101 : 3'b011;
										assign node695 = (inp[8]) ? 3'b111 : 3'b011;
									assign node698 = (inp[8]) ? node702 : node699;
										assign node699 = (inp[1]) ? 3'b101 : 3'b000;
										assign node702 = (inp[10]) ? 3'b111 : 3'b001;
								assign node705 = (inp[8]) ? node713 : node706;
									assign node706 = (inp[11]) ? node710 : node707;
										assign node707 = (inp[10]) ? 3'b011 : 3'b011;
										assign node710 = (inp[6]) ? 3'b111 : 3'b001;
									assign node713 = (inp[11]) ? node717 : node714;
										assign node714 = (inp[6]) ? 3'b001 : 3'b111;
										assign node717 = (inp[10]) ? 3'b111 : 3'b011;
							assign node720 = (inp[1]) ? node736 : node721;
								assign node721 = (inp[10]) ? node729 : node722;
									assign node722 = (inp[11]) ? node726 : node723;
										assign node723 = (inp[8]) ? 3'b101 : 3'b101;
										assign node726 = (inp[8]) ? 3'b101 : 3'b010;
									assign node729 = (inp[6]) ? node733 : node730;
										assign node730 = (inp[2]) ? 3'b001 : 3'b001;
										assign node733 = (inp[11]) ? 3'b100 : 3'b001;
								assign node736 = (inp[6]) ? node744 : node737;
									assign node737 = (inp[10]) ? node741 : node738;
										assign node738 = (inp[11]) ? 3'b111 : 3'b011;
										assign node741 = (inp[8]) ? 3'b101 : 3'b001;
									assign node744 = (inp[11]) ? node748 : node745;
										assign node745 = (inp[2]) ? 3'b111 : 3'b011;
										assign node748 = (inp[10]) ? 3'b011 : 3'b111;
					assign node751 = (inp[6]) ? node813 : node752;
						assign node752 = (inp[7]) ? node782 : node753;
							assign node753 = (inp[10]) ? node769 : node754;
								assign node754 = (inp[5]) ? node762 : node755;
									assign node755 = (inp[11]) ? node759 : node756;
										assign node756 = (inp[1]) ? 3'b001 : 3'b110;
										assign node759 = (inp[1]) ? 3'b110 : 3'b010;
									assign node762 = (inp[11]) ? node766 : node763;
										assign node763 = (inp[1]) ? 3'b110 : 3'b010;
										assign node766 = (inp[1]) ? 3'b010 : 3'b010;
								assign node769 = (inp[5]) ? node777 : node770;
									assign node770 = (inp[11]) ? node774 : node771;
										assign node771 = (inp[1]) ? 3'b110 : 3'b010;
										assign node774 = (inp[8]) ? 3'b010 : 3'b010;
									assign node777 = (inp[1]) ? node779 : 3'b100;
										assign node779 = (inp[8]) ? 3'b010 : 3'b100;
							assign node782 = (inp[1]) ? node798 : node783;
								assign node783 = (inp[5]) ? node791 : node784;
									assign node784 = (inp[10]) ? node788 : node785;
										assign node785 = (inp[8]) ? 3'b001 : 3'b001;
										assign node788 = (inp[11]) ? 3'b010 : 3'b110;
									assign node791 = (inp[10]) ? node795 : node792;
										assign node792 = (inp[2]) ? 3'b110 : 3'b110;
										assign node795 = (inp[8]) ? 3'b000 : 3'b100;
								assign node798 = (inp[5]) ? node806 : node799;
									assign node799 = (inp[10]) ? node803 : node800;
										assign node800 = (inp[8]) ? 3'b101 : 3'b001;
										assign node803 = (inp[11]) ? 3'b000 : 3'b001;
									assign node806 = (inp[10]) ? node810 : node807;
										assign node807 = (inp[2]) ? 3'b001 : 3'b000;
										assign node810 = (inp[8]) ? 3'b110 : 3'b010;
						assign node813 = (inp[10]) ? node843 : node814;
							assign node814 = (inp[5]) ? node828 : node815;
								assign node815 = (inp[1]) ? node823 : node816;
									assign node816 = (inp[11]) ? node820 : node817;
										assign node817 = (inp[7]) ? 3'b111 : 3'b101;
										assign node820 = (inp[7]) ? 3'b101 : 3'b011;
									assign node823 = (inp[7]) ? 3'b011 : node824;
										assign node824 = (inp[11]) ? 3'b101 : 3'b011;
								assign node828 = (inp[7]) ? node836 : node829;
									assign node829 = (inp[1]) ? node833 : node830;
										assign node830 = (inp[11]) ? 3'b111 : 3'b011;
										assign node833 = (inp[8]) ? 3'b001 : 3'b001;
									assign node836 = (inp[2]) ? node840 : node837;
										assign node837 = (inp[1]) ? 3'b001 : 3'b001;
										assign node840 = (inp[8]) ? 3'b101 : 3'b101;
							assign node843 = (inp[5]) ? node857 : node844;
								assign node844 = (inp[7]) ? node852 : node845;
									assign node845 = (inp[1]) ? node849 : node846;
										assign node846 = (inp[8]) ? 3'b001 : 3'b110;
										assign node849 = (inp[11]) ? 3'b001 : 3'b100;
									assign node852 = (inp[11]) ? node854 : 3'b101;
										assign node854 = (inp[1]) ? 3'b101 : 3'b001;
								assign node857 = (inp[7]) ? node865 : node858;
									assign node858 = (inp[1]) ? node862 : node859;
										assign node859 = (inp[2]) ? 3'b110 : 3'b010;
										assign node862 = (inp[11]) ? 3'b110 : 3'b111;
									assign node865 = (inp[1]) ? node869 : node866;
										assign node866 = (inp[11]) ? 3'b110 : 3'b000;
										assign node869 = (inp[8]) ? 3'b001 : 3'b000;
		assign node872 = (inp[4]) ? node1288 : node873;
			assign node873 = (inp[9]) ? node1105 : node874;
				assign node874 = (inp[6]) ? node982 : node875;
					assign node875 = (inp[0]) ? node927 : node876;
						assign node876 = (inp[7]) ? node902 : node877;
							assign node877 = (inp[5]) ? node893 : node878;
								assign node878 = (inp[11]) ? node886 : node879;
									assign node879 = (inp[8]) ? node883 : node880;
										assign node880 = (inp[1]) ? 3'b100 : 3'b100;
										assign node883 = (inp[2]) ? 3'b100 : 3'b000;
									assign node886 = (inp[10]) ? node890 : node887;
										assign node887 = (inp[1]) ? 3'b010 : 3'b000;
										assign node890 = (inp[1]) ? 3'b100 : 3'b000;
								assign node893 = (inp[10]) ? 3'b000 : node894;
									assign node894 = (inp[1]) ? node898 : node895;
										assign node895 = (inp[11]) ? 3'b000 : 3'b100;
										assign node898 = (inp[11]) ? 3'b100 : 3'b000;
							assign node902 = (inp[11]) ? node916 : node903;
								assign node903 = (inp[1]) ? node911 : node904;
									assign node904 = (inp[8]) ? node908 : node905;
										assign node905 = (inp[2]) ? 3'b100 : 3'b100;
										assign node908 = (inp[10]) ? 3'b000 : 3'b000;
									assign node911 = (inp[5]) ? 3'b110 : node912;
										assign node912 = (inp[8]) ? 3'b010 : 3'b110;
								assign node916 = (inp[1]) ? node922 : node917;
									assign node917 = (inp[10]) ? 3'b100 : node918;
										assign node918 = (inp[5]) ? 3'b100 : 3'b110;
									assign node922 = (inp[5]) ? 3'b000 : node923;
										assign node923 = (inp[2]) ? 3'b100 : 3'b100;
						assign node927 = (inp[7]) ? node951 : node928;
							assign node928 = (inp[1]) ? node942 : node929;
								assign node929 = (inp[10]) ? node935 : node930;
									assign node930 = (inp[5]) ? 3'b010 : node931;
										assign node931 = (inp[8]) ? 3'b110 : 3'b010;
									assign node935 = (inp[5]) ? node939 : node936;
										assign node936 = (inp[2]) ? 3'b010 : 3'b010;
										assign node939 = (inp[2]) ? 3'b100 : 3'b100;
								assign node942 = (inp[10]) ? node944 : 3'b110;
									assign node944 = (inp[5]) ? node948 : node945;
										assign node945 = (inp[11]) ? 3'b010 : 3'b110;
										assign node948 = (inp[2]) ? 3'b010 : 3'b100;
							assign node951 = (inp[1]) ? node967 : node952;
								assign node952 = (inp[11]) ? node960 : node953;
									assign node953 = (inp[10]) ? node957 : node954;
										assign node954 = (inp[8]) ? 3'b000 : 3'b010;
										assign node957 = (inp[2]) ? 3'b010 : 3'b010;
									assign node960 = (inp[2]) ? node964 : node961;
										assign node961 = (inp[8]) ? 3'b100 : 3'b010;
										assign node964 = (inp[10]) ? 3'b110 : 3'b100;
								assign node967 = (inp[5]) ? node975 : node968;
									assign node968 = (inp[8]) ? node972 : node969;
										assign node969 = (inp[2]) ? 3'b101 : 3'b101;
										assign node972 = (inp[10]) ? 3'b001 : 3'b011;
									assign node975 = (inp[10]) ? node979 : node976;
										assign node976 = (inp[2]) ? 3'b001 : 3'b100;
										assign node979 = (inp[8]) ? 3'b110 : 3'b010;
					assign node982 = (inp[0]) ? node1042 : node983;
						assign node983 = (inp[7]) ? node1011 : node984;
							assign node984 = (inp[1]) ? node998 : node985;
								assign node985 = (inp[10]) ? node993 : node986;
									assign node986 = (inp[11]) ? node990 : node987;
										assign node987 = (inp[2]) ? 3'b000 : 3'b000;
										assign node990 = (inp[5]) ? 3'b000 : 3'b100;
									assign node993 = (inp[2]) ? node995 : 3'b100;
										assign node995 = (inp[5]) ? 3'b100 : 3'b000;
								assign node998 = (inp[10]) ? node1004 : node999;
									assign node999 = (inp[5]) ? 3'b110 : node1000;
										assign node1000 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1004 = (inp[5]) ? node1008 : node1005;
										assign node1005 = (inp[11]) ? 3'b110 : 3'b110;
										assign node1008 = (inp[11]) ? 3'b010 : 3'b010;
							assign node1011 = (inp[10]) ? node1027 : node1012;
								assign node1012 = (inp[1]) ? node1020 : node1013;
									assign node1013 = (inp[5]) ? node1017 : node1014;
										assign node1014 = (inp[11]) ? 3'b101 : 3'b010;
										assign node1017 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1020 = (inp[11]) ? node1024 : node1021;
										assign node1021 = (inp[8]) ? 3'b111 : 3'b101;
										assign node1024 = (inp[5]) ? 3'b001 : 3'b101;
								assign node1027 = (inp[8]) ? node1035 : node1028;
									assign node1028 = (inp[1]) ? node1032 : node1029;
										assign node1029 = (inp[2]) ? 3'b110 : 3'b110;
										assign node1032 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1035 = (inp[11]) ? node1039 : node1036;
										assign node1036 = (inp[5]) ? 3'b010 : 3'b011;
										assign node1039 = (inp[1]) ? 3'b010 : 3'b110;
						assign node1042 = (inp[1]) ? node1074 : node1043;
							assign node1043 = (inp[7]) ? node1059 : node1044;
								assign node1044 = (inp[11]) ? node1052 : node1045;
									assign node1045 = (inp[5]) ? node1049 : node1046;
										assign node1046 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1049 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1052 = (inp[10]) ? node1056 : node1053;
										assign node1053 = (inp[5]) ? 3'b110 : 3'b011;
										assign node1056 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1059 = (inp[8]) ? node1067 : node1060;
									assign node1060 = (inp[10]) ? node1064 : node1061;
										assign node1061 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1064 = (inp[11]) ? 3'b110 : 3'b101;
									assign node1067 = (inp[5]) ? node1071 : node1068;
										assign node1068 = (inp[11]) ? 3'b001 : 3'b010;
										assign node1071 = (inp[11]) ? 3'b110 : 3'b101;
							assign node1074 = (inp[7]) ? node1090 : node1075;
								assign node1075 = (inp[10]) ? node1083 : node1076;
									assign node1076 = (inp[5]) ? node1080 : node1077;
										assign node1077 = (inp[8]) ? 3'b011 : 3'b101;
										assign node1080 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1083 = (inp[11]) ? node1087 : node1084;
										assign node1084 = (inp[5]) ? 3'b001 : 3'b000;
										assign node1087 = (inp[5]) ? 3'b110 : 3'b101;
								assign node1090 = (inp[5]) ? node1098 : node1091;
									assign node1091 = (inp[11]) ? node1095 : node1092;
										assign node1092 = (inp[8]) ? 3'b011 : 3'b111;
										assign node1095 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1098 = (inp[11]) ? node1102 : node1099;
										assign node1099 = (inp[10]) ? 3'b001 : 3'b011;
										assign node1102 = (inp[10]) ? 3'b001 : 3'b101;
				assign node1105 = (inp[6]) ? node1173 : node1106;
					assign node1106 = (inp[0]) ? node1120 : node1107;
						assign node1107 = (inp[1]) ? node1109 : 3'b000;
							assign node1109 = (inp[5]) ? 3'b000 : node1110;
								assign node1110 = (inp[10]) ? 3'b000 : node1111;
									assign node1111 = (inp[2]) ? node1115 : node1112;
										assign node1112 = (inp[7]) ? 3'b000 : 3'b000;
										assign node1115 = (inp[11]) ? 3'b100 : 3'b000;
						assign node1120 = (inp[10]) ? node1152 : node1121;
							assign node1121 = (inp[1]) ? node1137 : node1122;
								assign node1122 = (inp[5]) ? node1130 : node1123;
									assign node1123 = (inp[2]) ? node1127 : node1124;
										assign node1124 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1127 = (inp[8]) ? 3'b010 : 3'b100;
									assign node1130 = (inp[2]) ? node1134 : node1131;
										assign node1131 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1134 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1137 = (inp[7]) ? node1145 : node1138;
									assign node1138 = (inp[5]) ? node1142 : node1139;
										assign node1139 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1142 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1145 = (inp[5]) ? node1149 : node1146;
										assign node1146 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1149 = (inp[2]) ? 3'b010 : 3'b000;
							assign node1152 = (inp[5]) ? node1166 : node1153;
								assign node1153 = (inp[2]) ? node1159 : node1154;
									assign node1154 = (inp[7]) ? node1156 : 3'b000;
										assign node1156 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1159 = (inp[8]) ? node1163 : node1160;
										assign node1160 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1163 = (inp[11]) ? 3'b100 : 3'b100;
								assign node1166 = (inp[11]) ? 3'b000 : node1167;
									assign node1167 = (inp[7]) ? node1169 : 3'b000;
										assign node1169 = (inp[1]) ? 3'b100 : 3'b000;
					assign node1173 = (inp[0]) ? node1227 : node1174;
						assign node1174 = (inp[1]) ? node1198 : node1175;
							assign node1175 = (inp[7]) ? node1185 : node1176;
								assign node1176 = (inp[10]) ? 3'b000 : node1177;
									assign node1177 = (inp[5]) ? node1181 : node1178;
										assign node1178 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1181 = (inp[8]) ? 3'b000 : 3'b000;
								assign node1185 = (inp[10]) ? node1193 : node1186;
									assign node1186 = (inp[5]) ? node1190 : node1187;
										assign node1187 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1190 = (inp[11]) ? 3'b100 : 3'b100;
									assign node1193 = (inp[5]) ? 3'b000 : node1194;
										assign node1194 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1198 = (inp[10]) ? node1214 : node1199;
								assign node1199 = (inp[5]) ? node1207 : node1200;
									assign node1200 = (inp[2]) ? node1204 : node1201;
										assign node1201 = (inp[11]) ? 3'b010 : 3'b010;
										assign node1204 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1207 = (inp[7]) ? node1211 : node1208;
										assign node1208 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1211 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1214 = (inp[7]) ? node1220 : node1215;
									assign node1215 = (inp[5]) ? 3'b000 : node1216;
										assign node1216 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1220 = (inp[5]) ? node1224 : node1221;
										assign node1221 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1224 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1227 = (inp[5]) ? node1257 : node1228;
							assign node1228 = (inp[10]) ? node1244 : node1229;
								assign node1229 = (inp[11]) ? node1237 : node1230;
									assign node1230 = (inp[1]) ? node1234 : node1231;
										assign node1231 = (inp[7]) ? 3'b001 : 3'b110;
										assign node1234 = (inp[2]) ? 3'b001 : 3'b001;
									assign node1237 = (inp[7]) ? node1241 : node1238;
										assign node1238 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1241 = (inp[1]) ? 3'b001 : 3'b110;
								assign node1244 = (inp[11]) ? node1252 : node1245;
									assign node1245 = (inp[7]) ? node1249 : node1246;
										assign node1246 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1249 = (inp[8]) ? 3'b000 : 3'b110;
									assign node1252 = (inp[2]) ? node1254 : 3'b010;
										assign node1254 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1257 = (inp[10]) ? node1273 : node1258;
								assign node1258 = (inp[11]) ? node1266 : node1259;
									assign node1259 = (inp[7]) ? node1263 : node1260;
										assign node1260 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1263 = (inp[8]) ? 3'b110 : 3'b110;
									assign node1266 = (inp[1]) ? node1270 : node1267;
										assign node1267 = (inp[7]) ? 3'b010 : 3'b110;
										assign node1270 = (inp[7]) ? 3'b000 : 3'b010;
								assign node1273 = (inp[7]) ? node1281 : node1274;
									assign node1274 = (inp[11]) ? node1278 : node1275;
										assign node1275 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1278 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1281 = (inp[11]) ? node1285 : node1282;
										assign node1282 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1285 = (inp[1]) ? 3'b010 : 3'b100;
			assign node1288 = (inp[9]) ? node1464 : node1289;
				assign node1289 = (inp[6]) ? node1353 : node1290;
					assign node1290 = (inp[0]) ? node1308 : node1291;
						assign node1291 = (inp[1]) ? node1293 : 3'b000;
							assign node1293 = (inp[7]) ? node1295 : 3'b000;
								assign node1295 = (inp[5]) ? node1303 : node1296;
									assign node1296 = (inp[10]) ? node1300 : node1297;
										assign node1297 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1300 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1303 = (inp[11]) ? 3'b000 : node1304;
										assign node1304 = (inp[8]) ? 3'b000 : 3'b000;
						assign node1308 = (inp[1]) ? node1324 : node1309;
							assign node1309 = (inp[7]) ? node1311 : 3'b000;
								assign node1311 = (inp[5]) ? node1319 : node1312;
									assign node1312 = (inp[10]) ? node1316 : node1313;
										assign node1313 = (inp[11]) ? 3'b100 : 3'b001;
										assign node1316 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1319 = (inp[10]) ? 3'b000 : node1320;
										assign node1320 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1324 = (inp[7]) ? node1338 : node1325;
								assign node1325 = (inp[5]) ? node1333 : node1326;
									assign node1326 = (inp[10]) ? node1330 : node1327;
										assign node1327 = (inp[11]) ? 3'b100 : 3'b001;
										assign node1330 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1333 = (inp[10]) ? 3'b000 : node1334;
										assign node1334 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1338 = (inp[8]) ? node1346 : node1339;
									assign node1339 = (inp[5]) ? node1343 : node1340;
										assign node1340 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1343 = (inp[10]) ? 3'b000 : 3'b100;
									assign node1346 = (inp[5]) ? node1350 : node1347;
										assign node1347 = (inp[10]) ? 3'b010 : 3'b000;
										assign node1350 = (inp[10]) ? 3'b100 : 3'b010;
					assign node1353 = (inp[0]) ? node1405 : node1354;
						assign node1354 = (inp[7]) ? node1378 : node1355;
							assign node1355 = (inp[10]) ? node1371 : node1356;
								assign node1356 = (inp[8]) ? node1364 : node1357;
									assign node1357 = (inp[2]) ? node1361 : node1358;
										assign node1358 = (inp[5]) ? 3'b000 : 3'b000;
										assign node1361 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1364 = (inp[1]) ? node1368 : node1365;
										assign node1365 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1368 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1371 = (inp[5]) ? 3'b000 : node1372;
									assign node1372 = (inp[8]) ? node1374 : 3'b000;
										assign node1374 = (inp[1]) ? 3'b000 : 3'b100;
							assign node1378 = (inp[10]) ? node1394 : node1379;
								assign node1379 = (inp[1]) ? node1387 : node1380;
									assign node1380 = (inp[11]) ? node1384 : node1381;
										assign node1381 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1384 = (inp[5]) ? 3'b100 : 3'b110;
									assign node1387 = (inp[11]) ? node1391 : node1388;
										assign node1388 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1391 = (inp[5]) ? 3'b100 : 3'b010;
								assign node1394 = (inp[5]) ? node1400 : node1395;
									assign node1395 = (inp[11]) ? 3'b000 : node1396;
										assign node1396 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1400 = (inp[1]) ? node1402 : 3'b000;
										assign node1402 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1405 = (inp[7]) ? node1435 : node1406;
							assign node1406 = (inp[1]) ? node1422 : node1407;
								assign node1407 = (inp[8]) ? node1415 : node1408;
									assign node1408 = (inp[10]) ? node1412 : node1409;
										assign node1409 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1412 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1415 = (inp[5]) ? node1419 : node1416;
										assign node1416 = (inp[10]) ? 3'b010 : 3'b000;
										assign node1419 = (inp[10]) ? 3'b000 : 3'b010;
								assign node1422 = (inp[10]) ? node1428 : node1423;
									assign node1423 = (inp[11]) ? 3'b010 : node1424;
										assign node1424 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1428 = (inp[5]) ? node1432 : node1429;
										assign node1429 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1432 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1435 = (inp[10]) ? node1451 : node1436;
								assign node1436 = (inp[5]) ? node1444 : node1437;
									assign node1437 = (inp[8]) ? node1441 : node1438;
										assign node1438 = (inp[1]) ? 3'b001 : 3'b110;
										assign node1441 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1444 = (inp[8]) ? node1448 : node1445;
										assign node1445 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1448 = (inp[11]) ? 3'b110 : 3'b110;
								assign node1451 = (inp[11]) ? node1459 : node1452;
									assign node1452 = (inp[5]) ? node1456 : node1453;
										assign node1453 = (inp[8]) ? 3'b110 : 3'b110;
										assign node1456 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1459 = (inp[8]) ? 3'b010 : node1460;
										assign node1460 = (inp[5]) ? 3'b000 : 3'b010;
				assign node1464 = (inp[6]) ? node1478 : node1465;
					assign node1465 = (inp[7]) ? node1467 : 3'b000;
						assign node1467 = (inp[11]) ? 3'b000 : node1468;
							assign node1468 = (inp[0]) ? node1470 : 3'b000;
								assign node1470 = (inp[5]) ? 3'b000 : node1471;
									assign node1471 = (inp[10]) ? 3'b000 : node1472;
										assign node1472 = (inp[1]) ? 3'b100 : 3'b010;
					assign node1478 = (inp[0]) ? node1488 : node1479;
						assign node1479 = (inp[7]) ? node1481 : 3'b000;
							assign node1481 = (inp[5]) ? 3'b000 : node1482;
								assign node1482 = (inp[1]) ? node1484 : 3'b000;
									assign node1484 = (inp[10]) ? 3'b000 : 3'b100;
						assign node1488 = (inp[5]) ? node1516 : node1489;
							assign node1489 = (inp[1]) ? node1501 : node1490;
								assign node1490 = (inp[11]) ? node1496 : node1491;
									assign node1491 = (inp[7]) ? node1493 : 3'b000;
										assign node1493 = (inp[10]) ? 3'b000 : 3'b010;
									assign node1496 = (inp[10]) ? 3'b000 : node1497;
										assign node1497 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1501 = (inp[7]) ? node1509 : node1502;
									assign node1502 = (inp[10]) ? node1506 : node1503;
										assign node1503 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1506 = (inp[8]) ? 3'b000 : 3'b000;
									assign node1509 = (inp[10]) ? node1513 : node1510;
										assign node1510 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1513 = (inp[11]) ? 3'b100 : 3'b000;
							assign node1516 = (inp[10]) ? 3'b000 : node1517;
								assign node1517 = (inp[11]) ? 3'b000 : node1518;
									assign node1518 = (inp[7]) ? node1520 : 3'b000;
										assign node1520 = (inp[2]) ? 3'b100 : 3'b100;

endmodule