module dtc_split66_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node618;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node784;
	wire [3-1:0] node786;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node797;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node840;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node920;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node978;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node992;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1063;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1094;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;

	assign outp = (inp[6]) ? node362 : node1;
		assign node1 = (inp[9]) ? node321 : node2;
			assign node2 = (inp[0]) ? node242 : node3;
				assign node3 = (inp[7]) ? node99 : node4;
					assign node4 = (inp[10]) ? node70 : node5;
						assign node5 = (inp[1]) ? node45 : node6;
							assign node6 = (inp[11]) ? node28 : node7;
								assign node7 = (inp[8]) ? node13 : node8;
									assign node8 = (inp[3]) ? node10 : 3'b010;
										assign node10 = (inp[2]) ? 3'b100 : 3'b010;
									assign node13 = (inp[2]) ? node21 : node14;
										assign node14 = (inp[5]) ? 3'b110 : node15;
											assign node15 = (inp[3]) ? 3'b110 : node16;
												assign node16 = (inp[4]) ? 3'b110 : 3'b001;
										assign node21 = (inp[3]) ? node23 : 3'b110;
											assign node23 = (inp[5]) ? 3'b010 : node24;
												assign node24 = (inp[4]) ? 3'b010 : 3'b110;
								assign node28 = (inp[8]) ? node38 : node29;
									assign node29 = (inp[3]) ? node35 : node30;
										assign node30 = (inp[2]) ? 3'b100 : node31;
											assign node31 = (inp[4]) ? 3'b100 : 3'b010;
										assign node35 = (inp[2]) ? 3'b000 : 3'b100;
									assign node38 = (inp[4]) ? node40 : 3'b010;
										assign node40 = (inp[3]) ? node42 : 3'b010;
											assign node42 = (inp[2]) ? 3'b100 : 3'b010;
							assign node45 = (inp[8]) ? node55 : node46;
								assign node46 = (inp[11]) ? 3'b000 : node47;
									assign node47 = (inp[2]) ? node49 : 3'b100;
										assign node49 = (inp[4]) ? 3'b000 : node50;
											assign node50 = (inp[3]) ? 3'b000 : 3'b100;
								assign node55 = (inp[11]) ? node63 : node56;
									assign node56 = (inp[2]) ? node58 : 3'b010;
										assign node58 = (inp[3]) ? 3'b100 : node59;
											assign node59 = (inp[4]) ? 3'b100 : 3'b010;
									assign node63 = (inp[2]) ? node65 : 3'b100;
										assign node65 = (inp[3]) ? 3'b000 : node66;
											assign node66 = (inp[4]) ? 3'b000 : 3'b100;
						assign node70 = (inp[1]) ? 3'b000 : node71;
							assign node71 = (inp[8]) ? node81 : node72;
								assign node72 = (inp[2]) ? 3'b000 : node73;
									assign node73 = (inp[4]) ? 3'b000 : node74;
										assign node74 = (inp[5]) ? 3'b000 : node75;
											assign node75 = (inp[11]) ? 3'b000 : 3'b100;
								assign node81 = (inp[11]) ? node93 : node82;
									assign node82 = (inp[5]) ? node84 : 3'b100;
										assign node84 = (inp[2]) ? node88 : node85;
											assign node85 = (inp[3]) ? 3'b100 : 3'b010;
											assign node88 = (inp[3]) ? node90 : 3'b100;
												assign node90 = (inp[4]) ? 3'b000 : 3'b100;
									assign node93 = (inp[3]) ? 3'b000 : node94;
										assign node94 = (inp[2]) ? 3'b000 : 3'b100;
					assign node99 = (inp[10]) ? node167 : node100;
						assign node100 = (inp[1]) ? node138 : node101;
							assign node101 = (inp[8]) ? node123 : node102;
								assign node102 = (inp[11]) ? node114 : node103;
									assign node103 = (inp[5]) ? node111 : node104;
										assign node104 = (inp[2]) ? 3'b001 : node105;
											assign node105 = (inp[4]) ? 3'b001 : node106;
												assign node106 = (inp[3]) ? 3'b001 : 3'b101;
										assign node111 = (inp[2]) ? 3'b110 : 3'b001;
									assign node114 = (inp[2]) ? node118 : node115;
										assign node115 = (inp[3]) ? 3'b110 : 3'b001;
										assign node118 = (inp[3]) ? node120 : 3'b110;
											assign node120 = (inp[4]) ? 3'b010 : 3'b110;
								assign node123 = (inp[11]) ? node133 : node124;
									assign node124 = (inp[3]) ? 3'b101 : node125;
										assign node125 = (inp[5]) ? node127 : 3'b011;
											assign node127 = (inp[4]) ? 3'b101 : node128;
												assign node128 = (inp[2]) ? 3'b101 : 3'b011;
									assign node133 = (inp[3]) ? 3'b001 : node134;
										assign node134 = (inp[2]) ? 3'b001 : 3'b101;
							assign node138 = (inp[8]) ? node148 : node139;
								assign node139 = (inp[11]) ? node145 : node140;
									assign node140 = (inp[3]) ? node142 : 3'b110;
										assign node142 = (inp[2]) ? 3'b010 : 3'b110;
									assign node145 = (inp[3]) ? 3'b100 : 3'b010;
								assign node148 = (inp[11]) ? node158 : node149;
									assign node149 = (inp[3]) ? node155 : node150;
										assign node150 = (inp[4]) ? 3'b001 : node151;
											assign node151 = (inp[2]) ? 3'b001 : 3'b101;
										assign node155 = (inp[2]) ? 3'b110 : 3'b001;
									assign node158 = (inp[2]) ? node160 : 3'b110;
										assign node160 = (inp[3]) ? node162 : 3'b110;
											assign node162 = (inp[5]) ? 3'b010 : node163;
												assign node163 = (inp[4]) ? 3'b010 : 3'b110;
						assign node167 = (inp[1]) ? node205 : node168;
							assign node168 = (inp[8]) ? node194 : node169;
								assign node169 = (inp[11]) ? node185 : node170;
									assign node170 = (inp[3]) ? node178 : node171;
										assign node171 = (inp[2]) ? 3'b010 : node172;
											assign node172 = (inp[4]) ? node174 : 3'b110;
												assign node174 = (inp[5]) ? 3'b010 : 3'b110;
										assign node178 = (inp[5]) ? node180 : 3'b010;
											assign node180 = (inp[4]) ? node182 : 3'b010;
												assign node182 = (inp[2]) ? 3'b100 : 3'b010;
									assign node185 = (inp[4]) ? node187 : 3'b100;
										assign node187 = (inp[2]) ? node189 : 3'b010;
											assign node189 = (inp[5]) ? node191 : 3'b100;
												assign node191 = (inp[3]) ? 3'b000 : 3'b100;
								assign node194 = (inp[11]) ? node200 : node195;
									assign node195 = (inp[2]) ? 3'b110 : node196;
										assign node196 = (inp[3]) ? 3'b110 : 3'b001;
									assign node200 = (inp[2]) ? 3'b010 : node201;
										assign node201 = (inp[3]) ? 3'b010 : 3'b110;
							assign node205 = (inp[11]) ? node221 : node206;
								assign node206 = (inp[8]) ? node212 : node207;
									assign node207 = (inp[3]) ? node209 : 3'b100;
										assign node209 = (inp[4]) ? 3'b000 : 3'b100;
									assign node212 = (inp[2]) ? node214 : 3'b010;
										assign node214 = (inp[3]) ? node216 : 3'b010;
											assign node216 = (inp[5]) ? 3'b100 : node217;
												assign node217 = (inp[4]) ? 3'b100 : 3'b010;
								assign node221 = (inp[8]) ? node229 : node222;
									assign node222 = (inp[4]) ? 3'b000 : node223;
										assign node223 = (inp[2]) ? 3'b000 : node224;
											assign node224 = (inp[5]) ? 3'b000 : 3'b100;
									assign node229 = (inp[5]) ? node231 : 3'b100;
										assign node231 = (inp[4]) ? node237 : node232;
											assign node232 = (inp[3]) ? 3'b100 : node233;
												assign node233 = (inp[2]) ? 3'b100 : 3'b010;
											assign node237 = (inp[3]) ? node239 : 3'b100;
												assign node239 = (inp[2]) ? 3'b000 : 3'b100;
				assign node242 = (inp[7]) ? node258 : node243;
					assign node243 = (inp[1]) ? 3'b000 : node244;
						assign node244 = (inp[2]) ? 3'b000 : node245;
							assign node245 = (inp[10]) ? 3'b000 : node246;
								assign node246 = (inp[11]) ? 3'b000 : node247;
									assign node247 = (inp[8]) ? node249 : 3'b000;
										assign node249 = (inp[4]) ? node251 : 3'b100;
											assign node251 = (inp[3]) ? 3'b000 : 3'b100;
					assign node258 = (inp[10]) ? node310 : node259;
						assign node259 = (inp[1]) ? node289 : node260;
							assign node260 = (inp[8]) ? node274 : node261;
								assign node261 = (inp[11]) ? node269 : node262;
									assign node262 = (inp[2]) ? node264 : 3'b010;
										assign node264 = (inp[5]) ? 3'b100 : node265;
											assign node265 = (inp[4]) ? 3'b100 : 3'b010;
									assign node269 = (inp[2]) ? node271 : 3'b100;
										assign node271 = (inp[4]) ? 3'b000 : 3'b100;
								assign node274 = (inp[11]) ? node282 : node275;
									assign node275 = (inp[2]) ? node277 : 3'b110;
										assign node277 = (inp[4]) ? 3'b010 : node278;
											assign node278 = (inp[3]) ? 3'b010 : 3'b110;
									assign node282 = (inp[2]) ? node284 : 3'b010;
										assign node284 = (inp[4]) ? 3'b100 : node285;
											assign node285 = (inp[3]) ? 3'b100 : 3'b010;
							assign node289 = (inp[8]) ? node297 : node290;
								assign node290 = (inp[2]) ? 3'b000 : node291;
									assign node291 = (inp[11]) ? 3'b000 : node292;
										assign node292 = (inp[3]) ? 3'b000 : 3'b100;
								assign node297 = (inp[11]) ? node303 : node298;
									assign node298 = (inp[3]) ? 3'b100 : node299;
										assign node299 = (inp[2]) ? 3'b100 : 3'b010;
									assign node303 = (inp[2]) ? 3'b000 : node304;
										assign node304 = (inp[4]) ? node306 : 3'b100;
											assign node306 = (inp[3]) ? 3'b000 : 3'b100;
						assign node310 = (inp[11]) ? 3'b000 : node311;
							assign node311 = (inp[1]) ? 3'b000 : node312;
								assign node312 = (inp[8]) ? node314 : 3'b000;
									assign node314 = (inp[2]) ? node316 : 3'b100;
										assign node316 = (inp[3]) ? 3'b000 : 3'b100;
			assign node321 = (inp[0]) ? 3'b000 : node322;
				assign node322 = (inp[10]) ? 3'b000 : node323;
					assign node323 = (inp[7]) ? node325 : 3'b000;
						assign node325 = (inp[1]) ? node349 : node326;
							assign node326 = (inp[8]) ? node334 : node327;
								assign node327 = (inp[3]) ? 3'b000 : node328;
									assign node328 = (inp[11]) ? 3'b000 : node329;
										assign node329 = (inp[2]) ? 3'b000 : 3'b100;
								assign node334 = (inp[11]) ? node340 : node335;
									assign node335 = (inp[2]) ? 3'b100 : node336;
										assign node336 = (inp[4]) ? 3'b100 : 3'b010;
									assign node340 = (inp[2]) ? 3'b000 : node341;
										assign node341 = (inp[3]) ? node343 : 3'b100;
											assign node343 = (inp[5]) ? 3'b000 : node344;
												assign node344 = (inp[4]) ? 3'b000 : 3'b100;
							assign node349 = (inp[2]) ? 3'b000 : node350;
								assign node350 = (inp[4]) ? 3'b000 : node351;
									assign node351 = (inp[3]) ? 3'b000 : node352;
										assign node352 = (inp[11]) ? 3'b000 : node353;
											assign node353 = (inp[8]) ? 3'b100 : 3'b000;
		assign node362 = (inp[9]) ? node800 : node363;
			assign node363 = (inp[0]) ? node557 : node364;
				assign node364 = (inp[7]) ? node494 : node365;
					assign node365 = (inp[10]) ? node435 : node366;
						assign node366 = (inp[1]) ? node390 : node367;
							assign node367 = (inp[11]) ? node375 : node368;
								assign node368 = (inp[8]) ? 3'b111 : node369;
									assign node369 = (inp[3]) ? 3'b011 : node370;
										assign node370 = (inp[2]) ? 3'b011 : 3'b111;
								assign node375 = (inp[8]) ? node385 : node376;
									assign node376 = (inp[2]) ? 3'b101 : node377;
										assign node377 = (inp[3]) ? node379 : 3'b011;
											assign node379 = (inp[4]) ? 3'b101 : node380;
												assign node380 = (inp[5]) ? 3'b101 : 3'b011;
									assign node385 = (inp[2]) ? 3'b011 : node386;
										assign node386 = (inp[3]) ? 3'b011 : 3'b111;
							assign node390 = (inp[8]) ? node414 : node391;
								assign node391 = (inp[11]) ? node403 : node392;
									assign node392 = (inp[2]) ? node400 : node393;
										assign node393 = (inp[5]) ? 3'b101 : node394;
											assign node394 = (inp[3]) ? 3'b101 : node395;
												assign node395 = (inp[4]) ? 3'b101 : 3'b011;
										assign node400 = (inp[3]) ? 3'b001 : 3'b101;
									assign node403 = (inp[2]) ? node409 : node404;
										assign node404 = (inp[3]) ? 3'b001 : node405;
											assign node405 = (inp[4]) ? 3'b001 : 3'b101;
										assign node409 = (inp[4]) ? node411 : 3'b001;
											assign node411 = (inp[3]) ? 3'b110 : 3'b001;
								assign node414 = (inp[11]) ? node426 : node415;
									assign node415 = (inp[4]) ? node421 : node416;
										assign node416 = (inp[3]) ? 3'b011 : node417;
											assign node417 = (inp[5]) ? 3'b111 : 3'b011;
										assign node421 = (inp[3]) ? node423 : 3'b011;
											assign node423 = (inp[2]) ? 3'b101 : 3'b011;
									assign node426 = (inp[2]) ? node430 : node427;
										assign node427 = (inp[3]) ? 3'b101 : 3'b011;
										assign node430 = (inp[4]) ? node432 : 3'b101;
											assign node432 = (inp[3]) ? 3'b001 : 3'b101;
						assign node435 = (inp[1]) ? node457 : node436;
							assign node436 = (inp[8]) ? node448 : node437;
								assign node437 = (inp[11]) ? node443 : node438;
									assign node438 = (inp[2]) ? 3'b001 : node439;
										assign node439 = (inp[3]) ? 3'b001 : 3'b101;
									assign node443 = (inp[3]) ? 3'b110 : node444;
										assign node444 = (inp[2]) ? 3'b110 : 3'b001;
								assign node448 = (inp[11]) ? node450 : 3'b101;
									assign node450 = (inp[2]) ? 3'b001 : node451;
										assign node451 = (inp[4]) ? node453 : 3'b101;
											assign node453 = (inp[3]) ? 3'b001 : 3'b101;
							assign node457 = (inp[8]) ? node477 : node458;
								assign node458 = (inp[11]) ? node466 : node459;
									assign node459 = (inp[2]) ? node461 : 3'b110;
										assign node461 = (inp[4]) ? node463 : 3'b110;
											assign node463 = (inp[3]) ? 3'b010 : 3'b110;
									assign node466 = (inp[4]) ? node468 : 3'b010;
										assign node468 = (inp[2]) ? node474 : node469;
											assign node469 = (inp[5]) ? 3'b010 : node470;
												assign node470 = (inp[3]) ? 3'b010 : 3'b110;
											assign node474 = (inp[3]) ? 3'b100 : 3'b010;
								assign node477 = (inp[11]) ? node483 : node478;
									assign node478 = (inp[3]) ? 3'b001 : node479;
										assign node479 = (inp[2]) ? 3'b001 : 3'b101;
									assign node483 = (inp[3]) ? node487 : node484;
										assign node484 = (inp[2]) ? 3'b110 : 3'b001;
										assign node487 = (inp[2]) ? node489 : 3'b110;
											assign node489 = (inp[5]) ? node491 : 3'b110;
												assign node491 = (inp[4]) ? 3'b010 : 3'b110;
					assign node494 = (inp[10]) ? node512 : node495;
						assign node495 = (inp[8]) ? 3'b111 : node496;
							assign node496 = (inp[1]) ? node498 : 3'b111;
								assign node498 = (inp[11]) ? node506 : node499;
									assign node499 = (inp[2]) ? node501 : 3'b111;
										assign node501 = (inp[4]) ? node503 : 3'b111;
											assign node503 = (inp[3]) ? 3'b011 : 3'b111;
									assign node506 = (inp[3]) ? 3'b011 : node507;
										assign node507 = (inp[2]) ? 3'b011 : 3'b111;
						assign node512 = (inp[1]) ? node534 : node513;
							assign node513 = (inp[8]) ? node529 : node514;
								assign node514 = (inp[2]) ? node522 : node515;
									assign node515 = (inp[11]) ? 3'b011 : node516;
										assign node516 = (inp[5]) ? node518 : 3'b111;
											assign node518 = (inp[3]) ? 3'b011 : 3'b111;
									assign node522 = (inp[11]) ? node524 : 3'b011;
										assign node524 = (inp[4]) ? 3'b101 : node525;
											assign node525 = (inp[5]) ? 3'b101 : 3'b011;
								assign node529 = (inp[2]) ? node531 : 3'b111;
									assign node531 = (inp[11]) ? 3'b011 : 3'b111;
							assign node534 = (inp[8]) ? node546 : node535;
								assign node535 = (inp[11]) ? node541 : node536;
									assign node536 = (inp[3]) ? 3'b101 : node537;
										assign node537 = (inp[2]) ? 3'b101 : 3'b011;
									assign node541 = (inp[2]) ? 3'b001 : node542;
										assign node542 = (inp[3]) ? 3'b001 : 3'b101;
								assign node546 = (inp[11]) ? node552 : node547;
									assign node547 = (inp[2]) ? 3'b011 : node548;
										assign node548 = (inp[3]) ? 3'b011 : 3'b111;
									assign node552 = (inp[2]) ? 3'b101 : node553;
										assign node553 = (inp[3]) ? 3'b101 : 3'b011;
				assign node557 = (inp[7]) ? node667 : node558;
					assign node558 = (inp[10]) ? node602 : node559;
						assign node559 = (inp[1]) ? node583 : node560;
							assign node560 = (inp[8]) ? node572 : node561;
								assign node561 = (inp[2]) ? node565 : node562;
									assign node562 = (inp[11]) ? 3'b110 : 3'b001;
									assign node565 = (inp[11]) ? node567 : 3'b110;
										assign node567 = (inp[3]) ? 3'b010 : node568;
											assign node568 = (inp[4]) ? 3'b010 : 3'b110;
								assign node572 = (inp[11]) ? node578 : node573;
									assign node573 = (inp[2]) ? node575 : 3'b101;
										assign node575 = (inp[3]) ? 3'b001 : 3'b101;
									assign node578 = (inp[2]) ? node580 : 3'b001;
										assign node580 = (inp[3]) ? 3'b110 : 3'b001;
							assign node583 = (inp[11]) ? node593 : node584;
								assign node584 = (inp[2]) ? node590 : node585;
									assign node585 = (inp[8]) ? 3'b001 : node586;
										assign node586 = (inp[3]) ? 3'b010 : 3'b110;
									assign node590 = (inp[8]) ? 3'b110 : 3'b010;
								assign node593 = (inp[8]) ? node599 : node594;
									assign node594 = (inp[2]) ? 3'b100 : node595;
										assign node595 = (inp[5]) ? 3'b100 : 3'b010;
									assign node599 = (inp[2]) ? 3'b010 : 3'b110;
						assign node602 = (inp[1]) ? node640 : node603;
							assign node603 = (inp[8]) ? node623 : node604;
								assign node604 = (inp[2]) ? node608 : node605;
									assign node605 = (inp[11]) ? 3'b100 : 3'b010;
									assign node608 = (inp[5]) ? node618 : node609;
										assign node609 = (inp[4]) ? 3'b100 : node610;
											assign node610 = (inp[3]) ? node614 : node611;
												assign node611 = (inp[11]) ? 3'b100 : 3'b010;
												assign node614 = (inp[11]) ? 3'b000 : 3'b100;
										assign node618 = (inp[3]) ? node620 : 3'b100;
											assign node620 = (inp[11]) ? 3'b000 : 3'b100;
								assign node623 = (inp[11]) ? node629 : node624;
									assign node624 = (inp[3]) ? node626 : 3'b110;
										assign node626 = (inp[2]) ? 3'b010 : 3'b110;
									assign node629 = (inp[2]) ? node637 : node630;
										assign node630 = (inp[3]) ? 3'b010 : node631;
											assign node631 = (inp[5]) ? 3'b010 : node632;
												assign node632 = (inp[4]) ? 3'b010 : 3'b110;
										assign node637 = (inp[3]) ? 3'b100 : 3'b010;
							assign node640 = (inp[8]) ? node656 : node641;
								assign node641 = (inp[11]) ? 3'b000 : node642;
									assign node642 = (inp[2]) ? node648 : node643;
										assign node643 = (inp[5]) ? node645 : 3'b100;
											assign node645 = (inp[4]) ? 3'b000 : 3'b100;
										assign node648 = (inp[4]) ? 3'b000 : node649;
											assign node649 = (inp[5]) ? 3'b000 : node650;
												assign node650 = (inp[3]) ? 3'b000 : 3'b100;
								assign node656 = (inp[11]) ? node660 : node657;
									assign node657 = (inp[2]) ? 3'b100 : 3'b010;
									assign node660 = (inp[2]) ? node662 : 3'b100;
										assign node662 = (inp[3]) ? 3'b000 : node663;
											assign node663 = (inp[4]) ? 3'b000 : 3'b100;
					assign node667 = (inp[10]) ? node731 : node668;
						assign node668 = (inp[1]) ? node710 : node669;
							assign node669 = (inp[8]) ? node693 : node670;
								assign node670 = (inp[11]) ? node682 : node671;
									assign node671 = (inp[2]) ? node679 : node672;
										assign node672 = (inp[3]) ? 3'b011 : node673;
											assign node673 = (inp[5]) ? 3'b011 : node674;
												assign node674 = (inp[4]) ? 3'b011 : 3'b111;
										assign node679 = (inp[3]) ? 3'b101 : 3'b011;
									assign node682 = (inp[4]) ? node688 : node683;
										assign node683 = (inp[2]) ? 3'b101 : node684;
											assign node684 = (inp[5]) ? 3'b101 : 3'b011;
										assign node688 = (inp[5]) ? node690 : 3'b101;
											assign node690 = (inp[2]) ? 3'b001 : 3'b101;
								assign node693 = (inp[11]) ? node699 : node694;
									assign node694 = (inp[2]) ? node696 : 3'b111;
										assign node696 = (inp[3]) ? 3'b011 : 3'b111;
									assign node699 = (inp[2]) ? node705 : node700;
										assign node700 = (inp[4]) ? 3'b011 : node701;
											assign node701 = (inp[3]) ? 3'b011 : 3'b111;
										assign node705 = (inp[4]) ? node707 : 3'b011;
											assign node707 = (inp[3]) ? 3'b101 : 3'b011;
							assign node710 = (inp[8]) ? node722 : node711;
								assign node711 = (inp[2]) ? node715 : node712;
									assign node712 = (inp[11]) ? 3'b001 : 3'b101;
									assign node715 = (inp[11]) ? node717 : 3'b001;
										assign node717 = (inp[3]) ? 3'b110 : node718;
											assign node718 = (inp[4]) ? 3'b110 : 3'b001;
								assign node722 = (inp[2]) ? node726 : node723;
									assign node723 = (inp[11]) ? 3'b101 : 3'b011;
									assign node726 = (inp[11]) ? node728 : 3'b101;
										assign node728 = (inp[3]) ? 3'b001 : 3'b101;
						assign node731 = (inp[1]) ? node775 : node732;
							assign node732 = (inp[8]) ? node750 : node733;
								assign node733 = (inp[11]) ? node743 : node734;
									assign node734 = (inp[2]) ? node736 : 3'b001;
										assign node736 = (inp[3]) ? node738 : 3'b001;
											assign node738 = (inp[5]) ? 3'b110 : node739;
												assign node739 = (inp[4]) ? 3'b110 : 3'b001;
									assign node743 = (inp[3]) ? node747 : node744;
										assign node744 = (inp[2]) ? 3'b110 : 3'b001;
										assign node747 = (inp[2]) ? 3'b010 : 3'b110;
								assign node750 = (inp[11]) ? node762 : node751;
									assign node751 = (inp[3]) ? node757 : node752;
										assign node752 = (inp[4]) ? 3'b101 : node753;
											assign node753 = (inp[2]) ? 3'b101 : 3'b011;
										assign node757 = (inp[4]) ? node759 : 3'b101;
											assign node759 = (inp[2]) ? 3'b001 : 3'b101;
									assign node762 = (inp[5]) ? node768 : node763;
										assign node763 = (inp[3]) ? 3'b001 : node764;
											assign node764 = (inp[2]) ? 3'b001 : 3'b101;
										assign node768 = (inp[2]) ? node770 : 3'b101;
											assign node770 = (inp[3]) ? node772 : 3'b001;
												assign node772 = (inp[4]) ? 3'b110 : 3'b001;
							assign node775 = (inp[8]) ? node789 : node776;
								assign node776 = (inp[11]) ? node784 : node777;
									assign node777 = (inp[2]) ? node779 : 3'b110;
										assign node779 = (inp[4]) ? 3'b010 : node780;
											assign node780 = (inp[3]) ? 3'b010 : 3'b110;
									assign node784 = (inp[2]) ? node786 : 3'b010;
										assign node786 = (inp[5]) ? 3'b100 : 3'b010;
								assign node789 = (inp[11]) ? node795 : node790;
									assign node790 = (inp[3]) ? node792 : 3'b001;
										assign node792 = (inp[2]) ? 3'b110 : 3'b001;
									assign node795 = (inp[3]) ? node797 : 3'b110;
										assign node797 = (inp[2]) ? 3'b010 : 3'b110;
			assign node800 = (inp[0]) ? node1020 : node801;
				assign node801 = (inp[7]) ? node901 : node802;
					assign node802 = (inp[10]) ? node862 : node803;
						assign node803 = (inp[8]) ? node835 : node804;
							assign node804 = (inp[1]) ? node816 : node805;
								assign node805 = (inp[11]) ? node809 : node806;
									assign node806 = (inp[3]) ? 3'b010 : 3'b110;
									assign node809 = (inp[2]) ? 3'b100 : node810;
										assign node810 = (inp[4]) ? node812 : 3'b010;
											assign node812 = (inp[3]) ? 3'b100 : 3'b010;
								assign node816 = (inp[11]) ? node828 : node817;
									assign node817 = (inp[5]) ? node823 : node818;
										assign node818 = (inp[2]) ? 3'b100 : node819;
											assign node819 = (inp[3]) ? 3'b100 : 3'b010;
										assign node823 = (inp[2]) ? node825 : 3'b100;
											assign node825 = (inp[3]) ? 3'b000 : 3'b100;
									assign node828 = (inp[3]) ? 3'b000 : node829;
										assign node829 = (inp[4]) ? 3'b000 : node830;
											assign node830 = (inp[2]) ? 3'b000 : 3'b100;
							assign node835 = (inp[11]) ? node849 : node836;
								assign node836 = (inp[1]) ? node844 : node837;
									assign node837 = (inp[2]) ? 3'b110 : node838;
										assign node838 = (inp[4]) ? node840 : 3'b001;
											assign node840 = (inp[3]) ? 3'b110 : 3'b001;
									assign node844 = (inp[3]) ? 3'b010 : node845;
										assign node845 = (inp[2]) ? 3'b010 : 3'b110;
								assign node849 = (inp[1]) ? node857 : node850;
									assign node850 = (inp[2]) ? 3'b010 : node851;
										assign node851 = (inp[4]) ? node853 : 3'b110;
											assign node853 = (inp[3]) ? 3'b010 : 3'b110;
									assign node857 = (inp[3]) ? 3'b100 : node858;
										assign node858 = (inp[2]) ? 3'b100 : 3'b010;
						assign node862 = (inp[1]) ? node888 : node863;
							assign node863 = (inp[2]) ? node875 : node864;
								assign node864 = (inp[8]) ? node872 : node865;
									assign node865 = (inp[11]) ? 3'b000 : node866;
										assign node866 = (inp[3]) ? node868 : 3'b100;
											assign node868 = (inp[4]) ? 3'b000 : 3'b100;
									assign node872 = (inp[11]) ? 3'b100 : 3'b010;
								assign node875 = (inp[8]) ? node877 : 3'b000;
									assign node877 = (inp[11]) ? node881 : node878;
										assign node878 = (inp[3]) ? 3'b100 : 3'b010;
										assign node881 = (inp[5]) ? 3'b000 : node882;
											assign node882 = (inp[3]) ? 3'b000 : node883;
												assign node883 = (inp[4]) ? 3'b000 : 3'b100;
							assign node888 = (inp[8]) ? node890 : 3'b000;
								assign node890 = (inp[2]) ? 3'b000 : node891;
									assign node891 = (inp[11]) ? 3'b000 : node892;
										assign node892 = (inp[3]) ? node894 : 3'b100;
											assign node894 = (inp[5]) ? 3'b000 : node895;
												assign node895 = (inp[4]) ? 3'b000 : 3'b100;
					assign node901 = (inp[10]) ? node965 : node902;
						assign node902 = (inp[1]) ? node938 : node903;
							assign node903 = (inp[11]) ? node927 : node904;
								assign node904 = (inp[8]) ? node920 : node905;
									assign node905 = (inp[2]) ? node913 : node906;
										assign node906 = (inp[3]) ? node908 : 3'b101;
											assign node908 = (inp[4]) ? node910 : 3'b101;
												assign node910 = (inp[5]) ? 3'b001 : 3'b101;
										assign node913 = (inp[3]) ? 3'b001 : node914;
											assign node914 = (inp[4]) ? 3'b001 : node915;
												assign node915 = (inp[5]) ? 3'b001 : 3'b101;
									assign node920 = (inp[2]) ? node922 : 3'b011;
										assign node922 = (inp[5]) ? 3'b101 : node923;
											assign node923 = (inp[3]) ? 3'b101 : 3'b011;
								assign node927 = (inp[8]) ? node931 : node928;
									assign node928 = (inp[2]) ? 3'b110 : 3'b001;
									assign node931 = (inp[2]) ? node933 : 3'b101;
										assign node933 = (inp[3]) ? 3'b001 : node934;
											assign node934 = (inp[4]) ? 3'b001 : 3'b101;
							assign node938 = (inp[8]) ? node954 : node939;
								assign node939 = (inp[2]) ? node951 : node940;
									assign node940 = (inp[11]) ? node948 : node941;
										assign node941 = (inp[3]) ? node943 : 3'b001;
											assign node943 = (inp[4]) ? 3'b110 : node944;
												assign node944 = (inp[5]) ? 3'b110 : 3'b001;
										assign node948 = (inp[3]) ? 3'b010 : 3'b110;
									assign node951 = (inp[11]) ? 3'b010 : 3'b110;
								assign node954 = (inp[11]) ? node962 : node955;
									assign node955 = (inp[2]) ? 3'b001 : node956;
										assign node956 = (inp[4]) ? node958 : 3'b101;
											assign node958 = (inp[3]) ? 3'b001 : 3'b101;
									assign node962 = (inp[2]) ? 3'b110 : 3'b001;
						assign node965 = (inp[1]) ? node999 : node966;
							assign node966 = (inp[11]) ? node982 : node967;
								assign node967 = (inp[8]) ? node973 : node968;
									assign node968 = (inp[2]) ? node970 : 3'b110;
										assign node970 = (inp[3]) ? 3'b010 : 3'b110;
									assign node973 = (inp[2]) ? node975 : 3'b001;
										assign node975 = (inp[3]) ? 3'b110 : node976;
											assign node976 = (inp[5]) ? node978 : 3'b001;
												assign node978 = (inp[4]) ? 3'b110 : 3'b001;
								assign node982 = (inp[4]) ? node988 : node983;
									assign node983 = (inp[8]) ? node985 : 3'b010;
										assign node985 = (inp[2]) ? 3'b010 : 3'b110;
									assign node988 = (inp[8]) ? node992 : node989;
										assign node989 = (inp[2]) ? 3'b100 : 3'b010;
										assign node992 = (inp[2]) ? node994 : 3'b110;
											assign node994 = (inp[3]) ? 3'b010 : node995;
												assign node995 = (inp[5]) ? 3'b010 : 3'b110;
							assign node999 = (inp[8]) ? node1013 : node1000;
								assign node1000 = (inp[11]) ? node1006 : node1001;
									assign node1001 = (inp[4]) ? 3'b100 : node1002;
										assign node1002 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1006 = (inp[2]) ? 3'b000 : node1007;
										assign node1007 = (inp[4]) ? node1009 : 3'b100;
											assign node1009 = (inp[3]) ? 3'b000 : 3'b100;
								assign node1013 = (inp[2]) ? node1017 : node1014;
									assign node1014 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1017 = (inp[11]) ? 3'b100 : 3'b010;
				assign node1020 = (inp[7]) ? node1046 : node1021;
					assign node1021 = (inp[10]) ? 3'b000 : node1022;
						assign node1022 = (inp[8]) ? node1024 : 3'b000;
							assign node1024 = (inp[1]) ? 3'b000 : node1025;
								assign node1025 = (inp[11]) ? node1037 : node1026;
									assign node1026 = (inp[3]) ? node1034 : node1027;
										assign node1027 = (inp[5]) ? 3'b100 : node1028;
											assign node1028 = (inp[2]) ? 3'b100 : node1029;
												assign node1029 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1034 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1037 = (inp[2]) ? 3'b000 : node1038;
										assign node1038 = (inp[4]) ? 3'b000 : node1039;
											assign node1039 = (inp[3]) ? 3'b000 : 3'b100;
					assign node1046 = (inp[10]) ? node1110 : node1047;
						assign node1047 = (inp[1]) ? node1087 : node1048;
							assign node1048 = (inp[8]) ? node1066 : node1049;
								assign node1049 = (inp[11]) ? node1059 : node1050;
									assign node1050 = (inp[2]) ? node1056 : node1051;
										assign node1051 = (inp[4]) ? 3'b010 : node1052;
											assign node1052 = (inp[3]) ? 3'b010 : 3'b110;
										assign node1056 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1059 = (inp[4]) ? node1061 : 3'b100;
										assign node1061 = (inp[2]) ? node1063 : 3'b100;
											assign node1063 = (inp[3]) ? 3'b000 : 3'b100;
								assign node1066 = (inp[11]) ? node1074 : node1067;
									assign node1067 = (inp[2]) ? 3'b110 : node1068;
										assign node1068 = (inp[5]) ? 3'b110 : node1069;
											assign node1069 = (inp[3]) ? 3'b110 : 3'b001;
									assign node1074 = (inp[2]) ? node1080 : node1075;
										assign node1075 = (inp[3]) ? 3'b010 : node1076;
											assign node1076 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1080 = (inp[5]) ? node1082 : 3'b010;
											assign node1082 = (inp[4]) ? node1084 : 3'b010;
												assign node1084 = (inp[3]) ? 3'b100 : 3'b010;
							assign node1087 = (inp[11]) ? node1103 : node1088;
								assign node1088 = (inp[8]) ? node1098 : node1089;
									assign node1089 = (inp[2]) ? node1091 : 3'b100;
										assign node1091 = (inp[3]) ? 3'b000 : node1092;
											assign node1092 = (inp[5]) ? node1094 : 3'b100;
												assign node1094 = (inp[4]) ? 3'b000 : 3'b100;
									assign node1098 = (inp[3]) ? node1100 : 3'b010;
										assign node1100 = (inp[2]) ? 3'b100 : 3'b010;
								assign node1103 = (inp[8]) ? node1105 : 3'b000;
									assign node1105 = (inp[2]) ? node1107 : 3'b100;
										assign node1107 = (inp[3]) ? 3'b000 : 3'b100;
						assign node1110 = (inp[1]) ? node1132 : node1111;
							assign node1111 = (inp[8]) ? node1121 : node1112;
								assign node1112 = (inp[11]) ? 3'b000 : node1113;
									assign node1113 = (inp[4]) ? 3'b000 : node1114;
										assign node1114 = (inp[3]) ? 3'b000 : node1115;
											assign node1115 = (inp[2]) ? 3'b000 : 3'b100;
								assign node1121 = (inp[11]) ? node1127 : node1122;
									assign node1122 = (inp[3]) ? 3'b100 : node1123;
										assign node1123 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1127 = (inp[2]) ? 3'b000 : node1128;
										assign node1128 = (inp[3]) ? 3'b000 : 3'b100;
							assign node1132 = (inp[3]) ? 3'b000 : node1133;
								assign node1133 = (inp[2]) ? 3'b000 : node1134;
									assign node1134 = (inp[5]) ? 3'b000 : node1135;
										assign node1135 = (inp[8]) ? node1137 : 3'b000;
											assign node1137 = (inp[11]) ? 3'b000 : 3'b100;

endmodule