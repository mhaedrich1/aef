module dtc_split25_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node13;
	wire [1-1:0] node17;
	wire [1-1:0] node18;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node23;
	wire [1-1:0] node25;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node37;
	wire [1-1:0] node38;
	wire [1-1:0] node40;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node44;
	wire [1-1:0] node49;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node63;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node77;
	wire [1-1:0] node80;
	wire [1-1:0] node83;
	wire [1-1:0] node84;
	wire [1-1:0] node86;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node98;
	wire [1-1:0] node99;
	wire [1-1:0] node100;
	wire [1-1:0] node102;
	wire [1-1:0] node104;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node118;
	wire [1-1:0] node120;
	wire [1-1:0] node123;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node135;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node142;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node147;
	wire [1-1:0] node149;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node156;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node169;
	wire [1-1:0] node172;
	wire [1-1:0] node173;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node184;
	wire [1-1:0] node186;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node196;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node205;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node211;
	wire [1-1:0] node212;
	wire [1-1:0] node216;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node227;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node249;
	wire [1-1:0] node250;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node273;
	wire [1-1:0] node275;
	wire [1-1:0] node278;
	wire [1-1:0] node281;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node285;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node290;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node307;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node312;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node317;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node328;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node335;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node342;
	wire [1-1:0] node344;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node372;
	wire [1-1:0] node373;
	wire [1-1:0] node375;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node383;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node401;
	wire [1-1:0] node403;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node426;
	wire [1-1:0] node427;
	wire [1-1:0] node429;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node443;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node454;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node461;
	wire [1-1:0] node463;
	wire [1-1:0] node465;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node471;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node483;
	wire [1-1:0] node485;
	wire [1-1:0] node487;
	wire [1-1:0] node490;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node501;
	wire [1-1:0] node502;
	wire [1-1:0] node504;
	wire [1-1:0] node507;
	wire [1-1:0] node508;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node514;
	wire [1-1:0] node516;
	wire [1-1:0] node517;
	wire [1-1:0] node519;
	wire [1-1:0] node521;
	wire [1-1:0] node524;
	wire [1-1:0] node525;
	wire [1-1:0] node529;
	wire [1-1:0] node530;
	wire [1-1:0] node531;
	wire [1-1:0] node533;
	wire [1-1:0] node535;
	wire [1-1:0] node538;
	wire [1-1:0] node539;
	wire [1-1:0] node541;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node548;
	wire [1-1:0] node549;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node558;
	wire [1-1:0] node559;
	wire [1-1:0] node561;
	wire [1-1:0] node564;
	wire [1-1:0] node567;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node570;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node580;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node592;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node599;
	wire [1-1:0] node600;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node605;
	wire [1-1:0] node608;
	wire [1-1:0] node609;
	wire [1-1:0] node613;
	wire [1-1:0] node614;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node619;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node628;
	wire [1-1:0] node631;
	wire [1-1:0] node632;
	wire [1-1:0] node633;
	wire [1-1:0] node635;
	wire [1-1:0] node639;
	wire [1-1:0] node640;
	wire [1-1:0] node641;
	wire [1-1:0] node646;
	wire [1-1:0] node647;
	wire [1-1:0] node648;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node657;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node661;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node668;
	wire [1-1:0] node671;
	wire [1-1:0] node672;
	wire [1-1:0] node673;
	wire [1-1:0] node675;
	wire [1-1:0] node680;
	wire [1-1:0] node681;
	wire [1-1:0] node682;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node691;
	wire [1-1:0] node692;
	wire [1-1:0] node693;
	wire [1-1:0] node694;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node702;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node714;
	wire [1-1:0] node716;
	wire [1-1:0] node718;
	wire [1-1:0] node719;
	wire [1-1:0] node721;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node728;
	wire [1-1:0] node729;
	wire [1-1:0] node731;
	wire [1-1:0] node735;
	wire [1-1:0] node736;
	wire [1-1:0] node738;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node744;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node754;
	wire [1-1:0] node755;
	wire [1-1:0] node757;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node764;
	wire [1-1:0] node767;
	wire [1-1:0] node768;
	wire [1-1:0] node772;
	wire [1-1:0] node773;
	wire [1-1:0] node774;
	wire [1-1:0] node775;
	wire [1-1:0] node777;
	wire [1-1:0] node780;
	wire [1-1:0] node781;
	wire [1-1:0] node787;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node792;
	wire [1-1:0] node794;
	wire [1-1:0] node795;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node814;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node822;
	wire [1-1:0] node824;
	wire [1-1:0] node825;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node831;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node844;
	wire [1-1:0] node846;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node852;
	wire [1-1:0] node853;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node861;
	wire [1-1:0] node862;
	wire [1-1:0] node864;
	wire [1-1:0] node868;
	wire [1-1:0] node869;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node879;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node886;
	wire [1-1:0] node887;
	wire [1-1:0] node888;
	wire [1-1:0] node893;
	wire [1-1:0] node894;
	wire [1-1:0] node895;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node899;
	wire [1-1:0] node902;
	wire [1-1:0] node908;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node914;
	wire [1-1:0] node918;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node923;

	assign outp = (inp[3]) ? node452 : node1;
		assign node1 = (inp[9]) ? node179 : node2;
			assign node2 = (inp[0]) ? node68 : node3;
				assign node3 = (inp[11]) ? node17 : node4;
					assign node4 = (inp[7]) ? node6 : 1'b1;
						assign node6 = (inp[4]) ? node8 : 1'b1;
							assign node8 = (inp[12]) ? node10 : 1'b1;
								assign node10 = (inp[10]) ? node12 : 1'b1;
									assign node12 = (inp[5]) ? 1'b0 : node13;
										assign node13 = (inp[8]) ? 1'b0 : 1'b1;
					assign node17 = (inp[12]) ? node37 : node18;
						assign node18 = (inp[7]) ? node20 : 1'b1;
							assign node20 = (inp[8]) ? node22 : 1'b1;
								assign node22 = (inp[6]) ? node28 : node23;
									assign node23 = (inp[10]) ? node25 : 1'b1;
										assign node25 = (inp[5]) ? 1'b0 : 1'b1;
									assign node28 = (inp[2]) ? node32 : node29;
										assign node29 = (inp[5]) ? 1'b0 : 1'b1;
										assign node32 = (inp[1]) ? 1'b0 : node33;
											assign node33 = (inp[4]) ? 1'b0 : 1'b1;
						assign node37 = (inp[6]) ? node49 : node38;
							assign node38 = (inp[1]) ? node40 : 1'b1;
								assign node40 = (inp[5]) ? node42 : 1'b1;
									assign node42 = (inp[2]) ? 1'b0 : node43;
										assign node43 = (inp[10]) ? 1'b1 : node44;
											assign node44 = (inp[4]) ? 1'b0 : 1'b1;
							assign node49 = (inp[8]) ? node59 : node50;
								assign node50 = (inp[7]) ? node52 : 1'b1;
									assign node52 = (inp[10]) ? node54 : 1'b1;
										assign node54 = (inp[1]) ? 1'b0 : node55;
											assign node55 = (inp[4]) ? 1'b0 : 1'b1;
								assign node59 = (inp[4]) ? 1'b0 : node60;
									assign node60 = (inp[1]) ? 1'b0 : node61;
										assign node61 = (inp[7]) ? node63 : 1'b1;
											assign node63 = (inp[10]) ? 1'b0 : 1'b1;
				assign node68 = (inp[1]) ? node114 : node69;
					assign node69 = (inp[6]) ? node83 : node70;
						assign node70 = (inp[10]) ? node72 : 1'b1;
							assign node72 = (inp[12]) ? node80 : node73;
								assign node73 = (inp[2]) ? node75 : 1'b1;
									assign node75 = (inp[4]) ? node77 : 1'b1;
										assign node77 = (inp[11]) ? 1'b0 : 1'b1;
								assign node80 = (inp[5]) ? 1'b0 : 1'b1;
						assign node83 = (inp[8]) ? node95 : node84;
							assign node84 = (inp[2]) ? node86 : 1'b1;
								assign node86 = (inp[11]) ? node88 : 1'b1;
									assign node88 = (inp[7]) ? 1'b0 : node89;
										assign node89 = (inp[4]) ? node91 : 1'b1;
											assign node91 = (inp[12]) ? 1'b0 : 1'b1;
							assign node95 = (inp[11]) ? node109 : node96;
								assign node96 = (inp[4]) ? node98 : 1'b1;
									assign node98 = (inp[5]) ? 1'b0 : node99;
										assign node99 = (inp[12]) ? 1'b0 : node100;
											assign node100 = (inp[7]) ? node102 : 1'b1;
												assign node102 = (inp[2]) ? node104 : 1'b1;
													assign node104 = (inp[10]) ? 1'b0 : 1'b1;
								assign node109 = (inp[5]) ? 1'b0 : node110;
									assign node110 = (inp[2]) ? 1'b0 : 1'b1;
					assign node114 = (inp[11]) ? node140 : node115;
						assign node115 = (inp[12]) ? node123 : node116;
							assign node116 = (inp[7]) ? node118 : 1'b1;
								assign node118 = (inp[4]) ? node120 : 1'b1;
									assign node120 = (inp[8]) ? 1'b0 : 1'b1;
							assign node123 = (inp[5]) ? node131 : node124;
								assign node124 = (inp[2]) ? node126 : 1'b1;
									assign node126 = (inp[8]) ? 1'b0 : node127;
										assign node127 = (inp[7]) ? 1'b0 : 1'b1;
								assign node131 = (inp[10]) ? 1'b0 : node132;
									assign node132 = (inp[6]) ? 1'b0 : node133;
										assign node133 = (inp[7]) ? node135 : 1'b1;
											assign node135 = (inp[2]) ? 1'b0 : 1'b1;
						assign node140 = (inp[4]) ? node164 : node141;
							assign node141 = (inp[10]) ? node153 : node142;
								assign node142 = (inp[8]) ? node144 : 1'b1;
									assign node144 = (inp[5]) ? 1'b0 : node145;
										assign node145 = (inp[12]) ? node147 : 1'b1;
											assign node147 = (inp[6]) ? node149 : 1'b1;
												assign node149 = (inp[2]) ? 1'b0 : 1'b1;
								assign node153 = (inp[7]) ? node159 : node154;
									assign node154 = (inp[2]) ? node156 : 1'b1;
										assign node156 = (inp[5]) ? 1'b0 : 1'b1;
									assign node159 = (inp[12]) ? 1'b0 : node160;
										assign node160 = (inp[6]) ? 1'b0 : 1'b1;
							assign node164 = (inp[6]) ? 1'b0 : node165;
								assign node165 = (inp[7]) ? 1'b0 : node166;
									assign node166 = (inp[10]) ? node172 : node167;
										assign node167 = (inp[2]) ? node169 : 1'b1;
											assign node169 = (inp[12]) ? 1'b0 : 1'b1;
										assign node172 = (inp[8]) ? 1'b0 : node173;
											assign node173 = (inp[2]) ? 1'b0 : 1'b1;
			assign node179 = (inp[7]) ? node307 : node180;
				assign node180 = (inp[10]) ? node236 : node181;
					assign node181 = (inp[12]) ? node193 : node182;
						assign node182 = (inp[11]) ? node184 : 1'b1;
							assign node184 = (inp[8]) ? node186 : 1'b1;
								assign node186 = (inp[1]) ? node188 : 1'b1;
									assign node188 = (inp[0]) ? 1'b0 : node189;
										assign node189 = (inp[4]) ? 1'b0 : 1'b1;
						assign node193 = (inp[4]) ? node205 : node194;
							assign node194 = (inp[1]) ? node196 : 1'b1;
								assign node196 = (inp[0]) ? node198 : 1'b1;
									assign node198 = (inp[2]) ? 1'b0 : node199;
										assign node199 = (inp[5]) ? node201 : 1'b1;
											assign node201 = (inp[8]) ? 1'b0 : 1'b1;
							assign node205 = (inp[2]) ? node223 : node206;
								assign node206 = (inp[11]) ? node216 : node207;
									assign node207 = (inp[1]) ? node209 : 1'b1;
										assign node209 = (inp[0]) ? node211 : 1'b1;
											assign node211 = (inp[8]) ? 1'b0 : node212;
												assign node212 = (inp[6]) ? 1'b0 : 1'b1;
									assign node216 = (inp[8]) ? node218 : 1'b1;
										assign node218 = (inp[6]) ? 1'b0 : node219;
											assign node219 = (inp[5]) ? 1'b0 : 1'b1;
								assign node223 = (inp[8]) ? 1'b0 : node224;
									assign node224 = (inp[11]) ? node230 : node225;
										assign node225 = (inp[6]) ? node227 : 1'b1;
											assign node227 = (inp[1]) ? 1'b0 : 1'b1;
										assign node230 = (inp[0]) ? 1'b0 : node231;
											assign node231 = (inp[5]) ? 1'b0 : 1'b1;
					assign node236 = (inp[5]) ? node268 : node237;
						assign node237 = (inp[2]) ? node249 : node238;
							assign node238 = (inp[8]) ? node240 : 1'b1;
								assign node240 = (inp[6]) ? node242 : 1'b1;
									assign node242 = (inp[12]) ? node244 : 1'b1;
										assign node244 = (inp[0]) ? 1'b0 : node245;
											assign node245 = (inp[4]) ? 1'b1 : 1'b0;
							assign node249 = (inp[1]) ? node259 : node250;
								assign node250 = (inp[6]) ? node252 : 1'b1;
									assign node252 = (inp[0]) ? node254 : 1'b1;
										assign node254 = (inp[8]) ? 1'b0 : node255;
											assign node255 = (inp[12]) ? 1'b0 : 1'b1;
								assign node259 = (inp[11]) ? 1'b0 : node260;
									assign node260 = (inp[4]) ? node262 : 1'b1;
										assign node262 = (inp[0]) ? 1'b0 : node263;
											assign node263 = (inp[6]) ? 1'b1 : 1'b0;
						assign node268 = (inp[0]) ? node296 : node269;
							assign node269 = (inp[6]) ? node281 : node270;
								assign node270 = (inp[12]) ? node278 : node271;
									assign node271 = (inp[2]) ? node273 : 1'b1;
										assign node273 = (inp[1]) ? node275 : 1'b1;
											assign node275 = (inp[8]) ? 1'b0 : 1'b1;
									assign node278 = (inp[8]) ? 1'b0 : 1'b1;
								assign node281 = (inp[11]) ? 1'b0 : node282;
									assign node282 = (inp[4]) ? node288 : node283;
										assign node283 = (inp[2]) ? node285 : 1'b1;
											assign node285 = (inp[1]) ? 1'b0 : 1'b1;
										assign node288 = (inp[8]) ? 1'b0 : node289;
											assign node289 = (inp[2]) ? 1'b0 : node290;
												assign node290 = (inp[12]) ? 1'b0 : 1'b1;
							assign node296 = (inp[1]) ? 1'b0 : node297;
								assign node297 = (inp[12]) ? 1'b0 : node298;
									assign node298 = (inp[4]) ? node300 : 1'b1;
										assign node300 = (inp[2]) ? 1'b0 : node301;
											assign node301 = (inp[11]) ? 1'b0 : 1'b1;
				assign node307 = (inp[1]) ? node367 : node308;
					assign node308 = (inp[10]) ? node340 : node309;
						assign node309 = (inp[5]) ? node325 : node310;
							assign node310 = (inp[12]) ? node312 : 1'b1;
								assign node312 = (inp[8]) ? node314 : 1'b1;
									assign node314 = (inp[4]) ? node320 : node315;
										assign node315 = (inp[6]) ? node317 : 1'b1;
											assign node317 = (inp[11]) ? 1'b0 : 1'b1;
										assign node320 = (inp[0]) ? 1'b0 : node321;
											assign node321 = (inp[11]) ? 1'b0 : 1'b1;
							assign node325 = (inp[4]) ? node331 : node326;
								assign node326 = (inp[11]) ? node328 : 1'b1;
									assign node328 = (inp[0]) ? 1'b0 : 1'b1;
								assign node331 = (inp[2]) ? 1'b0 : node332;
									assign node332 = (inp[0]) ? 1'b0 : node333;
										assign node333 = (inp[12]) ? node335 : 1'b1;
											assign node335 = (inp[8]) ? 1'b0 : 1'b1;
						assign node340 = (inp[6]) ? node356 : node341;
							assign node341 = (inp[8]) ? node347 : node342;
								assign node342 = (inp[5]) ? node344 : 1'b1;
									assign node344 = (inp[4]) ? 1'b0 : 1'b1;
								assign node347 = (inp[12]) ? 1'b0 : node348;
									assign node348 = (inp[4]) ? node350 : 1'b1;
										assign node350 = (inp[11]) ? 1'b0 : node351;
											assign node351 = (inp[5]) ? 1'b1 : 1'b0;
							assign node356 = (inp[2]) ? 1'b0 : node357;
								assign node357 = (inp[5]) ? 1'b0 : node358;
									assign node358 = (inp[12]) ? node360 : 1'b1;
										assign node360 = (inp[11]) ? 1'b0 : node361;
											assign node361 = (inp[0]) ? 1'b1 : 1'b0;
					assign node367 = (inp[11]) ? node421 : node368;
						assign node368 = (inp[2]) ? node396 : node369;
							assign node369 = (inp[0]) ? node379 : node370;
								assign node370 = (inp[8]) ? node372 : 1'b1;
									assign node372 = (inp[5]) ? 1'b0 : node373;
										assign node373 = (inp[12]) ? node375 : 1'b1;
											assign node375 = (inp[4]) ? 1'b0 : 1'b1;
								assign node379 = (inp[6]) ? node391 : node380;
									assign node380 = (inp[4]) ? node386 : node381;
										assign node381 = (inp[10]) ? node383 : 1'b1;
											assign node383 = (inp[5]) ? 1'b0 : 1'b1;
										assign node386 = (inp[5]) ? 1'b0 : node387;
											assign node387 = (inp[10]) ? 1'b0 : 1'b1;
									assign node391 = (inp[5]) ? 1'b0 : node392;
										assign node392 = (inp[12]) ? 1'b0 : 1'b1;
							assign node396 = (inp[0]) ? node412 : node397;
								assign node397 = (inp[12]) ? 1'b0 : node398;
									assign node398 = (inp[5]) ? node406 : node399;
										assign node399 = (inp[6]) ? node401 : 1'b1;
											assign node401 = (inp[4]) ? node403 : 1'b1;
												assign node403 = (inp[10]) ? 1'b0 : 1'b1;
										assign node406 = (inp[4]) ? 1'b0 : node407;
											assign node407 = (inp[10]) ? 1'b0 : 1'b1;
								assign node412 = (inp[4]) ? 1'b0 : node413;
									assign node413 = (inp[10]) ? 1'b0 : node414;
										assign node414 = (inp[5]) ? 1'b0 : node415;
											assign node415 = (inp[8]) ? 1'b0 : 1'b1;
						assign node421 = (inp[5]) ? node443 : node422;
							assign node422 = (inp[0]) ? 1'b0 : node423;
								assign node423 = (inp[6]) ? node433 : node424;
									assign node424 = (inp[4]) ? node426 : 1'b1;
										assign node426 = (inp[12]) ? 1'b0 : node427;
											assign node427 = (inp[10]) ? node429 : 1'b1;
												assign node429 = (inp[8]) ? 1'b0 : 1'b1;
									assign node433 = (inp[4]) ? 1'b0 : node434;
										assign node434 = (inp[12]) ? 1'b0 : node435;
											assign node435 = (inp[8]) ? 1'b0 : node436;
												assign node436 = (inp[10]) ? 1'b0 : 1'b1;
							assign node443 = (inp[4]) ? 1'b0 : node444;
								assign node444 = (inp[2]) ? 1'b0 : node445;
									assign node445 = (inp[12]) ? 1'b0 : node446;
										assign node446 = (inp[8]) ? 1'b0 : 1'b1;
		assign node452 = (inp[0]) ? node710 : node453;
			assign node453 = (inp[12]) ? node587 : node454;
				assign node454 = (inp[7]) ? node512 : node455;
					assign node455 = (inp[10]) ? node479 : node456;
						assign node456 = (inp[2]) ? node458 : 1'b1;
							assign node458 = (inp[9]) ? node468 : node459;
								assign node459 = (inp[5]) ? node461 : 1'b1;
									assign node461 = (inp[4]) ? node463 : 1'b1;
										assign node463 = (inp[11]) ? node465 : 1'b1;
											assign node465 = (inp[1]) ? 1'b0 : 1'b1;
								assign node468 = (inp[4]) ? node476 : node469;
									assign node469 = (inp[6]) ? node471 : 1'b1;
										assign node471 = (inp[5]) ? node473 : 1'b1;
											assign node473 = (inp[11]) ? 1'b0 : 1'b1;
									assign node476 = (inp[1]) ? 1'b0 : 1'b1;
						assign node479 = (inp[5]) ? node501 : node480;
							assign node480 = (inp[11]) ? node490 : node481;
								assign node481 = (inp[2]) ? node483 : 1'b1;
									assign node483 = (inp[1]) ? node485 : 1'b1;
										assign node485 = (inp[4]) ? node487 : 1'b1;
											assign node487 = (inp[9]) ? 1'b0 : 1'b1;
								assign node490 = (inp[4]) ? node492 : 1'b1;
									assign node492 = (inp[6]) ? 1'b0 : node493;
										assign node493 = (inp[1]) ? node495 : 1'b1;
											assign node495 = (inp[8]) ? 1'b0 : node496;
												assign node496 = (inp[9]) ? 1'b0 : 1'b1;
							assign node501 = (inp[6]) ? node507 : node502;
								assign node502 = (inp[8]) ? node504 : 1'b1;
									assign node504 = (inp[4]) ? 1'b0 : 1'b1;
								assign node507 = (inp[9]) ? 1'b0 : node508;
									assign node508 = (inp[1]) ? 1'b0 : 1'b1;
					assign node512 = (inp[4]) ? node554 : node513;
						assign node513 = (inp[8]) ? node529 : node514;
							assign node514 = (inp[11]) ? node516 : 1'b1;
								assign node516 = (inp[1]) ? node524 : node517;
									assign node517 = (inp[2]) ? node519 : 1'b1;
										assign node519 = (inp[5]) ? node521 : 1'b1;
											assign node521 = (inp[9]) ? 1'b0 : 1'b1;
									assign node524 = (inp[5]) ? 1'b0 : node525;
										assign node525 = (inp[10]) ? 1'b0 : 1'b1;
							assign node529 = (inp[1]) ? node545 : node530;
								assign node530 = (inp[9]) ? node538 : node531;
									assign node531 = (inp[11]) ? node533 : 1'b1;
										assign node533 = (inp[2]) ? node535 : 1'b1;
											assign node535 = (inp[5]) ? 1'b0 : 1'b1;
									assign node538 = (inp[2]) ? 1'b0 : node539;
										assign node539 = (inp[11]) ? node541 : 1'b1;
											assign node541 = (inp[10]) ? 1'b0 : 1'b1;
								assign node545 = (inp[11]) ? 1'b0 : node546;
									assign node546 = (inp[2]) ? node548 : 1'b1;
										assign node548 = (inp[6]) ? 1'b0 : node549;
											assign node549 = (inp[5]) ? 1'b0 : 1'b1;
						assign node554 = (inp[10]) ? node580 : node555;
							assign node555 = (inp[6]) ? node567 : node556;
								assign node556 = (inp[8]) ? node558 : 1'b1;
									assign node558 = (inp[9]) ? node564 : node559;
										assign node559 = (inp[11]) ? node561 : 1'b1;
											assign node561 = (inp[5]) ? 1'b0 : 1'b1;
										assign node564 = (inp[1]) ? 1'b0 : 1'b1;
								assign node567 = (inp[9]) ? 1'b0 : node568;
									assign node568 = (inp[5]) ? node574 : node569;
										assign node569 = (inp[1]) ? 1'b1 : node570;
											assign node570 = (inp[11]) ? 1'b0 : 1'b1;
										assign node574 = (inp[11]) ? 1'b0 : node575;
											assign node575 = (inp[2]) ? 1'b0 : 1'b1;
							assign node580 = (inp[9]) ? 1'b0 : node581;
								assign node581 = (inp[6]) ? 1'b0 : node582;
									assign node582 = (inp[2]) ? 1'b0 : 1'b1;
				assign node587 = (inp[1]) ? node657 : node588;
					assign node588 = (inp[8]) ? node624 : node589;
						assign node589 = (inp[11]) ? node599 : node590;
							assign node590 = (inp[2]) ? node592 : 1'b1;
								assign node592 = (inp[9]) ? node594 : 1'b1;
									assign node594 = (inp[10]) ? 1'b0 : node595;
										assign node595 = (inp[6]) ? 1'b0 : 1'b1;
							assign node599 = (inp[10]) ? node613 : node600;
								assign node600 = (inp[5]) ? node602 : 1'b1;
									assign node602 = (inp[2]) ? node608 : node603;
										assign node603 = (inp[6]) ? node605 : 1'b1;
											assign node605 = (inp[4]) ? 1'b0 : 1'b1;
										assign node608 = (inp[7]) ? 1'b0 : node609;
											assign node609 = (inp[9]) ? 1'b0 : 1'b1;
								assign node613 = (inp[6]) ? 1'b0 : node614;
									assign node614 = (inp[7]) ? node616 : 1'b1;
										assign node616 = (inp[2]) ? 1'b0 : node617;
											assign node617 = (inp[9]) ? node619 : 1'b1;
												assign node619 = (inp[5]) ? 1'b0 : 1'b1;
						assign node624 = (inp[10]) ? node646 : node625;
							assign node625 = (inp[6]) ? node631 : node626;
								assign node626 = (inp[5]) ? node628 : 1'b1;
									assign node628 = (inp[7]) ? 1'b0 : 1'b1;
								assign node631 = (inp[11]) ? node639 : node632;
									assign node632 = (inp[4]) ? 1'b0 : node633;
										assign node633 = (inp[7]) ? node635 : 1'b1;
											assign node635 = (inp[5]) ? 1'b0 : 1'b1;
									assign node639 = (inp[7]) ? 1'b0 : node640;
										assign node640 = (inp[9]) ? 1'b0 : node641;
											assign node641 = (inp[2]) ? 1'b0 : 1'b1;
							assign node646 = (inp[5]) ? 1'b0 : node647;
								assign node647 = (inp[9]) ? 1'b0 : node648;
									assign node648 = (inp[2]) ? node650 : 1'b1;
										assign node650 = (inp[6]) ? 1'b0 : node651;
											assign node651 = (inp[11]) ? 1'b0 : 1'b1;
					assign node657 = (inp[2]) ? node691 : node658;
						assign node658 = (inp[7]) ? node680 : node659;
							assign node659 = (inp[8]) ? node671 : node660;
								assign node660 = (inp[4]) ? node668 : node661;
									assign node661 = (inp[9]) ? node663 : 1'b1;
										assign node663 = (inp[11]) ? node665 : 1'b1;
											assign node665 = (inp[6]) ? 1'b0 : 1'b1;
									assign node668 = (inp[10]) ? 1'b0 : 1'b1;
								assign node671 = (inp[9]) ? 1'b0 : node672;
									assign node672 = (inp[6]) ? 1'b0 : node673;
										assign node673 = (inp[11]) ? node675 : 1'b1;
											assign node675 = (inp[5]) ? 1'b0 : 1'b1;
							assign node680 = (inp[4]) ? 1'b0 : node681;
								assign node681 = (inp[6]) ? 1'b0 : node682;
									assign node682 = (inp[9]) ? node684 : 1'b1;
										assign node684 = (inp[5]) ? 1'b0 : node685;
											assign node685 = (inp[10]) ? 1'b0 : 1'b1;
						assign node691 = (inp[10]) ? 1'b0 : node692;
							assign node692 = (inp[8]) ? 1'b0 : node693;
								assign node693 = (inp[4]) ? node697 : node694;
									assign node694 = (inp[6]) ? 1'b0 : 1'b1;
									assign node697 = (inp[9]) ? 1'b0 : node698;
										assign node698 = (inp[11]) ? 1'b0 : node699;
											assign node699 = (inp[5]) ? 1'b0 : node700;
												assign node700 = (inp[7]) ? node702 : 1'b1;
													assign node702 = (inp[6]) ? 1'b0 : 1'b1;
			assign node710 = (inp[11]) ? node838 : node711;
				assign node711 = (inp[9]) ? node787 : node712;
					assign node712 = (inp[1]) ? node748 : node713;
						assign node713 = (inp[10]) ? node725 : node714;
							assign node714 = (inp[4]) ? node716 : 1'b1;
								assign node716 = (inp[7]) ? node718 : 1'b1;
									assign node718 = (inp[5]) ? 1'b0 : node719;
										assign node719 = (inp[12]) ? node721 : 1'b1;
											assign node721 = (inp[8]) ? 1'b0 : 1'b1;
							assign node725 = (inp[5]) ? node735 : node726;
								assign node726 = (inp[7]) ? node728 : 1'b1;
									assign node728 = (inp[12]) ? 1'b0 : node729;
										assign node729 = (inp[8]) ? node731 : 1'b1;
											assign node731 = (inp[6]) ? 1'b0 : 1'b1;
								assign node735 = (inp[6]) ? node741 : node736;
									assign node736 = (inp[12]) ? node738 : 1'b1;
										assign node738 = (inp[8]) ? 1'b0 : 1'b1;
									assign node741 = (inp[4]) ? 1'b0 : node742;
										assign node742 = (inp[12]) ? node744 : 1'b0;
											assign node744 = (inp[7]) ? 1'b0 : 1'b1;
						assign node748 = (inp[8]) ? node772 : node749;
							assign node749 = (inp[6]) ? node761 : node750;
								assign node750 = (inp[12]) ? node752 : 1'b1;
									assign node752 = (inp[2]) ? node754 : 1'b1;
										assign node754 = (inp[10]) ? 1'b0 : node755;
											assign node755 = (inp[4]) ? node757 : 1'b1;
												assign node757 = (inp[7]) ? 1'b0 : 1'b1;
								assign node761 = (inp[2]) ? node767 : node762;
									assign node762 = (inp[5]) ? node764 : 1'b1;
										assign node764 = (inp[12]) ? 1'b1 : 1'b0;
									assign node767 = (inp[5]) ? 1'b0 : node768;
										assign node768 = (inp[7]) ? 1'b0 : 1'b1;
							assign node772 = (inp[10]) ? 1'b0 : node773;
								assign node773 = (inp[6]) ? 1'b0 : node774;
									assign node774 = (inp[7]) ? node780 : node775;
										assign node775 = (inp[5]) ? node777 : 1'b1;
											assign node777 = (inp[2]) ? 1'b0 : 1'b1;
										assign node780 = (inp[12]) ? 1'b0 : node781;
											assign node781 = (inp[5]) ? 1'b0 : 1'b1;
					assign node787 = (inp[8]) ? node819 : node788;
						assign node788 = (inp[7]) ? node810 : node789;
							assign node789 = (inp[2]) ? node799 : node790;
								assign node790 = (inp[6]) ? node792 : 1'b1;
									assign node792 = (inp[1]) ? node794 : 1'b1;
										assign node794 = (inp[12]) ? 1'b0 : node795;
											assign node795 = (inp[4]) ? 1'b0 : 1'b1;
								assign node799 = (inp[5]) ? 1'b0 : node800;
									assign node800 = (inp[4]) ? node804 : node801;
										assign node801 = (inp[1]) ? 1'b0 : 1'b1;
										assign node804 = (inp[10]) ? 1'b0 : node805;
											assign node805 = (inp[6]) ? 1'b0 : 1'b1;
							assign node810 = (inp[12]) ? 1'b0 : node811;
								assign node811 = (inp[6]) ? 1'b0 : node812;
									assign node812 = (inp[5]) ? node814 : 1'b1;
										assign node814 = (inp[1]) ? 1'b0 : 1'b1;
						assign node819 = (inp[12]) ? 1'b0 : node820;
							assign node820 = (inp[10]) ? 1'b0 : node821;
								assign node821 = (inp[2]) ? node829 : node822;
									assign node822 = (inp[1]) ? node824 : 1'b1;
										assign node824 = (inp[5]) ? 1'b0 : node825;
											assign node825 = (inp[4]) ? 1'b0 : 1'b1;
									assign node829 = (inp[6]) ? 1'b0 : node830;
										assign node830 = (inp[1]) ? 1'b0 : node831;
											assign node831 = (inp[4]) ? 1'b0 : 1'b1;
				assign node838 = (inp[5]) ? node908 : node839;
					assign node839 = (inp[4]) ? node893 : node840;
						assign node840 = (inp[1]) ? node868 : node841;
							assign node841 = (inp[10]) ? node849 : node842;
								assign node842 = (inp[12]) ? node844 : 1'b1;
									assign node844 = (inp[9]) ? node846 : 1'b1;
										assign node846 = (inp[2]) ? 1'b0 : 1'b1;
								assign node849 = (inp[2]) ? node861 : node850;
									assign node850 = (inp[6]) ? node852 : 1'b1;
										assign node852 = (inp[12]) ? 1'b0 : node853;
											assign node853 = (inp[7]) ? node855 : 1'b1;
												assign node855 = (inp[9]) ? 1'b0 : node856;
													assign node856 = (inp[8]) ? 1'b0 : 1'b1;
									assign node861 = (inp[9]) ? 1'b0 : node862;
										assign node862 = (inp[6]) ? node864 : 1'b0;
											assign node864 = (inp[7]) ? 1'b0 : 1'b1;
							assign node868 = (inp[12]) ? node886 : node869;
								assign node869 = (inp[8]) ? node879 : node870;
									assign node870 = (inp[10]) ? 1'b0 : node871;
										assign node871 = (inp[9]) ? node873 : 1'b1;
											assign node873 = (inp[2]) ? 1'b0 : node874;
												assign node874 = (inp[6]) ? 1'b0 : 1'b1;
									assign node879 = (inp[2]) ? node881 : 1'b0;
										assign node881 = (inp[7]) ? 1'b0 : node882;
											assign node882 = (inp[9]) ? 1'b0 : 1'b1;
								assign node886 = (inp[2]) ? 1'b0 : node887;
									assign node887 = (inp[6]) ? 1'b0 : node888;
										assign node888 = (inp[8]) ? 1'b0 : 1'b1;
						assign node893 = (inp[12]) ? 1'b0 : node894;
							assign node894 = (inp[2]) ? 1'b0 : node895;
								assign node895 = (inp[10]) ? 1'b0 : node896;
									assign node896 = (inp[6]) ? node902 : node897;
										assign node897 = (inp[1]) ? node899 : 1'b1;
											assign node899 = (inp[7]) ? 1'b0 : 1'b1;
										assign node902 = (inp[8]) ? 1'b0 : 1'b1;
					assign node908 = (inp[1]) ? 1'b0 : node909;
						assign node909 = (inp[2]) ? 1'b0 : node910;
							assign node910 = (inp[6]) ? node918 : node911;
								assign node911 = (inp[4]) ? 1'b0 : node912;
									assign node912 = (inp[12]) ? node914 : 1'b1;
										assign node914 = (inp[10]) ? 1'b0 : 1'b1;
								assign node918 = (inp[8]) ? 1'b0 : node919;
									assign node919 = (inp[9]) ? 1'b0 : node920;
										assign node920 = (inp[10]) ? 1'b0 : node921;
											assign node921 = (inp[12]) ? node923 : 1'b1;
												assign node923 = (inp[4]) ? 1'b0 : 1'b1;

endmodule