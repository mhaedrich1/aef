module dtc_split75_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node444;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node630;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node681;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node753;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node798;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1032;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1104;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1120;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1167;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1198;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1277;
	wire [3-1:0] node1279;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1288;
	wire [3-1:0] node1290;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1301;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1319;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1327;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1341;
	wire [3-1:0] node1343;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1357;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1370;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1391;
	wire [3-1:0] node1393;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1399;
	wire [3-1:0] node1402;
	wire [3-1:0] node1404;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1411;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1427;
	wire [3-1:0] node1428;
	wire [3-1:0] node1432;
	wire [3-1:0] node1434;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1444;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1462;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1470;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;
	wire [3-1:0] node1523;
	wire [3-1:0] node1525;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1531;
	wire [3-1:0] node1534;
	wire [3-1:0] node1536;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1548;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1558;
	wire [3-1:0] node1561;
	wire [3-1:0] node1562;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1575;
	wire [3-1:0] node1577;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1583;
	wire [3-1:0] node1585;
	wire [3-1:0] node1588;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1597;
	wire [3-1:0] node1599;
	wire [3-1:0] node1602;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1609;
	wire [3-1:0] node1610;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1614;
	wire [3-1:0] node1619;
	wire [3-1:0] node1621;
	wire [3-1:0] node1624;
	wire [3-1:0] node1626;
	wire [3-1:0] node1628;
	wire [3-1:0] node1631;
	wire [3-1:0] node1632;
	wire [3-1:0] node1633;
	wire [3-1:0] node1635;
	wire [3-1:0] node1637;
	wire [3-1:0] node1642;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1647;
	wire [3-1:0] node1649;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1654;
	wire [3-1:0] node1657;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1670;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1677;
	wire [3-1:0] node1679;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1687;
	wire [3-1:0] node1688;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1696;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;

	assign outp = (inp[10]) ? node876 : node1;
		assign node1 = (inp[9]) ? node467 : node2;
			assign node2 = (inp[2]) ? node136 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[3]) ? node86 : node5;
						assign node5 = (inp[5]) ? node45 : node6;
							assign node6 = (inp[6]) ? node20 : node7;
								assign node7 = (inp[7]) ? node15 : node8;
									assign node8 = (inp[8]) ? node10 : 3'b000;
										assign node10 = (inp[4]) ? 3'b000 : node11;
											assign node11 = (inp[1]) ? 3'b100 : 3'b111;
									assign node15 = (inp[4]) ? 3'b100 : node16;
										assign node16 = (inp[8]) ? 3'b000 : 3'b100;
								assign node20 = (inp[11]) ? node34 : node21;
									assign node21 = (inp[7]) ? node29 : node22;
										assign node22 = (inp[1]) ? 3'b110 : node23;
											assign node23 = (inp[8]) ? 3'b111 : node24;
												assign node24 = (inp[4]) ? 3'b010 : 3'b111;
										assign node29 = (inp[8]) ? 3'b010 : node30;
											assign node30 = (inp[4]) ? 3'b110 : 3'b010;
									assign node34 = (inp[7]) ? node40 : node35;
										assign node35 = (inp[4]) ? 3'b000 : node36;
											assign node36 = (inp[8]) ? 3'b111 : 3'b000;
										assign node40 = (inp[4]) ? 3'b100 : node41;
											assign node41 = (inp[8]) ? 3'b000 : 3'b100;
							assign node45 = (inp[6]) ? node59 : node46;
								assign node46 = (inp[7]) ? node54 : node47;
									assign node47 = (inp[4]) ? 3'b010 : node48;
										assign node48 = (inp[8]) ? node50 : 3'b010;
											assign node50 = (inp[1]) ? 3'b110 : 3'b111;
									assign node54 = (inp[8]) ? node56 : 3'b110;
										assign node56 = (inp[4]) ? 3'b110 : 3'b010;
								assign node59 = (inp[11]) ? node73 : node60;
									assign node60 = (inp[7]) ? node68 : node61;
										assign node61 = (inp[8]) ? node63 : 3'b000;
											assign node63 = (inp[4]) ? 3'b000 : node64;
												assign node64 = (inp[1]) ? 3'b100 : 3'b111;
										assign node68 = (inp[4]) ? 3'b100 : node69;
											assign node69 = (inp[8]) ? 3'b000 : 3'b100;
									assign node73 = (inp[7]) ? node81 : node74;
										assign node74 = (inp[4]) ? 3'b010 : node75;
											assign node75 = (inp[8]) ? node77 : 3'b010;
												assign node77 = (inp[1]) ? 3'b110 : 3'b111;
										assign node81 = (inp[4]) ? 3'b110 : node82;
											assign node82 = (inp[1]) ? 3'b010 : 3'b110;
						assign node86 = (inp[1]) ? node88 : 3'b111;
							assign node88 = (inp[7]) ? node108 : node89;
								assign node89 = (inp[8]) ? node99 : node90;
									assign node90 = (inp[5]) ? node94 : node91;
										assign node91 = (inp[6]) ? 3'b010 : 3'b000;
										assign node94 = (inp[6]) ? node96 : 3'b010;
											assign node96 = (inp[11]) ? 3'b010 : 3'b000;
									assign node99 = (inp[4]) ? node101 : 3'b111;
										assign node101 = (inp[11]) ? node105 : node102;
											assign node102 = (inp[5]) ? 3'b000 : 3'b111;
											assign node105 = (inp[5]) ? 3'b010 : 3'b000;
								assign node108 = (inp[4]) ? node124 : node109;
									assign node109 = (inp[8]) ? node115 : node110;
										assign node110 = (inp[5]) ? 3'b100 : node111;
											assign node111 = (inp[6]) ? 3'b010 : 3'b100;
										assign node115 = (inp[11]) ? 3'b010 : node116;
											assign node116 = (inp[6]) ? node120 : node117;
												assign node117 = (inp[5]) ? 3'b010 : 3'b000;
												assign node120 = (inp[5]) ? 3'b000 : 3'b010;
									assign node124 = (inp[5]) ? node130 : node125;
										assign node125 = (inp[11]) ? 3'b100 : node126;
											assign node126 = (inp[6]) ? 3'b010 : 3'b100;
										assign node130 = (inp[6]) ? node132 : 3'b110;
											assign node132 = (inp[11]) ? 3'b110 : 3'b100;
				assign node136 = (inp[1]) ? node282 : node137;
					assign node137 = (inp[0]) ? node233 : node138;
						assign node138 = (inp[11]) ? node198 : node139;
							assign node139 = (inp[4]) ? node165 : node140;
								assign node140 = (inp[3]) ? node146 : node141;
									assign node141 = (inp[5]) ? 3'b000 : node142;
										assign node142 = (inp[8]) ? 3'b100 : 3'b000;
									assign node146 = (inp[7]) ? node158 : node147;
										assign node147 = (inp[8]) ? node153 : node148;
											assign node148 = (inp[5]) ? node150 : 3'b110;
												assign node150 = (inp[6]) ? 3'b000 : 3'b010;
											assign node153 = (inp[5]) ? node155 : 3'b100;
												assign node155 = (inp[6]) ? 3'b100 : 3'b110;
										assign node158 = (inp[6]) ? node160 : 3'b000;
											assign node160 = (inp[8]) ? node162 : 3'b000;
												assign node162 = (inp[5]) ? 3'b000 : 3'b010;
								assign node165 = (inp[5]) ? node183 : node166;
									assign node166 = (inp[8]) ? node176 : node167;
										assign node167 = (inp[3]) ? node171 : node168;
											assign node168 = (inp[7]) ? 3'b010 : 3'b100;
											assign node171 = (inp[6]) ? 3'b010 : node172;
												assign node172 = (inp[7]) ? 3'b100 : 3'b000;
										assign node176 = (inp[6]) ? node178 : 3'b000;
											assign node178 = (inp[7]) ? 3'b000 : node179;
												assign node179 = (inp[3]) ? 3'b110 : 3'b000;
									assign node183 = (inp[6]) ? node189 : node184;
										assign node184 = (inp[3]) ? node186 : 3'b100;
											assign node186 = (inp[7]) ? 3'b100 : 3'b010;
										assign node189 = (inp[3]) ? node195 : node190;
											assign node190 = (inp[7]) ? node192 : 3'b100;
												assign node192 = (inp[8]) ? 3'b010 : 3'b110;
											assign node195 = (inp[8]) ? 3'b000 : 3'b100;
							assign node198 = (inp[5]) ? node226 : node199;
								assign node199 = (inp[3]) ? node213 : node200;
									assign node200 = (inp[7]) ? node208 : node201;
										assign node201 = (inp[4]) ? node205 : node202;
											assign node202 = (inp[8]) ? 3'b100 : 3'b010;
											assign node205 = (inp[8]) ? 3'b010 : 3'b110;
										assign node208 = (inp[4]) ? node210 : 3'b010;
											assign node210 = (inp[8]) ? 3'b000 : 3'b100;
									assign node213 = (inp[7]) ? node219 : node214;
										assign node214 = (inp[8]) ? node216 : 3'b000;
											assign node216 = (inp[4]) ? 3'b000 : 3'b100;
										assign node219 = (inp[4]) ? node223 : node220;
											assign node220 = (inp[8]) ? 3'b000 : 3'b010;
											assign node223 = (inp[8]) ? 3'b010 : 3'b110;
								assign node226 = (inp[4]) ? node228 : 3'b010;
									assign node228 = (inp[3]) ? node230 : 3'b110;
										assign node230 = (inp[7]) ? 3'b110 : 3'b010;
						assign node233 = (inp[3]) ? 3'b110 : node234;
							assign node234 = (inp[5]) ? node262 : node235;
								assign node235 = (inp[11]) ? node251 : node236;
									assign node236 = (inp[6]) ? node244 : node237;
										assign node237 = (inp[8]) ? node241 : node238;
											assign node238 = (inp[7]) ? 3'b100 : 3'b000;
											assign node241 = (inp[7]) ? 3'b000 : 3'b110;
										assign node244 = (inp[7]) ? node246 : 3'b110;
											assign node246 = (inp[8]) ? 3'b010 : node247;
												assign node247 = (inp[4]) ? 3'b110 : 3'b010;
									assign node251 = (inp[7]) ? node257 : node252;
										assign node252 = (inp[8]) ? node254 : 3'b000;
											assign node254 = (inp[4]) ? 3'b000 : 3'b110;
										assign node257 = (inp[4]) ? 3'b100 : node258;
											assign node258 = (inp[8]) ? 3'b000 : 3'b100;
								assign node262 = (inp[7]) ? node272 : node263;
									assign node263 = (inp[4]) ? node267 : node264;
										assign node264 = (inp[8]) ? 3'b110 : 3'b010;
										assign node267 = (inp[11]) ? 3'b010 : node268;
											assign node268 = (inp[6]) ? 3'b000 : 3'b010;
									assign node272 = (inp[8]) ? node278 : node273;
										assign node273 = (inp[11]) ? 3'b110 : node274;
											assign node274 = (inp[6]) ? 3'b100 : 3'b110;
										assign node278 = (inp[4]) ? 3'b110 : 3'b010;
					assign node282 = (inp[7]) ? node400 : node283;
						assign node283 = (inp[11]) ? node361 : node284;
							assign node284 = (inp[3]) ? node324 : node285;
								assign node285 = (inp[0]) ? node305 : node286;
									assign node286 = (inp[4]) ? node296 : node287;
										assign node287 = (inp[6]) ? node293 : node288;
											assign node288 = (inp[8]) ? 3'b010 : node289;
												assign node289 = (inp[5]) ? 3'b110 : 3'b010;
											assign node293 = (inp[5]) ? 3'b110 : 3'b100;
										assign node296 = (inp[5]) ? node300 : node297;
											assign node297 = (inp[6]) ? 3'b010 : 3'b100;
											assign node300 = (inp[6]) ? node302 : 3'b000;
												assign node302 = (inp[8]) ? 3'b000 : 3'b100;
									assign node305 = (inp[5]) ? node319 : node306;
										assign node306 = (inp[6]) ? node314 : node307;
											assign node307 = (inp[8]) ? node311 : node308;
												assign node308 = (inp[4]) ? 3'b100 : 3'b000;
												assign node311 = (inp[4]) ? 3'b000 : 3'b100;
											assign node314 = (inp[8]) ? 3'b110 : node315;
												assign node315 = (inp[4]) ? 3'b100 : 3'b000;
										assign node319 = (inp[4]) ? node321 : 3'b000;
											assign node321 = (inp[8]) ? 3'b000 : 3'b010;
								assign node324 = (inp[8]) ? node346 : node325;
									assign node325 = (inp[4]) ? node339 : node326;
										assign node326 = (inp[0]) ? node334 : node327;
											assign node327 = (inp[5]) ? node331 : node328;
												assign node328 = (inp[6]) ? 3'b000 : 3'b010;
												assign node331 = (inp[6]) ? 3'b010 : 3'b100;
											assign node334 = (inp[5]) ? 3'b000 : node335;
												assign node335 = (inp[6]) ? 3'b110 : 3'b000;
										assign node339 = (inp[0]) ? node341 : 3'b010;
											assign node341 = (inp[5]) ? node343 : 3'b010;
												assign node343 = (inp[6]) ? 3'b000 : 3'b010;
									assign node346 = (inp[5]) ? node354 : node347;
										assign node347 = (inp[4]) ? node349 : 3'b110;
											assign node349 = (inp[0]) ? 3'b000 : node350;
												assign node350 = (inp[6]) ? 3'b100 : 3'b110;
										assign node354 = (inp[0]) ? node358 : node355;
											assign node355 = (inp[4]) ? 3'b010 : 3'b000;
											assign node358 = (inp[4]) ? 3'b010 : 3'b110;
							assign node361 = (inp[5]) ? node387 : node362;
								assign node362 = (inp[8]) ? node374 : node363;
									assign node363 = (inp[3]) ? node369 : node364;
										assign node364 = (inp[4]) ? node366 : 3'b010;
											assign node366 = (inp[0]) ? 3'b000 : 3'b010;
										assign node369 = (inp[0]) ? 3'b000 : node370;
											assign node370 = (inp[4]) ? 3'b010 : 3'b000;
									assign node374 = (inp[4]) ? node382 : node375;
										assign node375 = (inp[0]) ? node379 : node376;
											assign node376 = (inp[3]) ? 3'b000 : 3'b010;
											assign node379 = (inp[3]) ? 3'b110 : 3'b100;
										assign node382 = (inp[0]) ? node384 : 3'b100;
											assign node384 = (inp[3]) ? 3'b000 : 3'b010;
								assign node387 = (inp[4]) ? 3'b010 : node388;
									assign node388 = (inp[0]) ? node394 : node389;
										assign node389 = (inp[3]) ? 3'b110 : node390;
											assign node390 = (inp[8]) ? 3'b110 : 3'b010;
										assign node394 = (inp[3]) ? node396 : 3'b010;
											assign node396 = (inp[8]) ? 3'b110 : 3'b010;
						assign node400 = (inp[4]) ? node450 : node401;
							assign node401 = (inp[5]) ? node439 : node402;
								assign node402 = (inp[3]) ? node428 : node403;
									assign node403 = (inp[11]) ? node413 : node404;
										assign node404 = (inp[0]) ? node410 : node405;
											assign node405 = (inp[8]) ? 3'b010 : node406;
												assign node406 = (inp[6]) ? 3'b010 : 3'b000;
											assign node410 = (inp[8]) ? 3'b000 : 3'b010;
										assign node413 = (inp[6]) ? node421 : node414;
											assign node414 = (inp[0]) ? node418 : node415;
												assign node415 = (inp[8]) ? 3'b000 : 3'b010;
												assign node418 = (inp[8]) ? 3'b010 : 3'b000;
											assign node421 = (inp[0]) ? node425 : node422;
												assign node422 = (inp[8]) ? 3'b000 : 3'b010;
												assign node425 = (inp[8]) ? 3'b010 : 3'b000;
									assign node428 = (inp[0]) ? node430 : 3'b000;
										assign node430 = (inp[8]) ? node434 : node431;
											assign node431 = (inp[11]) ? 3'b010 : 3'b000;
											assign node434 = (inp[11]) ? 3'b000 : node435;
												assign node435 = (inp[6]) ? 3'b010 : 3'b000;
								assign node439 = (inp[11]) ? 3'b010 : node440;
									assign node440 = (inp[0]) ? 3'b000 : node441;
										assign node441 = (inp[3]) ? 3'b010 : node442;
											assign node442 = (inp[8]) ? node444 : 3'b010;
												assign node444 = (inp[6]) ? 3'b010 : 3'b000;
							assign node450 = (inp[5]) ? 3'b000 : node451;
								assign node451 = (inp[11]) ? 3'b000 : node452;
									assign node452 = (inp[8]) ? node458 : node453;
										assign node453 = (inp[6]) ? 3'b010 : node454;
											assign node454 = (inp[0]) ? 3'b000 : 3'b010;
										assign node458 = (inp[6]) ? 3'b000 : node459;
											assign node459 = (inp[3]) ? node461 : 3'b000;
												assign node461 = (inp[0]) ? 3'b010 : 3'b000;
			assign node467 = (inp[2]) ? node573 : node468;
				assign node468 = (inp[0]) ? 3'b010 : node469;
					assign node469 = (inp[1]) ? node493 : node470;
						assign node470 = (inp[7]) ? node472 : 3'b011;
							assign node472 = (inp[3]) ? 3'b011 : node473;
								assign node473 = (inp[8]) ? node487 : node474;
									assign node474 = (inp[5]) ? node482 : node475;
										assign node475 = (inp[11]) ? 3'b000 : node476;
											assign node476 = (inp[4]) ? node478 : 3'b011;
												assign node478 = (inp[6]) ? 3'b010 : 3'b000;
										assign node482 = (inp[6]) ? node484 : 3'b010;
											assign node484 = (inp[11]) ? 3'b010 : 3'b000;
									assign node487 = (inp[4]) ? node489 : 3'b011;
										assign node489 = (inp[11]) ? 3'b010 : 3'b000;
						assign node493 = (inp[3]) ? node547 : node494;
							assign node494 = (inp[5]) ? node526 : node495;
								assign node495 = (inp[6]) ? node507 : node496;
									assign node496 = (inp[7]) ? node502 : node497;
										assign node497 = (inp[4]) ? 3'b100 : node498;
											assign node498 = (inp[8]) ? 3'b000 : 3'b100;
										assign node502 = (inp[8]) ? node504 : 3'b000;
											assign node504 = (inp[4]) ? 3'b000 : 3'b100;
									assign node507 = (inp[11]) ? node519 : node508;
										assign node508 = (inp[7]) ? node514 : node509;
											assign node509 = (inp[4]) ? node511 : 3'b010;
												assign node511 = (inp[8]) ? 3'b010 : 3'b110;
											assign node514 = (inp[8]) ? 3'b110 : node515;
												assign node515 = (inp[4]) ? 3'b010 : 3'b110;
										assign node519 = (inp[7]) ? 3'b000 : node520;
											assign node520 = (inp[8]) ? node522 : 3'b100;
												assign node522 = (inp[4]) ? 3'b100 : 3'b000;
								assign node526 = (inp[7]) ? node536 : node527;
									assign node527 = (inp[11]) ? node531 : node528;
										assign node528 = (inp[6]) ? 3'b100 : 3'b110;
										assign node531 = (inp[4]) ? 3'b110 : node532;
											assign node532 = (inp[8]) ? 3'b010 : 3'b110;
									assign node536 = (inp[6]) ? node542 : node537;
										assign node537 = (inp[4]) ? 3'b010 : node538;
											assign node538 = (inp[8]) ? 3'b110 : 3'b010;
										assign node542 = (inp[11]) ? 3'b010 : node543;
											assign node543 = (inp[4]) ? 3'b000 : 3'b100;
							assign node547 = (inp[7]) ? node549 : 3'b011;
								assign node549 = (inp[4]) ? node559 : node550;
									assign node550 = (inp[8]) ? 3'b011 : node551;
										assign node551 = (inp[11]) ? node555 : node552;
											assign node552 = (inp[5]) ? 3'b000 : 3'b011;
											assign node555 = (inp[5]) ? 3'b010 : 3'b000;
									assign node559 = (inp[5]) ? node567 : node560;
										assign node560 = (inp[6]) ? node562 : 3'b000;
											assign node562 = (inp[11]) ? 3'b000 : node563;
												assign node563 = (inp[8]) ? 3'b011 : 3'b010;
										assign node567 = (inp[6]) ? node569 : 3'b010;
											assign node569 = (inp[11]) ? 3'b010 : 3'b000;
				assign node573 = (inp[0]) ? node787 : node574;
					assign node574 = (inp[1]) ? node686 : node575;
						assign node575 = (inp[11]) ? node643 : node576;
							assign node576 = (inp[3]) ? node604 : node577;
								assign node577 = (inp[7]) ? node593 : node578;
									assign node578 = (inp[8]) ? node582 : node579;
										assign node579 = (inp[4]) ? 3'b000 : 3'b100;
										assign node582 = (inp[4]) ? node590 : node583;
											assign node583 = (inp[6]) ? node587 : node584;
												assign node584 = (inp[5]) ? 3'b010 : 3'b000;
												assign node587 = (inp[5]) ? 3'b000 : 3'b010;
											assign node590 = (inp[5]) ? 3'b000 : 3'b100;
									assign node593 = (inp[4]) ? node599 : node594;
										assign node594 = (inp[8]) ? node596 : 3'b100;
											assign node596 = (inp[5]) ? 3'b100 : 3'b000;
										assign node599 = (inp[5]) ? node601 : 3'b100;
											assign node601 = (inp[6]) ? 3'b010 : 3'b000;
								assign node604 = (inp[7]) ? node626 : node605;
									assign node605 = (inp[4]) ? node619 : node606;
										assign node606 = (inp[8]) ? node614 : node607;
											assign node607 = (inp[6]) ? node611 : node608;
												assign node608 = (inp[5]) ? 3'b110 : 3'b100;
												assign node611 = (inp[5]) ? 3'b100 : 3'b010;
											assign node614 = (inp[6]) ? 3'b000 : node615;
												assign node615 = (inp[5]) ? 3'b010 : 3'b000;
										assign node619 = (inp[6]) ? node623 : node620;
											assign node620 = (inp[5]) ? 3'b110 : 3'b100;
											assign node623 = (inp[5]) ? 3'b100 : 3'b110;
									assign node626 = (inp[8]) ? node634 : node627;
										assign node627 = (inp[4]) ? 3'b000 : node628;
											assign node628 = (inp[5]) ? node630 : 3'b000;
												assign node630 = (inp[6]) ? 3'b000 : 3'b010;
										assign node634 = (inp[4]) ? node640 : node635;
											assign node635 = (inp[6]) ? 3'b100 : node636;
												assign node636 = (inp[5]) ? 3'b110 : 3'b100;
											assign node640 = (inp[5]) ? 3'b000 : 3'b110;
							assign node643 = (inp[5]) ? node671 : node644;
								assign node644 = (inp[3]) ? node658 : node645;
									assign node645 = (inp[7]) ? node651 : node646;
										assign node646 = (inp[8]) ? node648 : 3'b010;
											assign node648 = (inp[4]) ? 3'b100 : 3'b000;
										assign node651 = (inp[8]) ? node655 : node652;
											assign node652 = (inp[4]) ? 3'b000 : 3'b110;
											assign node655 = (inp[4]) ? 3'b110 : 3'b010;
									assign node658 = (inp[7]) ? node664 : node659;
										assign node659 = (inp[8]) ? node661 : 3'b100;
											assign node661 = (inp[4]) ? 3'b100 : 3'b000;
										assign node664 = (inp[8]) ? node668 : node665;
											assign node665 = (inp[4]) ? 3'b010 : 3'b000;
											assign node668 = (inp[4]) ? 3'b000 : 3'b100;
								assign node671 = (inp[4]) ? node681 : node672;
									assign node672 = (inp[7]) ? node676 : node673;
										assign node673 = (inp[8]) ? 3'b010 : 3'b110;
										assign node676 = (inp[8]) ? 3'b110 : node677;
											assign node677 = (inp[3]) ? 3'b010 : 3'b110;
									assign node681 = (inp[3]) ? node683 : 3'b010;
										assign node683 = (inp[7]) ? 3'b010 : 3'b110;
						assign node686 = (inp[7]) ? node740 : node687;
							assign node687 = (inp[4]) ? node717 : node688;
								assign node688 = (inp[11]) ? node706 : node689;
									assign node689 = (inp[3]) ? node699 : node690;
										assign node690 = (inp[8]) ? node696 : node691;
											assign node691 = (inp[5]) ? 3'b010 : node692;
												assign node692 = (inp[6]) ? 3'b100 : 3'b110;
											assign node696 = (inp[5]) ? 3'b100 : 3'b000;
										assign node699 = (inp[6]) ? 3'b100 : node700;
											assign node700 = (inp[5]) ? node702 : 3'b000;
												assign node702 = (inp[8]) ? 3'b100 : 3'b000;
									assign node706 = (inp[5]) ? node712 : node707;
										assign node707 = (inp[3]) ? node709 : 3'b100;
											assign node709 = (inp[8]) ? 3'b010 : 3'b110;
										assign node712 = (inp[8]) ? node714 : 3'b010;
											assign node714 = (inp[3]) ? 3'b110 : 3'b010;
								assign node717 = (inp[5]) ? node733 : node718;
									assign node718 = (inp[11]) ? node728 : node719;
										assign node719 = (inp[6]) ? node725 : node720;
											assign node720 = (inp[8]) ? 3'b010 : node721;
												assign node721 = (inp[3]) ? 3'b010 : 3'b000;
											assign node725 = (inp[8]) ? 3'b010 : 3'b110;
										assign node728 = (inp[3]) ? node730 : 3'b000;
											assign node730 = (inp[8]) ? 3'b000 : 3'b100;
									assign node733 = (inp[11]) ? 3'b010 : node734;
										assign node734 = (inp[3]) ? 3'b010 : node735;
											assign node735 = (inp[8]) ? 3'b010 : 3'b000;
							assign node740 = (inp[4]) ? node774 : node741;
								assign node741 = (inp[11]) ? node757 : node742;
									assign node742 = (inp[5]) ? node750 : node743;
										assign node743 = (inp[3]) ? node747 : node744;
											assign node744 = (inp[6]) ? 3'b000 : 3'b010;
											assign node747 = (inp[6]) ? 3'b010 : 3'b000;
										assign node750 = (inp[8]) ? 3'b000 : node751;
											assign node751 = (inp[3]) ? node753 : 3'b000;
												assign node753 = (inp[6]) ? 3'b010 : 3'b000;
									assign node757 = (inp[5]) ? 3'b010 : node758;
										assign node758 = (inp[6]) ? node766 : node759;
											assign node759 = (inp[3]) ? node763 : node760;
												assign node760 = (inp[8]) ? 3'b010 : 3'b000;
												assign node763 = (inp[8]) ? 3'b000 : 3'b010;
											assign node766 = (inp[8]) ? node770 : node767;
												assign node767 = (inp[3]) ? 3'b010 : 3'b000;
												assign node770 = (inp[3]) ? 3'b000 : 3'b010;
								assign node774 = (inp[6]) ? node776 : 3'b000;
									assign node776 = (inp[5]) ? 3'b000 : node777;
										assign node777 = (inp[11]) ? 3'b000 : node778;
											assign node778 = (inp[3]) ? node782 : node779;
												assign node779 = (inp[8]) ? 3'b010 : 3'b000;
												assign node782 = (inp[8]) ? 3'b000 : 3'b010;
					assign node787 = (inp[1]) ? node807 : node788;
						assign node788 = (inp[7]) ? node790 : 3'b010;
							assign node790 = (inp[3]) ? 3'b010 : node791;
								assign node791 = (inp[5]) ? node801 : node792;
									assign node792 = (inp[6]) ? node798 : node793;
										assign node793 = (inp[4]) ? 3'b000 : node794;
											assign node794 = (inp[8]) ? 3'b010 : 3'b000;
										assign node798 = (inp[11]) ? 3'b000 : 3'b010;
									assign node801 = (inp[11]) ? 3'b010 : node802;
										assign node802 = (inp[6]) ? 3'b000 : 3'b010;
						assign node807 = (inp[7]) ? node841 : node808;
							assign node808 = (inp[3]) ? 3'b010 : node809;
								assign node809 = (inp[11]) ? node827 : node810;
									assign node810 = (inp[8]) ? node818 : node811;
										assign node811 = (inp[4]) ? 3'b000 : node812;
											assign node812 = (inp[5]) ? 3'b100 : node813;
												assign node813 = (inp[6]) ? 3'b010 : 3'b100;
										assign node818 = (inp[5]) ? node822 : node819;
											assign node819 = (inp[6]) ? 3'b010 : 3'b000;
											assign node822 = (inp[4]) ? 3'b000 : node823;
												assign node823 = (inp[6]) ? 3'b000 : 3'b010;
									assign node827 = (inp[5]) ? node835 : node828;
										assign node828 = (inp[4]) ? node832 : node829;
											assign node829 = (inp[8]) ? 3'b000 : 3'b100;
											assign node832 = (inp[8]) ? 3'b100 : 3'b010;
										assign node835 = (inp[8]) ? 3'b010 : node836;
											assign node836 = (inp[4]) ? 3'b010 : 3'b110;
							assign node841 = (inp[4]) ? node867 : node842;
								assign node842 = (inp[5]) ? node858 : node843;
									assign node843 = (inp[3]) ? node851 : node844;
										assign node844 = (inp[6]) ? 3'b000 : node845;
											assign node845 = (inp[8]) ? 3'b000 : node846;
												assign node846 = (inp[11]) ? 3'b000 : 3'b010;
										assign node851 = (inp[8]) ? 3'b010 : node852;
											assign node852 = (inp[6]) ? node854 : 3'b000;
												assign node854 = (inp[11]) ? 3'b000 : 3'b010;
									assign node858 = (inp[11]) ? 3'b010 : node859;
										assign node859 = (inp[6]) ? node861 : 3'b010;
											assign node861 = (inp[3]) ? node863 : 3'b010;
												assign node863 = (inp[8]) ? 3'b010 : 3'b000;
								assign node867 = (inp[5]) ? 3'b000 : node868;
									assign node868 = (inp[3]) ? node870 : 3'b000;
										assign node870 = (inp[6]) ? node872 : 3'b000;
											assign node872 = (inp[11]) ? 3'b000 : 3'b010;
		assign node876 = (inp[9]) ? node1364 : node877;
			assign node877 = (inp[2]) ? node1021 : node878;
				assign node878 = (inp[0]) ? 3'b100 : node879;
					assign node879 = (inp[1]) ? node929 : node880;
						assign node880 = (inp[3]) ? 3'b101 : node881;
							assign node881 = (inp[7]) ? node907 : node882;
								assign node882 = (inp[8]) ? node898 : node883;
									assign node883 = (inp[4]) ? node891 : node884;
										assign node884 = (inp[5]) ? node886 : 3'b101;
											assign node886 = (inp[11]) ? 3'b000 : node887;
												assign node887 = (inp[6]) ? 3'b101 : 3'b000;
										assign node891 = (inp[5]) ? node893 : 3'b010;
											assign node893 = (inp[6]) ? node895 : 3'b000;
												assign node895 = (inp[11]) ? 3'b000 : 3'b010;
									assign node898 = (inp[4]) ? node900 : 3'b101;
										assign node900 = (inp[5]) ? node902 : 3'b101;
											assign node902 = (inp[6]) ? node904 : 3'b000;
												assign node904 = (inp[11]) ? 3'b000 : 3'b101;
								assign node907 = (inp[5]) ? node915 : node908;
									assign node908 = (inp[4]) ? node910 : 3'b010;
										assign node910 = (inp[8]) ? 3'b010 : node911;
											assign node911 = (inp[11]) ? 3'b110 : 3'b100;
									assign node915 = (inp[11]) ? node923 : node916;
										assign node916 = (inp[6]) ? node918 : 3'b100;
											assign node918 = (inp[8]) ? 3'b010 : node919;
												assign node919 = (inp[4]) ? 3'b110 : 3'b010;
										assign node923 = (inp[8]) ? node925 : 3'b100;
											assign node925 = (inp[4]) ? 3'b100 : 3'b000;
						assign node929 = (inp[7]) ? node985 : node930;
							assign node930 = (inp[3]) ? node960 : node931;
								assign node931 = (inp[5]) ? node947 : node932;
									assign node932 = (inp[8]) ? node942 : node933;
										assign node933 = (inp[4]) ? node939 : node934;
											assign node934 = (inp[11]) ? 3'b110 : node935;
												assign node935 = (inp[6]) ? 3'b100 : 3'b110;
											assign node939 = (inp[11]) ? 3'b010 : 3'b000;
										assign node942 = (inp[6]) ? node944 : 3'b110;
											assign node944 = (inp[11]) ? 3'b110 : 3'b100;
									assign node947 = (inp[4]) ? node953 : node948;
										assign node948 = (inp[6]) ? node950 : 3'b100;
											assign node950 = (inp[11]) ? 3'b000 : 3'b110;
										assign node953 = (inp[6]) ? node955 : 3'b000;
											assign node955 = (inp[11]) ? 3'b000 : node956;
												assign node956 = (inp[8]) ? 3'b110 : 3'b010;
								assign node960 = (inp[5]) ? node968 : node961;
									assign node961 = (inp[8]) ? 3'b101 : node962;
										assign node962 = (inp[4]) ? node964 : 3'b101;
											assign node964 = (inp[11]) ? 3'b010 : 3'b000;
									assign node968 = (inp[4]) ? node974 : node969;
										assign node969 = (inp[8]) ? 3'b101 : node970;
											assign node970 = (inp[6]) ? 3'b101 : 3'b000;
										assign node974 = (inp[8]) ? node980 : node975;
											assign node975 = (inp[6]) ? node977 : 3'b000;
												assign node977 = (inp[11]) ? 3'b000 : 3'b010;
											assign node980 = (inp[11]) ? 3'b000 : node981;
												assign node981 = (inp[6]) ? 3'b101 : 3'b000;
							assign node985 = (inp[5]) ? node1003 : node986;
								assign node986 = (inp[11]) ? node998 : node987;
									assign node987 = (inp[6]) ? node993 : node988;
										assign node988 = (inp[8]) ? 3'b010 : node989;
											assign node989 = (inp[4]) ? 3'b110 : 3'b010;
										assign node993 = (inp[8]) ? 3'b000 : node994;
											assign node994 = (inp[4]) ? 3'b100 : 3'b000;
									assign node998 = (inp[8]) ? 3'b010 : node999;
										assign node999 = (inp[4]) ? 3'b110 : 3'b010;
								assign node1003 = (inp[6]) ? node1009 : node1004;
									assign node1004 = (inp[4]) ? 3'b100 : node1005;
										assign node1005 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1009 = (inp[11]) ? node1015 : node1010;
										assign node1010 = (inp[8]) ? 3'b010 : node1011;
											assign node1011 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1015 = (inp[4]) ? 3'b100 : node1016;
											assign node1016 = (inp[8]) ? 3'b000 : 3'b100;
				assign node1021 = (inp[1]) ? node1181 : node1022;
					assign node1022 = (inp[0]) ? node1138 : node1023;
						assign node1023 = (inp[11]) ? node1097 : node1024;
							assign node1024 = (inp[4]) ? node1056 : node1025;
								assign node1025 = (inp[3]) ? node1039 : node1026;
									assign node1026 = (inp[8]) ? node1032 : node1027;
										assign node1027 = (inp[5]) ? 3'b010 : node1028;
											assign node1028 = (inp[7]) ? 3'b110 : 3'b100;
										assign node1032 = (inp[5]) ? node1034 : 3'b110;
											assign node1034 = (inp[6]) ? 3'b110 : node1035;
												assign node1035 = (inp[7]) ? 3'b110 : 3'b100;
									assign node1039 = (inp[7]) ? node1049 : node1040;
										assign node1040 = (inp[5]) ? node1044 : node1041;
											assign node1041 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1044 = (inp[6]) ? 3'b110 : node1045;
												assign node1045 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1049 = (inp[5]) ? node1053 : node1050;
											assign node1050 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1053 = (inp[6]) ? 3'b010 : 3'b000;
								assign node1056 = (inp[5]) ? node1074 : node1057;
									assign node1057 = (inp[8]) ? node1067 : node1058;
										assign node1058 = (inp[6]) ? node1064 : node1059;
											assign node1059 = (inp[7]) ? node1061 : 3'b010;
												assign node1061 = (inp[3]) ? 3'b010 : 3'b000;
											assign node1064 = (inp[7]) ? 3'b010 : 3'b000;
										assign node1067 = (inp[7]) ? 3'b010 : node1068;
											assign node1068 = (inp[3]) ? node1070 : 3'b010;
												assign node1070 = (inp[6]) ? 3'b100 : 3'b110;
									assign node1074 = (inp[8]) ? node1084 : node1075;
										assign node1075 = (inp[7]) ? node1079 : node1076;
											assign node1076 = (inp[6]) ? 3'b110 : 3'b000;
											assign node1079 = (inp[3]) ? 3'b110 : node1080;
												assign node1080 = (inp[6]) ? 3'b100 : 3'b110;
										assign node1084 = (inp[6]) ? node1090 : node1085;
											assign node1085 = (inp[7]) ? 3'b010 : node1086;
												assign node1086 = (inp[3]) ? 3'b000 : 3'b010;
											assign node1090 = (inp[7]) ? node1094 : node1091;
												assign node1091 = (inp[3]) ? 3'b110 : 3'b010;
												assign node1094 = (inp[3]) ? 3'b010 : 3'b000;
							assign node1097 = (inp[5]) ? node1125 : node1098;
								assign node1098 = (inp[7]) ? node1112 : node1099;
									assign node1099 = (inp[3]) ? node1107 : node1100;
										assign node1100 = (inp[8]) ? node1104 : node1101;
											assign node1101 = (inp[4]) ? 3'b100 : 3'b000;
											assign node1104 = (inp[4]) ? 3'b000 : 3'b110;
										assign node1107 = (inp[8]) ? 3'b110 : node1108;
											assign node1108 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1112 = (inp[8]) ? node1120 : node1113;
										assign node1113 = (inp[3]) ? node1117 : node1114;
											assign node1114 = (inp[4]) ? 3'b010 : 3'b000;
											assign node1117 = (inp[4]) ? 3'b100 : 3'b000;
										assign node1120 = (inp[3]) ? node1122 : 3'b100;
											assign node1122 = (inp[4]) ? 3'b000 : 3'b010;
								assign node1125 = (inp[4]) ? node1133 : node1126;
									assign node1126 = (inp[7]) ? 3'b000 : node1127;
										assign node1127 = (inp[3]) ? node1129 : 3'b000;
											assign node1129 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1133 = (inp[7]) ? 3'b100 : node1134;
										assign node1134 = (inp[3]) ? 3'b000 : 3'b100;
						assign node1138 = (inp[3]) ? 3'b100 : node1139;
							assign node1139 = (inp[5]) ? node1159 : node1140;
								assign node1140 = (inp[7]) ? node1150 : node1141;
									assign node1141 = (inp[8]) ? 3'b100 : node1142;
										assign node1142 = (inp[4]) ? node1144 : 3'b100;
											assign node1144 = (inp[11]) ? 3'b010 : node1145;
												assign node1145 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1150 = (inp[11]) ? node1154 : node1151;
										assign node1151 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1154 = (inp[8]) ? 3'b010 : node1155;
											assign node1155 = (inp[4]) ? 3'b110 : 3'b010;
								assign node1159 = (inp[7]) ? node1171 : node1160;
									assign node1160 = (inp[4]) ? node1164 : node1161;
										assign node1161 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1164 = (inp[11]) ? 3'b000 : node1165;
											assign node1165 = (inp[6]) ? node1167 : 3'b000;
												assign node1167 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1171 = (inp[11]) ? node1175 : node1172;
										assign node1172 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1175 = (inp[4]) ? 3'b100 : node1176;
											assign node1176 = (inp[8]) ? 3'b000 : 3'b100;
					assign node1181 = (inp[7]) ? node1293 : node1182;
						assign node1182 = (inp[4]) ? node1244 : node1183;
							assign node1183 = (inp[11]) ? node1215 : node1184;
								assign node1184 = (inp[8]) ? node1202 : node1185;
									assign node1185 = (inp[5]) ? node1195 : node1186;
										assign node1186 = (inp[0]) ? node1190 : node1187;
											assign node1187 = (inp[6]) ? 3'b110 : 3'b000;
											assign node1190 = (inp[6]) ? 3'b100 : node1191;
												assign node1191 = (inp[3]) ? 3'b100 : 3'b110;
										assign node1195 = (inp[0]) ? 3'b010 : node1196;
											assign node1196 = (inp[3]) ? node1198 : 3'b100;
												assign node1198 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1202 = (inp[0]) ? node1206 : node1203;
										assign node1203 = (inp[5]) ? 3'b000 : 3'b110;
										assign node1206 = (inp[3]) ? 3'b100 : node1207;
											assign node1207 = (inp[6]) ? node1211 : node1208;
												assign node1208 = (inp[5]) ? 3'b100 : 3'b110;
												assign node1211 = (inp[5]) ? 3'b110 : 3'b100;
								assign node1215 = (inp[3]) ? node1225 : node1216;
									assign node1216 = (inp[8]) ? node1218 : 3'b000;
										assign node1218 = (inp[5]) ? node1222 : node1219;
											assign node1219 = (inp[0]) ? 3'b110 : 3'b000;
											assign node1222 = (inp[0]) ? 3'b000 : 3'b100;
									assign node1225 = (inp[5]) ? node1231 : node1226;
										assign node1226 = (inp[8]) ? 3'b100 : node1227;
											assign node1227 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1231 = (inp[6]) ? node1237 : node1232;
											assign node1232 = (inp[8]) ? 3'b100 : node1233;
												assign node1233 = (inp[0]) ? 3'b000 : 3'b100;
											assign node1237 = (inp[8]) ? node1241 : node1238;
												assign node1238 = (inp[0]) ? 3'b000 : 3'b100;
												assign node1241 = (inp[0]) ? 3'b100 : 3'b000;
							assign node1244 = (inp[3]) ? node1262 : node1245;
								assign node1245 = (inp[11]) ? node1255 : node1246;
									assign node1246 = (inp[6]) ? node1248 : 3'b010;
										assign node1248 = (inp[8]) ? 3'b010 : node1249;
											assign node1249 = (inp[5]) ? 3'b010 : node1250;
												assign node1250 = (inp[0]) ? 3'b010 : 3'b000;
									assign node1255 = (inp[5]) ? 3'b000 : node1256;
										assign node1256 = (inp[0]) ? 3'b000 : node1257;
											assign node1257 = (inp[8]) ? 3'b010 : 3'b000;
								assign node1262 = (inp[8]) ? node1282 : node1263;
									assign node1263 = (inp[0]) ? node1271 : node1264;
										assign node1264 = (inp[6]) ? node1266 : 3'b000;
											assign node1266 = (inp[11]) ? 3'b000 : node1267;
												assign node1267 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1271 = (inp[5]) ? node1277 : node1272;
											assign node1272 = (inp[11]) ? 3'b010 : node1273;
												assign node1273 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1277 = (inp[6]) ? node1279 : 3'b000;
												assign node1279 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1282 = (inp[0]) ? node1288 : node1283;
										assign node1283 = (inp[11]) ? 3'b000 : node1284;
											assign node1284 = (inp[6]) ? 3'b010 : 3'b100;
										assign node1288 = (inp[5]) ? node1290 : 3'b100;
											assign node1290 = (inp[6]) ? 3'b100 : 3'b000;
						assign node1293 = (inp[5]) ? node1347 : node1294;
							assign node1294 = (inp[4]) ? node1322 : node1295;
								assign node1295 = (inp[11]) ? node1311 : node1296;
									assign node1296 = (inp[0]) ? node1298 : 3'b000;
										assign node1298 = (inp[8]) ? node1304 : node1299;
											assign node1299 = (inp[3]) ? node1301 : 3'b000;
												assign node1301 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1304 = (inp[3]) ? node1308 : node1305;
												assign node1305 = (inp[6]) ? 3'b010 : 3'b000;
												assign node1308 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1311 = (inp[8]) ? node1317 : node1312;
										assign node1312 = (inp[3]) ? node1314 : 3'b000;
											assign node1314 = (inp[0]) ? 3'b000 : 3'b010;
										assign node1317 = (inp[3]) ? node1319 : 3'b010;
											assign node1319 = (inp[0]) ? 3'b010 : 3'b000;
								assign node1322 = (inp[11]) ? 3'b000 : node1323;
									assign node1323 = (inp[8]) ? node1335 : node1324;
										assign node1324 = (inp[0]) ? node1330 : node1325;
											assign node1325 = (inp[6]) ? node1327 : 3'b000;
												assign node1327 = (inp[3]) ? 3'b010 : 3'b000;
											assign node1330 = (inp[3]) ? 3'b000 : node1331;
												assign node1331 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1335 = (inp[3]) ? node1341 : node1336;
											assign node1336 = (inp[0]) ? 3'b000 : node1337;
												assign node1337 = (inp[6]) ? 3'b010 : 3'b000;
											assign node1341 = (inp[0]) ? node1343 : 3'b010;
												assign node1343 = (inp[6]) ? 3'b010 : 3'b000;
							assign node1347 = (inp[11]) ? 3'b000 : node1348;
								assign node1348 = (inp[4]) ? 3'b000 : node1349;
									assign node1349 = (inp[0]) ? node1355 : node1350;
										assign node1350 = (inp[3]) ? 3'b000 : node1351;
											assign node1351 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1355 = (inp[3]) ? 3'b010 : node1356;
											assign node1356 = (inp[8]) ? 3'b000 : node1357;
												assign node1357 = (inp[6]) ? 3'b010 : 3'b000;
			assign node1364 = (inp[0]) ? node1642 : node1365;
				assign node1365 = (inp[2]) ? node1455 : node1366;
					assign node1366 = (inp[3]) ? node1432 : node1367;
						assign node1367 = (inp[1]) ? node1383 : node1368;
							assign node1368 = (inp[7]) ? node1370 : 3'b001;
								assign node1370 = (inp[4]) ? node1372 : 3'b001;
									assign node1372 = (inp[8]) ? node1376 : node1373;
										assign node1373 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1376 = (inp[5]) ? node1378 : 3'b001;
											assign node1378 = (inp[11]) ? 3'b000 : node1379;
												assign node1379 = (inp[6]) ? 3'b001 : 3'b000;
							assign node1383 = (inp[5]) ? node1407 : node1384;
								assign node1384 = (inp[11]) ? node1396 : node1385;
									assign node1385 = (inp[6]) ? node1391 : node1386;
										assign node1386 = (inp[7]) ? 3'b110 : node1387;
											assign node1387 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1391 = (inp[7]) ? node1393 : 3'b000;
											assign node1393 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1396 = (inp[7]) ? node1402 : node1397;
										assign node1397 = (inp[4]) ? node1399 : 3'b010;
											assign node1399 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1402 = (inp[4]) ? node1404 : 3'b110;
											assign node1404 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1407 = (inp[6]) ? node1419 : node1408;
									assign node1408 = (inp[7]) ? node1414 : node1409;
										assign node1409 = (inp[11]) ? node1411 : 3'b100;
											assign node1411 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1414 = (inp[8]) ? node1416 : 3'b000;
											assign node1416 = (inp[4]) ? 3'b000 : 3'b100;
									assign node1419 = (inp[11]) ? node1427 : node1420;
										assign node1420 = (inp[7]) ? 3'b110 : node1421;
											assign node1421 = (inp[8]) ? 3'b010 : node1422;
												assign node1422 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1427 = (inp[7]) ? 3'b000 : node1428;
											assign node1428 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1432 = (inp[7]) ? node1434 : 3'b001;
							assign node1434 = (inp[1]) ? node1436 : 3'b001;
								assign node1436 = (inp[8]) ? node1450 : node1437;
									assign node1437 = (inp[4]) ? node1441 : node1438;
										assign node1438 = (inp[5]) ? 3'b000 : 3'b001;
										assign node1441 = (inp[5]) ? node1447 : node1442;
											assign node1442 = (inp[6]) ? node1444 : 3'b010;
												assign node1444 = (inp[11]) ? 3'b010 : 3'b000;
											assign node1447 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1450 = (inp[5]) ? node1452 : 3'b001;
										assign node1452 = (inp[6]) ? 3'b000 : 3'b001;
					assign node1455 = (inp[1]) ? node1539 : node1456;
						assign node1456 = (inp[5]) ? node1496 : node1457;
							assign node1457 = (inp[7]) ? node1477 : node1458;
								assign node1458 = (inp[11]) ? node1470 : node1459;
									assign node1459 = (inp[6]) ? node1465 : node1460;
										assign node1460 = (inp[4]) ? node1462 : 3'b010;
											assign node1462 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1465 = (inp[8]) ? 3'b000 : node1466;
											assign node1466 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1470 = (inp[8]) ? 3'b010 : node1471;
										assign node1471 = (inp[3]) ? 3'b110 : node1472;
											assign node1472 = (inp[4]) ? 3'b000 : 3'b010;
								assign node1477 = (inp[3]) ? node1489 : node1478;
									assign node1478 = (inp[11]) ? node1482 : node1479;
										assign node1479 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1482 = (inp[8]) ? node1486 : node1483;
											assign node1483 = (inp[4]) ? 3'b000 : 3'b100;
											assign node1486 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1489 = (inp[6]) ? node1491 : 3'b110;
										assign node1491 = (inp[4]) ? 3'b000 : node1492;
											assign node1492 = (inp[11]) ? 3'b110 : 3'b100;
							assign node1496 = (inp[11]) ? node1528 : node1497;
								assign node1497 = (inp[6]) ? node1517 : node1498;
									assign node1498 = (inp[7]) ? node1506 : node1499;
										assign node1499 = (inp[3]) ? 3'b100 : node1500;
											assign node1500 = (inp[4]) ? 3'b010 : node1501;
												assign node1501 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1506 = (inp[3]) ? node1512 : node1507;
											assign node1507 = (inp[4]) ? node1509 : 3'b110;
												assign node1509 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1512 = (inp[8]) ? 3'b000 : node1513;
												assign node1513 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1517 = (inp[7]) ? node1523 : node1518;
										assign node1518 = (inp[3]) ? node1520 : 3'b010;
											assign node1520 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1523 = (inp[3]) ? node1525 : 3'b110;
											assign node1525 = (inp[4]) ? 3'b010 : 3'b110;
								assign node1528 = (inp[4]) ? node1534 : node1529;
									assign node1529 = (inp[8]) ? node1531 : 3'b100;
										assign node1531 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1534 = (inp[3]) ? node1536 : 3'b000;
										assign node1536 = (inp[7]) ? 3'b000 : 3'b100;
						assign node1539 = (inp[7]) ? node1609 : node1540;
							assign node1540 = (inp[5]) ? node1580 : node1541;
								assign node1541 = (inp[6]) ? node1561 : node1542;
									assign node1542 = (inp[11]) ? node1548 : node1543;
										assign node1543 = (inp[4]) ? 3'b000 : node1544;
											assign node1544 = (inp[3]) ? 3'b010 : 3'b000;
										assign node1548 = (inp[8]) ? node1554 : node1549;
											assign node1549 = (inp[4]) ? 3'b010 : node1550;
												assign node1550 = (inp[3]) ? 3'b100 : 3'b110;
											assign node1554 = (inp[4]) ? node1558 : node1555;
												assign node1555 = (inp[3]) ? 3'b000 : 3'b010;
												assign node1558 = (inp[3]) ? 3'b010 : 3'b100;
									assign node1561 = (inp[11]) ? node1567 : node1562;
										assign node1562 = (inp[4]) ? node1564 : 3'b010;
											assign node1564 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1567 = (inp[3]) ? node1575 : node1568;
											assign node1568 = (inp[8]) ? node1572 : node1569;
												assign node1569 = (inp[4]) ? 3'b010 : 3'b110;
												assign node1572 = (inp[4]) ? 3'b100 : 3'b010;
											assign node1575 = (inp[8]) ? node1577 : 3'b100;
												assign node1577 = (inp[4]) ? 3'b010 : 3'b000;
								assign node1580 = (inp[11]) ? node1602 : node1581;
									assign node1581 = (inp[4]) ? node1591 : node1582;
										assign node1582 = (inp[3]) ? node1588 : node1583;
											assign node1583 = (inp[8]) ? node1585 : 3'b000;
												assign node1585 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1588 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1591 = (inp[8]) ? node1597 : node1592;
											assign node1592 = (inp[6]) ? 3'b010 : node1593;
												assign node1593 = (inp[3]) ? 3'b000 : 3'b100;
											assign node1597 = (inp[3]) ? node1599 : 3'b000;
												assign node1599 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1602 = (inp[3]) ? node1604 : 3'b000;
										assign node1604 = (inp[4]) ? 3'b000 : node1605;
											assign node1605 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1609 = (inp[4]) ? node1631 : node1610;
								assign node1610 = (inp[11]) ? node1624 : node1611;
									assign node1611 = (inp[6]) ? node1619 : node1612;
										assign node1612 = (inp[5]) ? 3'b010 : node1613;
											assign node1613 = (inp[8]) ? 3'b000 : node1614;
												assign node1614 = (inp[3]) ? 3'b010 : 3'b000;
										assign node1619 = (inp[3]) ? node1621 : 3'b010;
											assign node1621 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1624 = (inp[8]) ? node1626 : 3'b000;
										assign node1626 = (inp[3]) ? node1628 : 3'b000;
											assign node1628 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1631 = (inp[5]) ? 3'b000 : node1632;
									assign node1632 = (inp[11]) ? 3'b000 : node1633;
										assign node1633 = (inp[3]) ? node1635 : 3'b000;
											assign node1635 = (inp[8]) ? node1637 : 3'b000;
												assign node1637 = (inp[6]) ? 3'b010 : 3'b000;
				assign node1642 = (inp[2]) ? node1644 : 3'b000;
					assign node1644 = (inp[3]) ? node1696 : node1645;
						assign node1645 = (inp[1]) ? node1661 : node1646;
							assign node1646 = (inp[8]) ? 3'b000 : node1647;
								assign node1647 = (inp[4]) ? node1649 : 3'b000;
									assign node1649 = (inp[7]) ? node1651 : 3'b000;
										assign node1651 = (inp[5]) ? node1657 : node1652;
											assign node1652 = (inp[6]) ? node1654 : 3'b010;
												assign node1654 = (inp[11]) ? 3'b010 : 3'b000;
											assign node1657 = (inp[6]) ? 3'b010 : 3'b000;
							assign node1661 = (inp[5]) ? node1687 : node1662;
								assign node1662 = (inp[4]) ? node1670 : node1663;
									assign node1663 = (inp[11]) ? 3'b010 : node1664;
										assign node1664 = (inp[8]) ? 3'b010 : node1665;
											assign node1665 = (inp[7]) ? 3'b010 : 3'b000;
									assign node1670 = (inp[7]) ? node1682 : node1671;
										assign node1671 = (inp[8]) ? node1677 : node1672;
											assign node1672 = (inp[11]) ? 3'b000 : node1673;
												assign node1673 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1677 = (inp[6]) ? node1679 : 3'b010;
												assign node1679 = (inp[11]) ? 3'b010 : 3'b000;
										assign node1682 = (inp[8]) ? 3'b000 : node1683;
											assign node1683 = (inp[6]) ? 3'b010 : 3'b000;
								assign node1687 = (inp[6]) ? node1691 : node1688;
									assign node1688 = (inp[7]) ? 3'b000 : 3'b100;
									assign node1691 = (inp[7]) ? 3'b000 : node1692;
										assign node1692 = (inp[11]) ? 3'b000 : 3'b010;
						assign node1696 = (inp[1]) ? node1698 : 3'b000;
							assign node1698 = (inp[8]) ? 3'b000 : node1699;
								assign node1699 = (inp[5]) ? 3'b000 : node1700;
									assign node1700 = (inp[4]) ? node1702 : 3'b000;
										assign node1702 = (inp[11]) ? 3'b000 : node1703;
											assign node1703 = (inp[7]) ? 3'b010 : 3'b000;

endmodule