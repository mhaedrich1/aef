module dtc_split125_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node14;
	wire [4-1:0] node18;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node22;
	wire [4-1:0] node26;
	wire [4-1:0] node27;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node42;
	wire [4-1:0] node45;
	wire [4-1:0] node47;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node69;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node83;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node99;
	wire [4-1:0] node101;
	wire [4-1:0] node103;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node121;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node159;
	wire [4-1:0] node162;
	wire [4-1:0] node165;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node176;
	wire [4-1:0] node177;
	wire [4-1:0] node179;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node191;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node210;
	wire [4-1:0] node212;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node231;
	wire [4-1:0] node233;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node241;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node251;
	wire [4-1:0] node254;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node264;
	wire [4-1:0] node266;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node299;
	wire [4-1:0] node302;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node316;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node344;
	wire [4-1:0] node346;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node367;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node387;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node400;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node415;
	wire [4-1:0] node417;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node439;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node451;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node465;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node511;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node532;
	wire [4-1:0] node533;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node545;
	wire [4-1:0] node548;
	wire [4-1:0] node549;
	wire [4-1:0] node551;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node578;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node586;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node594;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node632;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node642;
	wire [4-1:0] node643;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node671;
	wire [4-1:0] node674;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node684;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node722;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node750;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node766;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node787;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node805;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node817;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node847;
	wire [4-1:0] node849;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node857;
	wire [4-1:0] node860;
	wire [4-1:0] node862;
	wire [4-1:0] node865;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node878;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node885;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node897;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node907;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node920;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node937;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node946;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node953;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node972;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node981;
	wire [4-1:0] node984;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node997;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1004;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1013;
	wire [4-1:0] node1015;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1033;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1065;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1077;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1086;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1099;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1110;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1126;
	wire [4-1:0] node1128;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1134;
	wire [4-1:0] node1137;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1143;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1164;
	wire [4-1:0] node1166;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1179;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1191;
	wire [4-1:0] node1193;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1206;
	wire [4-1:0] node1209;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1231;
	wire [4-1:0] node1233;
	wire [4-1:0] node1235;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1277;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1295;
	wire [4-1:0] node1298;
	wire [4-1:0] node1300;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1309;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1356;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1396;
	wire [4-1:0] node1398;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1405;
	wire [4-1:0] node1408;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1415;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1420;
	wire [4-1:0] node1424;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1448;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1485;
	wire [4-1:0] node1487;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1504;
	wire [4-1:0] node1506;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1513;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1519;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1526;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1547;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1555;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1562;
	wire [4-1:0] node1564;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1573;
	wire [4-1:0] node1575;
	wire [4-1:0] node1576;
	wire [4-1:0] node1578;
	wire [4-1:0] node1581;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1588;
	wire [4-1:0] node1590;
	wire [4-1:0] node1593;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1601;
	wire [4-1:0] node1604;
	wire [4-1:0] node1605;
	wire [4-1:0] node1608;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1620;
	wire [4-1:0] node1622;
	wire [4-1:0] node1624;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1633;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1639;
	wire [4-1:0] node1642;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1656;
	wire [4-1:0] node1658;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1670;
	wire [4-1:0] node1673;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1684;
	wire [4-1:0] node1686;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1698;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1728;
	wire [4-1:0] node1730;
	wire [4-1:0] node1733;
	wire [4-1:0] node1734;
	wire [4-1:0] node1736;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1746;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1754;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1769;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1785;
	wire [4-1:0] node1788;
	wire [4-1:0] node1789;
	wire [4-1:0] node1793;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1804;
	wire [4-1:0] node1807;
	wire [4-1:0] node1810;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1818;
	wire [4-1:0] node1822;
	wire [4-1:0] node1824;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1831;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1861;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1871;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1882;
	wire [4-1:0] node1883;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1890;
	wire [4-1:0] node1891;
	wire [4-1:0] node1894;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1904;
	wire [4-1:0] node1906;
	wire [4-1:0] node1909;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1916;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1923;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1936;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1952;
	wire [4-1:0] node1956;
	wire [4-1:0] node1958;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1968;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1997;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2015;
	wire [4-1:0] node2018;
	wire [4-1:0] node2019;
	wire [4-1:0] node2020;
	wire [4-1:0] node2022;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2039;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2053;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2067;
	wire [4-1:0] node2073;
	wire [4-1:0] node2075;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2093;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2113;
	wire [4-1:0] node2115;
	wire [4-1:0] node2118;
	wire [4-1:0] node2119;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2127;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2155;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2165;
	wire [4-1:0] node2169;
	wire [4-1:0] node2171;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2177;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2191;
	wire [4-1:0] node2192;
	wire [4-1:0] node2194;
	wire [4-1:0] node2197;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2207;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2219;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2228;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2233;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2271;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2280;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2292;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2300;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;
	wire [4-1:0] node2315;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2327;
	wire [4-1:0] node2328;
	wire [4-1:0] node2331;
	wire [4-1:0] node2334;
	wire [4-1:0] node2335;
	wire [4-1:0] node2338;
	wire [4-1:0] node2340;
	wire [4-1:0] node2343;
	wire [4-1:0] node2344;
	wire [4-1:0] node2345;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2358;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2365;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2390;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2397;
	wire [4-1:0] node2398;
	wire [4-1:0] node2399;
	wire [4-1:0] node2401;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2410;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2416;
	wire [4-1:0] node2417;
	wire [4-1:0] node2422;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2426;
	wire [4-1:0] node2427;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2439;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2450;
	wire [4-1:0] node2452;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2462;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2466;
	wire [4-1:0] node2470;
	wire [4-1:0] node2472;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2479;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2487;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2493;
	wire [4-1:0] node2496;
	wire [4-1:0] node2499;
	wire [4-1:0] node2501;
	wire [4-1:0] node2503;
	wire [4-1:0] node2504;
	wire [4-1:0] node2506;
	wire [4-1:0] node2507;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2514;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2529;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2538;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2543;
	wire [4-1:0] node2547;
	wire [4-1:0] node2548;
	wire [4-1:0] node2549;
	wire [4-1:0] node2550;
	wire [4-1:0] node2554;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2565;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2574;
	wire [4-1:0] node2576;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2584;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2591;
	wire [4-1:0] node2594;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2600;
	wire [4-1:0] node2603;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2611;
	wire [4-1:0] node2615;
	wire [4-1:0] node2617;
	wire [4-1:0] node2619;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2625;
	wire [4-1:0] node2628;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2634;
	wire [4-1:0] node2636;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2643;
	wire [4-1:0] node2645;
	wire [4-1:0] node2648;
	wire [4-1:0] node2649;
	wire [4-1:0] node2652;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2663;
	wire [4-1:0] node2666;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2673;
	wire [4-1:0] node2676;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2682;
	wire [4-1:0] node2685;
	wire [4-1:0] node2687;
	wire [4-1:0] node2689;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2694;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2700;
	wire [4-1:0] node2702;
	wire [4-1:0] node2705;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2710;
	wire [4-1:0] node2711;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2728;
	wire [4-1:0] node2729;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2743;
	wire [4-1:0] node2746;
	wire [4-1:0] node2747;
	wire [4-1:0] node2751;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2757;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2762;
	wire [4-1:0] node2763;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2769;
	wire [4-1:0] node2772;
	wire [4-1:0] node2774;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2792;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2801;
	wire [4-1:0] node2804;
	wire [4-1:0] node2805;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2810;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2819;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2836;
	wire [4-1:0] node2839;
	wire [4-1:0] node2841;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2847;
	wire [4-1:0] node2848;
	wire [4-1:0] node2849;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2858;
	wire [4-1:0] node2861;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2867;
	wire [4-1:0] node2868;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2874;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2882;
	wire [4-1:0] node2885;
	wire [4-1:0] node2887;
	wire [4-1:0] node2890;
	wire [4-1:0] node2891;
	wire [4-1:0] node2892;
	wire [4-1:0] node2894;
	wire [4-1:0] node2898;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2908;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2915;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2921;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2928;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2939;
	wire [4-1:0] node2940;
	wire [4-1:0] node2941;
	wire [4-1:0] node2944;
	wire [4-1:0] node2947;
	wire [4-1:0] node2948;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2967;
	wire [4-1:0] node2971;
	wire [4-1:0] node2972;
	wire [4-1:0] node2974;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2982;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2985;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2996;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3005;
	wire [4-1:0] node3008;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3012;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3020;
	wire [4-1:0] node3022;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3030;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3046;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3052;
	wire [4-1:0] node3053;
	wire [4-1:0] node3057;
	wire [4-1:0] node3060;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3063;
	wire [4-1:0] node3064;
	wire [4-1:0] node3068;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3073;
	wire [4-1:0] node3077;
	wire [4-1:0] node3080;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3096;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3104;
	wire [4-1:0] node3107;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3113;
	wire [4-1:0] node3116;
	wire [4-1:0] node3117;
	wire [4-1:0] node3119;
	wire [4-1:0] node3122;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3140;
	wire [4-1:0] node3141;
	wire [4-1:0] node3143;
	wire [4-1:0] node3146;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3155;
	wire [4-1:0] node3156;
	wire [4-1:0] node3157;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3173;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3181;
	wire [4-1:0] node3184;
	wire [4-1:0] node3187;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3198;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3204;
	wire [4-1:0] node3205;
	wire [4-1:0] node3208;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3216;
	wire [4-1:0] node3217;
	wire [4-1:0] node3219;
	wire [4-1:0] node3222;
	wire [4-1:0] node3224;
	wire [4-1:0] node3228;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3233;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3239;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3251;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3261;
	wire [4-1:0] node3264;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3281;
	wire [4-1:0] node3282;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3289;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3300;
	wire [4-1:0] node3301;
	wire [4-1:0] node3304;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3313;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3323;
	wire [4-1:0] node3327;
	wire [4-1:0] node3328;
	wire [4-1:0] node3331;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3338;
	wire [4-1:0] node3341;
	wire [4-1:0] node3343;
	wire [4-1:0] node3346;
	wire [4-1:0] node3347;
	wire [4-1:0] node3349;
	wire [4-1:0] node3352;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3357;
	wire [4-1:0] node3358;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3365;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3374;
	wire [4-1:0] node3377;
	wire [4-1:0] node3379;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3386;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3396;
	wire [4-1:0] node3400;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3405;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3413;
	wire [4-1:0] node3414;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3421;
	wire [4-1:0] node3422;
	wire [4-1:0] node3424;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3430;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3437;
	wire [4-1:0] node3438;
	wire [4-1:0] node3440;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3447;
	wire [4-1:0] node3450;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3465;
	wire [4-1:0] node3466;
	wire [4-1:0] node3467;
	wire [4-1:0] node3471;
	wire [4-1:0] node3474;
	wire [4-1:0] node3475;
	wire [4-1:0] node3478;
	wire [4-1:0] node3479;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3490;
	wire [4-1:0] node3493;
	wire [4-1:0] node3495;
	wire [4-1:0] node3497;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3506;
	wire [4-1:0] node3510;
	wire [4-1:0] node3511;
	wire [4-1:0] node3513;
	wire [4-1:0] node3516;
	wire [4-1:0] node3518;
	wire [4-1:0] node3521;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3529;
	wire [4-1:0] node3531;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3541;
	wire [4-1:0] node3543;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3554;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3569;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3576;
	wire [4-1:0] node3579;
	wire [4-1:0] node3580;
	wire [4-1:0] node3581;
	wire [4-1:0] node3582;
	wire [4-1:0] node3584;
	wire [4-1:0] node3587;
	wire [4-1:0] node3590;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3597;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3606;
	wire [4-1:0] node3609;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3622;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3630;
	wire [4-1:0] node3631;
	wire [4-1:0] node3632;
	wire [4-1:0] node3635;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3642;
	wire [4-1:0] node3643;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3650;
	wire [4-1:0] node3653;
	wire [4-1:0] node3654;
	wire [4-1:0] node3657;
	wire [4-1:0] node3660;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3668;
	wire [4-1:0] node3671;
	wire [4-1:0] node3673;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3695;
	wire [4-1:0] node3696;
	wire [4-1:0] node3697;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3707;
	wire [4-1:0] node3708;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3716;
	wire [4-1:0] node3717;
	wire [4-1:0] node3720;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3727;
	wire [4-1:0] node3729;
	wire [4-1:0] node3732;
	wire [4-1:0] node3733;
	wire [4-1:0] node3734;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3741;
	wire [4-1:0] node3745;
	wire [4-1:0] node3746;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3757;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3763;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3769;
	wire [4-1:0] node3771;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3779;
	wire [4-1:0] node3780;
	wire [4-1:0] node3786;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3791;
	wire [4-1:0] node3792;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3799;
	wire [4-1:0] node3801;
	wire [4-1:0] node3805;
	wire [4-1:0] node3806;
	wire [4-1:0] node3807;
	wire [4-1:0] node3808;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3817;
	wire [4-1:0] node3820;
	wire [4-1:0] node3822;
	wire [4-1:0] node3824;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3831;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3839;
	wire [4-1:0] node3840;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3847;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3854;
	wire [4-1:0] node3856;
	wire [4-1:0] node3859;
	wire [4-1:0] node3862;
	wire [4-1:0] node3863;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3870;
	wire [4-1:0] node3871;
	wire [4-1:0] node3874;
	wire [4-1:0] node3876;
	wire [4-1:0] node3879;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3892;
	wire [4-1:0] node3893;
	wire [4-1:0] node3897;
	wire [4-1:0] node3899;
	wire [4-1:0] node3900;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3910;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3917;
	wire [4-1:0] node3920;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3931;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3942;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3951;
	wire [4-1:0] node3953;
	wire [4-1:0] node3956;
	wire [4-1:0] node3958;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3978;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3988;
	wire [4-1:0] node3991;
	wire [4-1:0] node3992;
	wire [4-1:0] node3995;
	wire [4-1:0] node3998;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4007;
	wire [4-1:0] node4010;
	wire [4-1:0] node4012;
	wire [4-1:0] node4014;
	wire [4-1:0] node4017;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4020;
	wire [4-1:0] node4023;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4031;
	wire [4-1:0] node4033;
	wire [4-1:0] node4035;
	wire [4-1:0] node4038;
	wire [4-1:0] node4039;
	wire [4-1:0] node4040;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4049;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4054;
	wire [4-1:0] node4055;
	wire [4-1:0] node4058;
	wire [4-1:0] node4061;
	wire [4-1:0] node4063;
	wire [4-1:0] node4066;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4072;
	wire [4-1:0] node4074;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4080;
	wire [4-1:0] node4083;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4090;
	wire [4-1:0] node4091;
	wire [4-1:0] node4093;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4100;
	wire [4-1:0] node4102;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4108;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4115;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4122;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4130;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4144;
	wire [4-1:0] node4148;
	wire [4-1:0] node4151;
	wire [4-1:0] node4152;
	wire [4-1:0] node4154;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4160;
	wire [4-1:0] node4161;
	wire [4-1:0] node4165;
	wire [4-1:0] node4167;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4173;
	wire [4-1:0] node4176;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4191;
	wire [4-1:0] node4194;
	wire [4-1:0] node4195;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4203;
	wire [4-1:0] node4204;
	wire [4-1:0] node4205;
	wire [4-1:0] node4206;
	wire [4-1:0] node4211;
	wire [4-1:0] node4213;
	wire [4-1:0] node4216;
	wire [4-1:0] node4217;
	wire [4-1:0] node4218;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4222;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4240;
	wire [4-1:0] node4243;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4249;
	wire [4-1:0] node4253;
	wire [4-1:0] node4254;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4267;
	wire [4-1:0] node4270;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4274;
	wire [4-1:0] node4279;
	wire [4-1:0] node4281;
	wire [4-1:0] node4282;
	wire [4-1:0] node4283;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4290;
	wire [4-1:0] node4292;
	wire [4-1:0] node4295;
	wire [4-1:0] node4296;
	wire [4-1:0] node4298;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4306;
	wire [4-1:0] node4308;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4314;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4322;
	wire [4-1:0] node4325;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4329;
	wire [4-1:0] node4332;
	wire [4-1:0] node4334;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4341;
	wire [4-1:0] node4343;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4353;
	wire [4-1:0] node4357;
	wire [4-1:0] node4360;
	wire [4-1:0] node4361;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4371;
	wire [4-1:0] node4374;
	wire [4-1:0] node4375;
	wire [4-1:0] node4376;
	wire [4-1:0] node4378;
	wire [4-1:0] node4381;
	wire [4-1:0] node4382;
	wire [4-1:0] node4385;
	wire [4-1:0] node4388;
	wire [4-1:0] node4390;
	wire [4-1:0] node4392;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4406;
	wire [4-1:0] node4408;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4416;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4424;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4428;
	wire [4-1:0] node4432;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4439;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4445;
	wire [4-1:0] node4448;
	wire [4-1:0] node4449;
	wire [4-1:0] node4450;
	wire [4-1:0] node4454;
	wire [4-1:0] node4457;
	wire [4-1:0] node4458;
	wire [4-1:0] node4460;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4466;
	wire [4-1:0] node4467;
	wire [4-1:0] node4468;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4473;
	wire [4-1:0] node4474;
	wire [4-1:0] node4478;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4484;
	wire [4-1:0] node4487;
	wire [4-1:0] node4489;
	wire [4-1:0] node4492;
	wire [4-1:0] node4494;
	wire [4-1:0] node4496;
	wire [4-1:0] node4498;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4512;
	wire [4-1:0] node4515;
	wire [4-1:0] node4518;
	wire [4-1:0] node4519;
	wire [4-1:0] node4520;
	wire [4-1:0] node4524;
	wire [4-1:0] node4526;
	wire [4-1:0] node4528;
	wire [4-1:0] node4531;
	wire [4-1:0] node4532;
	wire [4-1:0] node4533;
	wire [4-1:0] node4534;
	wire [4-1:0] node4536;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4543;
	wire [4-1:0] node4546;
	wire [4-1:0] node4547;
	wire [4-1:0] node4550;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4555;
	wire [4-1:0] node4558;
	wire [4-1:0] node4559;
	wire [4-1:0] node4562;
	wire [4-1:0] node4565;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4571;
	wire [4-1:0] node4573;
	wire [4-1:0] node4576;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4582;
	wire [4-1:0] node4583;
	wire [4-1:0] node4585;
	wire [4-1:0] node4588;
	wire [4-1:0] node4590;
	wire [4-1:0] node4592;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4600;
	wire [4-1:0] node4601;
	wire [4-1:0] node4603;
	wire [4-1:0] node4606;
	wire [4-1:0] node4608;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4615;
	wire [4-1:0] node4616;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4623;
	wire [4-1:0] node4624;
	wire [4-1:0] node4627;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4633;
	wire [4-1:0] node4636;
	wire [4-1:0] node4639;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4646;
	wire [4-1:0] node4649;
	wire [4-1:0] node4651;
	wire [4-1:0] node4654;
	wire [4-1:0] node4656;
	wire [4-1:0] node4658;
	wire [4-1:0] node4661;
	wire [4-1:0] node4662;
	wire [4-1:0] node4664;
	wire [4-1:0] node4666;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4672;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4682;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4689;
	wire [4-1:0] node4692;
	wire [4-1:0] node4694;
	wire [4-1:0] node4696;
	wire [4-1:0] node4699;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4703;
	wire [4-1:0] node4707;
	wire [4-1:0] node4708;
	wire [4-1:0] node4709;
	wire [4-1:0] node4713;
	wire [4-1:0] node4714;
	wire [4-1:0] node4717;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4727;
	wire [4-1:0] node4731;
	wire [4-1:0] node4732;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4740;
	wire [4-1:0] node4743;
	wire [4-1:0] node4746;
	wire [4-1:0] node4747;
	wire [4-1:0] node4749;
	wire [4-1:0] node4752;
	wire [4-1:0] node4753;
	wire [4-1:0] node4756;
	wire [4-1:0] node4759;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4765;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4772;
	wire [4-1:0] node4776;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4784;
	wire [4-1:0] node4787;
	wire [4-1:0] node4790;
	wire [4-1:0] node4791;
	wire [4-1:0] node4792;
	wire [4-1:0] node4793;
	wire [4-1:0] node4795;
	wire [4-1:0] node4799;
	wire [4-1:0] node4800;
	wire [4-1:0] node4801;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4810;
	wire [4-1:0] node4811;
	wire [4-1:0] node4814;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4821;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4825;
	wire [4-1:0] node4830;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4836;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4842;
	wire [4-1:0] node4844;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4855;
	wire [4-1:0] node4856;
	wire [4-1:0] node4860;
	wire [4-1:0] node4863;
	wire [4-1:0] node4865;
	wire [4-1:0] node4868;
	wire [4-1:0] node4870;
	wire [4-1:0] node4871;
	wire [4-1:0] node4872;
	wire [4-1:0] node4874;
	wire [4-1:0] node4875;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4879;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4885;
	wire [4-1:0] node4888;
	wire [4-1:0] node4891;
	wire [4-1:0] node4893;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4899;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4902;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4923;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4929;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4934;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4944;
	wire [4-1:0] node4945;
	wire [4-1:0] node4949;
	wire [4-1:0] node4951;
	wire [4-1:0] node4954;
	wire [4-1:0] node4956;
	wire [4-1:0] node4958;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4963;
	wire [4-1:0] node4965;
	wire [4-1:0] node4968;
	wire [4-1:0] node4970;

	assign outp = (inp[8]) ? node2526 : node1;
		assign node1 = (inp[15]) ? node1427 : node2;
			assign node2 = (inp[6]) ? node404 : node3;
				assign node3 = (inp[9]) ? node195 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[5]) ? node73 : node6;
							assign node6 = (inp[2]) ? 4'b1111 : node7;
								assign node7 = (inp[3]) ? node35 : node8;
									assign node8 = (inp[4]) ? node18 : node9;
										assign node9 = (inp[7]) ? 4'b1111 : node10;
											assign node10 = (inp[10]) ? node14 : node11;
												assign node11 = (inp[11]) ? 4'b1111 : 4'b0001;
												assign node14 = (inp[13]) ? 4'b1000 : 4'b0001;
										assign node18 = (inp[1]) ? node26 : node19;
											assign node19 = (inp[7]) ? 4'b0000 : node20;
												assign node20 = (inp[12]) ? node22 : 4'b1000;
													assign node22 = (inp[10]) ? 4'b1000 : 4'b0001;
											assign node26 = (inp[13]) ? node32 : node27;
												assign node27 = (inp[12]) ? node29 : 4'b0001;
													assign node29 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node32 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node35 = (inp[13]) ? node55 : node36;
										assign node36 = (inp[4]) ? node50 : node37;
											assign node37 = (inp[7]) ? node45 : node38;
												assign node38 = (inp[1]) ? node42 : node39;
													assign node39 = (inp[12]) ? 4'b1001 : 4'b0100;
													assign node42 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node45 = (inp[1]) ? node47 : 4'b0000;
													assign node47 = (inp[11]) ? 4'b0001 : 4'b1000;
											assign node50 = (inp[1]) ? node52 : 4'b0100;
												assign node52 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node55 = (inp[10]) ? node63 : node56;
											assign node56 = (inp[12]) ? node58 : 4'b1001;
												assign node58 = (inp[14]) ? node60 : 4'b0101;
													assign node60 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node63 = (inp[7]) ? node69 : node64;
												assign node64 = (inp[1]) ? 4'b1101 : node65;
													assign node65 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node69 = (inp[1]) ? 4'b1101 : 4'b0001;
							assign node73 = (inp[1]) ? node135 : node74;
								assign node74 = (inp[3]) ? node106 : node75;
									assign node75 = (inp[4]) ? node91 : node76;
										assign node76 = (inp[2]) ? node86 : node77;
											assign node77 = (inp[7]) ? node79 : 4'b0000;
												assign node79 = (inp[12]) ? node83 : node80;
													assign node80 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node83 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node86 = (inp[7]) ? 4'b1111 : node87;
												assign node87 = (inp[13]) ? 4'b1000 : 4'b1111;
										assign node91 = (inp[11]) ? node99 : node92;
											assign node92 = (inp[14]) ? node94 : 4'b0000;
												assign node94 = (inp[10]) ? node96 : 4'b1101;
													assign node96 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node99 = (inp[7]) ? node101 : 4'b0000;
												assign node101 = (inp[14]) ? node103 : 4'b0000;
													assign node103 = (inp[2]) ? 4'b1111 : 4'b0000;
									assign node106 = (inp[4]) ? node124 : node107;
										assign node107 = (inp[7]) ? node115 : node108;
											assign node108 = (inp[12]) ? 4'b1001 : node109;
												assign node109 = (inp[13]) ? 4'b1100 : node110;
													assign node110 = (inp[11]) ? 4'b0100 : 4'b0100;
											assign node115 = (inp[10]) ? node121 : node116;
												assign node116 = (inp[11]) ? 4'b1000 : node117;
													assign node117 = (inp[13]) ? 4'b0001 : 4'b1000;
												assign node121 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node124 = (inp[13]) ? node132 : node125;
											assign node125 = (inp[12]) ? node127 : 4'b0100;
												assign node127 = (inp[10]) ? 4'b0100 : node128;
													assign node128 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node132 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node135 = (inp[3]) ? node165 : node136;
									assign node136 = (inp[13]) ? node150 : node137;
										assign node137 = (inp[7]) ? node145 : node138;
											assign node138 = (inp[12]) ? node140 : 4'b0001;
												assign node140 = (inp[10]) ? 4'b0000 : node141;
													assign node141 = (inp[4]) ? 4'b1000 : 4'b1111;
											assign node145 = (inp[2]) ? 4'b1111 : node146;
												assign node146 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node150 = (inp[12]) ? node156 : node151;
											assign node151 = (inp[11]) ? 4'b1001 : node152;
												assign node152 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node156 = (inp[11]) ? node162 : node157;
												assign node157 = (inp[4]) ? node159 : 4'b0100;
													assign node159 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node162 = (inp[4]) ? 4'b0001 : 4'b1001;
									assign node165 = (inp[2]) ? node187 : node166;
										assign node166 = (inp[13]) ? node176 : node167;
											assign node167 = (inp[12]) ? node173 : node168;
												assign node168 = (inp[7]) ? node170 : 4'b0100;
													assign node170 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node173 = (inp[10]) ? 4'b0101 : 4'b1001;
											assign node176 = (inp[10]) ? node182 : node177;
												assign node177 = (inp[12]) ? node179 : 4'b1101;
													assign node179 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node182 = (inp[11]) ? 4'b1101 : node183;
													assign node183 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node187 = (inp[7]) ? node191 : node188;
											assign node188 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node191 = (inp[4]) ? 4'b0101 : 4'b0001;
					assign node195 = (inp[0]) ? 4'b0101 : node196;
						assign node196 = (inp[5]) ? node258 : node197;
							assign node197 = (inp[2]) ? 4'b0111 : node198;
								assign node198 = (inp[3]) ? node222 : node199;
									assign node199 = (inp[7]) ? node215 : node200;
										assign node200 = (inp[4]) ? node204 : node201;
											assign node201 = (inp[1]) ? 4'b0001 : 4'b0111;
											assign node204 = (inp[13]) ? node210 : node205;
												assign node205 = (inp[1]) ? 4'b1001 : node206;
													assign node206 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node210 = (inp[1]) ? node212 : 4'b0000;
													assign node212 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node215 = (inp[13]) ? node217 : 4'b0111;
											assign node217 = (inp[10]) ? node219 : 4'b0111;
												assign node219 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node222 = (inp[4]) ? node236 : node223;
										assign node223 = (inp[10]) ? node231 : node224;
											assign node224 = (inp[13]) ? 4'b1001 : node225;
												assign node225 = (inp[12]) ? 4'b0001 : node226;
													assign node226 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node231 = (inp[1]) ? node233 : 4'b1000;
												assign node233 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node236 = (inp[13]) ? node246 : node237;
											assign node237 = (inp[7]) ? node241 : node238;
												assign node238 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node241 = (inp[14]) ? node243 : 4'b1000;
													assign node243 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node246 = (inp[10]) ? node254 : node247;
												assign node247 = (inp[12]) ? node251 : node248;
													assign node248 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node251 = (inp[7]) ? 4'b1001 : 4'b1100;
												assign node254 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node258 = (inp[1]) ? node316 : node259;
								assign node259 = (inp[13]) ? node291 : node260;
									assign node260 = (inp[10]) ? node278 : node261;
										assign node261 = (inp[3]) ? node269 : node262;
											assign node262 = (inp[2]) ? node264 : 4'b0101;
												assign node264 = (inp[4]) ? node266 : 4'b0111;
													assign node266 = (inp[7]) ? 4'b0111 : 4'b0000;
											assign node269 = (inp[14]) ? node273 : node270;
												assign node270 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node273 = (inp[11]) ? 4'b1100 : node274;
													assign node274 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node278 = (inp[3]) ? node286 : node279;
											assign node279 = (inp[2]) ? 4'b0111 : node280;
												assign node280 = (inp[4]) ? node282 : 4'b1100;
													assign node282 = (inp[7]) ? 4'b1100 : 4'b0000;
											assign node286 = (inp[7]) ? 4'b1000 : node287;
												assign node287 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node291 = (inp[10]) ? node305 : node292;
										assign node292 = (inp[12]) ? node302 : node293;
											assign node293 = (inp[4]) ? node299 : node294;
												assign node294 = (inp[11]) ? node296 : 4'b0100;
													assign node296 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node299 = (inp[3]) ? 4'b1001 : 4'b0000;
											assign node302 = (inp[7]) ? 4'b1100 : 4'b1000;
										assign node305 = (inp[3]) ? node311 : node306;
											assign node306 = (inp[7]) ? node308 : 4'b0000;
												assign node308 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node311 = (inp[4]) ? 4'b0100 : node312;
												assign node312 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node316 = (inp[13]) ? node360 : node317;
									assign node317 = (inp[12]) ? node337 : node318;
										assign node318 = (inp[11]) ? node326 : node319;
											assign node319 = (inp[14]) ? node323 : node320;
												assign node320 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node323 = (inp[3]) ? 4'b1000 : 4'b1100;
											assign node326 = (inp[3]) ? node332 : node327;
												assign node327 = (inp[14]) ? 4'b1001 : node328;
													assign node328 = (inp[2]) ? 4'b0111 : 4'b1101;
												assign node332 = (inp[4]) ? node334 : 4'b1001;
													assign node334 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node337 = (inp[10]) ? node349 : node338;
											assign node338 = (inp[3]) ? node344 : node339;
												assign node339 = (inp[2]) ? 4'b0111 : node340;
													assign node340 = (inp[4]) ? 4'b0000 : 4'b0101;
												assign node344 = (inp[4]) ? node346 : 4'b0001;
													assign node346 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node349 = (inp[2]) ? node357 : node350;
												assign node350 = (inp[11]) ? node354 : node351;
													assign node351 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node354 = (inp[14]) ? 4'b1001 : 4'b1001;
												assign node357 = (inp[7]) ? 4'b0111 : 4'b1001;
									assign node360 = (inp[10]) ? node390 : node361;
										assign node361 = (inp[12]) ? node377 : node362;
											assign node362 = (inp[14]) ? node370 : node363;
												assign node363 = (inp[2]) ? node367 : node364;
													assign node364 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node367 = (inp[3]) ? 4'b0001 : 4'b0111;
												assign node370 = (inp[3]) ? node374 : node371;
													assign node371 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node374 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node377 = (inp[3]) ? node383 : node378;
												assign node378 = (inp[2]) ? node380 : 4'b1101;
													assign node380 = (inp[4]) ? 4'b1000 : 4'b0111;
												assign node383 = (inp[14]) ? node387 : node384;
													assign node384 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node387 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node390 = (inp[3]) ? node400 : node391;
											assign node391 = (inp[4]) ? node395 : node392;
												assign node392 = (inp[7]) ? 4'b0111 : 4'b0001;
												assign node395 = (inp[7]) ? 4'b0001 : node396;
													assign node396 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node400 = (inp[4]) ? 4'b0101 : 4'b0001;
				assign node404 = (inp[5]) ? node888 : node405;
					assign node405 = (inp[0]) ? node733 : node406;
						assign node406 = (inp[11]) ? node570 : node407;
							assign node407 = (inp[2]) ? node485 : node408;
								assign node408 = (inp[3]) ? node446 : node409;
									assign node409 = (inp[4]) ? node431 : node410;
										assign node410 = (inp[13]) ? node420 : node411;
											assign node411 = (inp[12]) ? node415 : node412;
												assign node412 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node415 = (inp[9]) ? node417 : 4'b1101;
													assign node417 = (inp[14]) ? 4'b0000 : 4'b1100;
											assign node420 = (inp[1]) ? node426 : node421;
												assign node421 = (inp[10]) ? 4'b0000 : node422;
													assign node422 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node426 = (inp[14]) ? 4'b1000 : node427;
													assign node427 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node431 = (inp[7]) ? node439 : node432;
											assign node432 = (inp[9]) ? 4'b0100 : node433;
												assign node433 = (inp[10]) ? 4'b1100 : node434;
													assign node434 = (inp[1]) ? 4'b0100 : 4'b1100;
											assign node439 = (inp[13]) ? node441 : 4'b0000;
												assign node441 = (inp[12]) ? 4'b0100 : node442;
													assign node442 = (inp[9]) ? 4'b1000 : 4'b0100;
									assign node446 = (inp[4]) ? node468 : node447;
										assign node447 = (inp[7]) ? node459 : node448;
											assign node448 = (inp[10]) ? node454 : node449;
												assign node449 = (inp[13]) ? node451 : 4'b0000;
													assign node451 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node454 = (inp[9]) ? 4'b0000 : node455;
													assign node455 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node459 = (inp[10]) ? node463 : node460;
												assign node460 = (inp[9]) ? 4'b1100 : 4'b0100;
												assign node463 = (inp[13]) ? node465 : 4'b1100;
													assign node465 = (inp[9]) ? 4'b0000 : 4'b1000;
										assign node468 = (inp[13]) ? node474 : node469;
											assign node469 = (inp[1]) ? 4'b1000 : node470;
												assign node470 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node474 = (inp[7]) ? node480 : node475;
												assign node475 = (inp[10]) ? node477 : 4'b1101;
													assign node477 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node480 = (inp[10]) ? 4'b1001 : node481;
													assign node481 = (inp[14]) ? 4'b1001 : 4'b0100;
								assign node485 = (inp[3]) ? node537 : node486;
									assign node486 = (inp[7]) ? node514 : node487;
										assign node487 = (inp[10]) ? node499 : node488;
											assign node488 = (inp[4]) ? node496 : node489;
												assign node489 = (inp[1]) ? node493 : node490;
													assign node490 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node493 = (inp[14]) ? 4'b1000 : 4'b0001;
												assign node496 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node499 = (inp[14]) ? node507 : node500;
												assign node500 = (inp[9]) ? node504 : node501;
													assign node501 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node504 = (inp[12]) ? 4'b1100 : 4'b1101;
												assign node507 = (inp[1]) ? node511 : node508;
													assign node508 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node511 = (inp[9]) ? 4'b0000 : 4'b1000;
										assign node514 = (inp[4]) ? node526 : node515;
											assign node515 = (inp[12]) ? node519 : node516;
												assign node516 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node519 = (inp[1]) ? node523 : node520;
													assign node520 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node523 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node526 = (inp[14]) ? node532 : node527;
												assign node527 = (inp[12]) ? node529 : 4'b0001;
													assign node529 = (inp[9]) ? 4'b0001 : 4'b1001;
												assign node532 = (inp[13]) ? 4'b1000 : node533;
													assign node533 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node537 = (inp[4]) ? node559 : node538;
										assign node538 = (inp[7]) ? node548 : node539;
											assign node539 = (inp[12]) ? node541 : 4'b0000;
												assign node541 = (inp[13]) ? node545 : node542;
													assign node542 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node545 = (inp[9]) ? 4'b1000 : 4'b0000;
											assign node548 = (inp[13]) ? node554 : node549;
												assign node549 = (inp[9]) ? node551 : 4'b1001;
													assign node551 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node554 = (inp[9]) ? node556 : 4'b1000;
													assign node556 = (inp[14]) ? 4'b0000 : 4'b0000;
										assign node559 = (inp[10]) ? node565 : node560;
											assign node560 = (inp[12]) ? node562 : 4'b0100;
												assign node562 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node565 = (inp[7]) ? 4'b0100 : node566;
												assign node566 = (inp[12]) ? 4'b0100 : 4'b1100;
							assign node570 = (inp[1]) ? node654 : node571;
								assign node571 = (inp[3]) ? node613 : node572;
									assign node572 = (inp[2]) ? node594 : node573;
										assign node573 = (inp[4]) ? node581 : node574;
											assign node574 = (inp[10]) ? node578 : node575;
												assign node575 = (inp[7]) ? 4'b0100 : 4'b1100;
												assign node578 = (inp[12]) ? 4'b1100 : 4'b1001;
											assign node581 = (inp[13]) ? node589 : node582;
												assign node582 = (inp[9]) ? node586 : node583;
													assign node583 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node586 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node589 = (inp[7]) ? 4'b1001 : node590;
													assign node590 = (inp[14]) ? 4'b1101 : 4'b0101;
										assign node594 = (inp[7]) ? node604 : node595;
											assign node595 = (inp[9]) ? 4'b0000 : node596;
												assign node596 = (inp[14]) ? node600 : node597;
													assign node597 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node600 = (inp[13]) ? 4'b1000 : 4'b1000;
											assign node604 = (inp[4]) ? node610 : node605;
												assign node605 = (inp[9]) ? node607 : 4'b1100;
													assign node607 = (inp[14]) ? 4'b0100 : 4'b1100;
												assign node610 = (inp[14]) ? 4'b1100 : 4'b0000;
									assign node613 = (inp[2]) ? node635 : node614;
										assign node614 = (inp[4]) ? node624 : node615;
											assign node615 = (inp[9]) ? node619 : node616;
												assign node616 = (inp[12]) ? 4'b0001 : 4'b1000;
												assign node619 = (inp[10]) ? 4'b1101 : node620;
													assign node620 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node624 = (inp[7]) ? node628 : node625;
												assign node625 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node628 = (inp[13]) ? node632 : node629;
													assign node629 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node632 = (inp[9]) ? 4'b0000 : 4'b1000;
										assign node635 = (inp[9]) ? node647 : node636;
											assign node636 = (inp[4]) ? node642 : node637;
												assign node637 = (inp[10]) ? node639 : 4'b0000;
													assign node639 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node642 = (inp[13]) ? 4'b1101 : node643;
													assign node643 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node647 = (inp[10]) ? node651 : node648;
												assign node648 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node651 = (inp[4]) ? 4'b1001 : 4'b1000;
								assign node654 = (inp[4]) ? node696 : node655;
									assign node655 = (inp[7]) ? node677 : node656;
										assign node656 = (inp[13]) ? node668 : node657;
											assign node657 = (inp[2]) ? node663 : node658;
												assign node658 = (inp[12]) ? node660 : 4'b0001;
													assign node660 = (inp[10]) ? 4'b0001 : 4'b0001;
												assign node663 = (inp[9]) ? 4'b1101 : node664;
													assign node664 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node668 = (inp[2]) ? node674 : node669;
												assign node669 = (inp[9]) ? node671 : 4'b1001;
													assign node671 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node674 = (inp[3]) ? 4'b1001 : 4'b0001;
										assign node677 = (inp[13]) ? node687 : node678;
											assign node678 = (inp[3]) ? node684 : node679;
												assign node679 = (inp[9]) ? 4'b1101 : node680;
													assign node680 = (inp[2]) ? 4'b1101 : 4'b0101;
												assign node684 = (inp[2]) ? 4'b0001 : 4'b1101;
											assign node687 = (inp[3]) ? node691 : node688;
												assign node688 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node691 = (inp[10]) ? 4'b1001 : node692;
													assign node692 = (inp[2]) ? 4'b1001 : 4'b0001;
									assign node696 = (inp[13]) ? node716 : node697;
										assign node697 = (inp[12]) ? node705 : node698;
											assign node698 = (inp[7]) ? node700 : 4'b1001;
												assign node700 = (inp[10]) ? 4'b0001 : node701;
													assign node701 = (inp[3]) ? 4'b0001 : 4'b1001;
											assign node705 = (inp[3]) ? node713 : node706;
												assign node706 = (inp[9]) ? node710 : node707;
													assign node707 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node710 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node713 = (inp[10]) ? 4'b1101 : 4'b1001;
										assign node716 = (inp[3]) ? node730 : node717;
											assign node717 = (inp[2]) ? node725 : node718;
												assign node718 = (inp[7]) ? node722 : node719;
													assign node719 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node722 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node725 = (inp[12]) ? node727 : 4'b1001;
													assign node727 = (inp[9]) ? 4'b1001 : 4'b0001;
											assign node730 = (inp[9]) ? 4'b0101 : 4'b1101;
						assign node733 = (inp[2]) ? node885 : node734;
							assign node734 = (inp[1]) ? node812 : node735;
								assign node735 = (inp[14]) ? node773 : node736;
									assign node736 = (inp[3]) ? node750 : node737;
										assign node737 = (inp[7]) ? node747 : node738;
											assign node738 = (inp[9]) ? node740 : 4'b1000;
												assign node740 = (inp[4]) ? node744 : node741;
													assign node741 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node744 = (inp[11]) ? 4'b0000 : 4'b0000;
											assign node747 = (inp[9]) ? 4'b0101 : 4'b1101;
										assign node750 = (inp[7]) ? node760 : node751;
											assign node751 = (inp[9]) ? node757 : node752;
												assign node752 = (inp[4]) ? node754 : 4'b0100;
													assign node754 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node757 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node760 = (inp[4]) ? node766 : node761;
												assign node761 = (inp[12]) ? 4'b1000 : node762;
													assign node762 = (inp[9]) ? 4'b0000 : 4'b0000;
												assign node766 = (inp[10]) ? node770 : node767;
													assign node767 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node770 = (inp[9]) ? 4'b0100 : 4'b0100;
									assign node773 = (inp[11]) ? node797 : node774;
										assign node774 = (inp[10]) ? node790 : node775;
											assign node775 = (inp[12]) ? node783 : node776;
												assign node776 = (inp[13]) ? node780 : node777;
													assign node777 = (inp[7]) ? 4'b1001 : 4'b1001;
													assign node780 = (inp[9]) ? 4'b1001 : 4'b0001;
												assign node783 = (inp[13]) ? node787 : node784;
													assign node784 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node787 = (inp[9]) ? 4'b1101 : 4'b0101;
											assign node790 = (inp[3]) ? 4'b1001 : node791;
												assign node791 = (inp[13]) ? 4'b0001 : node792;
													assign node792 = (inp[4]) ? 4'b1001 : 4'b0001;
										assign node797 = (inp[3]) ? node805 : node798;
											assign node798 = (inp[10]) ? node800 : 4'b0101;
												assign node800 = (inp[7]) ? 4'b1000 : node801;
													assign node801 = (inp[13]) ? 4'b0000 : 4'b0000;
											assign node805 = (inp[13]) ? node807 : 4'b0100;
												assign node807 = (inp[7]) ? 4'b1000 : node808;
													assign node808 = (inp[9]) ? 4'b0100 : 4'b1100;
								assign node812 = (inp[11]) ? node852 : node813;
									assign node813 = (inp[14]) ? node829 : node814;
										assign node814 = (inp[10]) ? node820 : node815;
											assign node815 = (inp[7]) ? node817 : 4'b0101;
												assign node817 = (inp[3]) ? 4'b0101 : 4'b1101;
											assign node820 = (inp[13]) ? node824 : node821;
												assign node821 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node824 = (inp[9]) ? node826 : 4'b1101;
													assign node826 = (inp[12]) ? 4'b0001 : 4'b0001;
										assign node829 = (inp[4]) ? node843 : node830;
											assign node830 = (inp[10]) ? node836 : node831;
												assign node831 = (inp[9]) ? node833 : 4'b0000;
													assign node833 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node836 = (inp[7]) ? node840 : node837;
													assign node837 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node840 = (inp[3]) ? 4'b1000 : 4'b0101;
											assign node843 = (inp[3]) ? node847 : node844;
												assign node844 = (inp[9]) ? 4'b0000 : 4'b1000;
												assign node847 = (inp[10]) ? node849 : 4'b1100;
													assign node849 = (inp[13]) ? 4'b0100 : 4'b0100;
									assign node852 = (inp[9]) ? node872 : node853;
										assign node853 = (inp[4]) ? node865 : node854;
											assign node854 = (inp[14]) ? node860 : node855;
												assign node855 = (inp[10]) ? node857 : 4'b0001;
													assign node857 = (inp[7]) ? 4'b1101 : 4'b0001;
												assign node860 = (inp[3]) ? node862 : 4'b1101;
													assign node862 = (inp[13]) ? 4'b1001 : 4'b1001;
											assign node865 = (inp[3]) ? node867 : 4'b0001;
												assign node867 = (inp[12]) ? node869 : 4'b0101;
													assign node869 = (inp[13]) ? 4'b0101 : 4'b1001;
										assign node872 = (inp[7]) ? node878 : node873;
											assign node873 = (inp[13]) ? 4'b0101 : node874;
												assign node874 = (inp[4]) ? 4'b1101 : 4'b0101;
											assign node878 = (inp[13]) ? node880 : 4'b0101;
												assign node880 = (inp[12]) ? node882 : 4'b0001;
													assign node882 = (inp[10]) ? 4'b0101 : 4'b1001;
							assign node885 = (inp[9]) ? 4'b0101 : 4'b1101;
					assign node888 = (inp[3]) ? node1196 : node889;
						assign node889 = (inp[13]) ? node1039 : node890;
							assign node890 = (inp[7]) ? node966 : node891;
								assign node891 = (inp[0]) ? node925 : node892;
									assign node892 = (inp[1]) ? node910 : node893;
										assign node893 = (inp[10]) ? node897 : node894;
											assign node894 = (inp[9]) ? 4'b0101 : 4'b0000;
											assign node897 = (inp[4]) ? node903 : node898;
												assign node898 = (inp[11]) ? node900 : 4'b0001;
													assign node900 = (inp[9]) ? 4'b1001 : 4'b0001;
												assign node903 = (inp[2]) ? node907 : node904;
													assign node904 = (inp[14]) ? 4'b0001 : 4'b0100;
													assign node907 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node910 = (inp[9]) ? node918 : node911;
											assign node911 = (inp[2]) ? 4'b0001 : node912;
												assign node912 = (inp[10]) ? 4'b0001 : node913;
													assign node913 = (inp[14]) ? 4'b0001 : 4'b1001;
											assign node918 = (inp[4]) ? 4'b0000 : node919;
												assign node919 = (inp[10]) ? 4'b1001 : node920;
													assign node920 = (inp[12]) ? 4'b1100 : 4'b0001;
									assign node925 = (inp[9]) ? node949 : node926;
										assign node926 = (inp[1]) ? node940 : node927;
											assign node927 = (inp[12]) ? node933 : node928;
												assign node928 = (inp[11]) ? 4'b0000 : node929;
													assign node929 = (inp[2]) ? 4'b1001 : 4'b0100;
												assign node933 = (inp[10]) ? node937 : node934;
													assign node934 = (inp[14]) ? 4'b1001 : 4'b1100;
													assign node937 = (inp[4]) ? 4'b0101 : 4'b0000;
											assign node940 = (inp[10]) ? node946 : node941;
												assign node941 = (inp[12]) ? 4'b1101 : node942;
													assign node942 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node946 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node949 = (inp[4]) ? node957 : node950;
											assign node950 = (inp[2]) ? 4'b0101 : node951;
												assign node951 = (inp[11]) ? node953 : 4'b0101;
													assign node953 = (inp[1]) ? 4'b0001 : 4'b1100;
											assign node957 = (inp[10]) ? node963 : node958;
												assign node958 = (inp[12]) ? 4'b0001 : node959;
													assign node959 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node963 = (inp[11]) ? 4'b0101 : 4'b0100;
								assign node966 = (inp[4]) ? node1000 : node967;
									assign node967 = (inp[0]) ? node987 : node968;
										assign node968 = (inp[12]) ? node978 : node969;
											assign node969 = (inp[14]) ? node975 : node970;
												assign node970 = (inp[11]) ? node972 : 4'b0001;
													assign node972 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node975 = (inp[2]) ? 4'b0100 : 4'b1100;
											assign node978 = (inp[10]) ? node984 : node979;
												assign node979 = (inp[9]) ? node981 : 4'b0101;
													assign node981 = (inp[14]) ? 4'b1100 : 4'b0100;
												assign node984 = (inp[9]) ? 4'b0101 : 4'b1101;
										assign node987 = (inp[2]) ? node997 : node988;
											assign node988 = (inp[1]) ? node992 : node989;
												assign node989 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node992 = (inp[11]) ? 4'b0101 : node993;
													assign node993 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node997 = (inp[9]) ? 4'b0101 : 4'b1101;
									assign node1000 = (inp[2]) ? node1018 : node1001;
										assign node1001 = (inp[12]) ? node1007 : node1002;
											assign node1002 = (inp[11]) ? node1004 : 4'b0000;
												assign node1004 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node1007 = (inp[1]) ? node1013 : node1008;
												assign node1008 = (inp[11]) ? node1010 : 4'b0000;
													assign node1010 = (inp[0]) ? 4'b1001 : 4'b0000;
												assign node1013 = (inp[10]) ? node1015 : 4'b1001;
													assign node1015 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node1018 = (inp[12]) ? node1030 : node1019;
											assign node1019 = (inp[1]) ? node1025 : node1020;
												assign node1020 = (inp[0]) ? 4'b0000 : node1021;
													assign node1021 = (inp[9]) ? 4'b1001 : 4'b0101;
												assign node1025 = (inp[10]) ? node1027 : 4'b0101;
													assign node1027 = (inp[0]) ? 4'b0101 : 4'b0001;
											assign node1030 = (inp[0]) ? node1036 : node1031;
												assign node1031 = (inp[10]) ? node1033 : 4'b0101;
													assign node1033 = (inp[9]) ? 4'b0001 : 4'b1001;
												assign node1036 = (inp[9]) ? 4'b0101 : 4'b1101;
							assign node1039 = (inp[4]) ? node1117 : node1040;
								assign node1040 = (inp[11]) ? node1080 : node1041;
									assign node1041 = (inp[0]) ? node1061 : node1042;
										assign node1042 = (inp[7]) ? node1054 : node1043;
											assign node1043 = (inp[9]) ? node1049 : node1044;
												assign node1044 = (inp[14]) ? 4'b1001 : node1045;
													assign node1045 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node1049 = (inp[1]) ? node1051 : 4'b1001;
													assign node1051 = (inp[10]) ? 4'b1001 : 4'b0000;
											assign node1054 = (inp[12]) ? node1056 : 4'b0001;
												assign node1056 = (inp[1]) ? 4'b1000 : node1057;
													assign node1057 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node1061 = (inp[14]) ? node1071 : node1062;
											assign node1062 = (inp[7]) ? node1068 : node1063;
												assign node1063 = (inp[2]) ? node1065 : 4'b0000;
													assign node1065 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node1068 = (inp[12]) ? 4'b1101 : 4'b1000;
											assign node1071 = (inp[2]) ? node1077 : node1072;
												assign node1072 = (inp[1]) ? 4'b0000 : node1073;
													assign node1073 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node1077 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node1080 = (inp[10]) ? node1102 : node1081;
										assign node1081 = (inp[12]) ? node1091 : node1082;
											assign node1082 = (inp[0]) ? node1086 : node1083;
												assign node1083 = (inp[14]) ? 4'b0101 : 4'b1001;
												assign node1086 = (inp[9]) ? node1088 : 4'b0001;
													assign node1088 = (inp[14]) ? 4'b0001 : 4'b0101;
											assign node1091 = (inp[1]) ? node1095 : node1092;
												assign node1092 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node1095 = (inp[0]) ? node1099 : node1096;
													assign node1096 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node1099 = (inp[9]) ? 4'b1001 : 4'b0001;
										assign node1102 = (inp[1]) ? node1110 : node1103;
											assign node1103 = (inp[9]) ? node1105 : 4'b1101;
												assign node1105 = (inp[2]) ? 4'b1000 : node1106;
													assign node1106 = (inp[14]) ? 4'b1001 : 4'b0001;
											assign node1110 = (inp[9]) ? node1112 : 4'b1001;
												assign node1112 = (inp[14]) ? 4'b0101 : node1113;
													assign node1113 = (inp[0]) ? 4'b0001 : 4'b0101;
								assign node1117 = (inp[1]) ? node1161 : node1118;
									assign node1118 = (inp[11]) ? node1140 : node1119;
										assign node1119 = (inp[14]) ? node1131 : node1120;
											assign node1120 = (inp[12]) ? node1126 : node1121;
												assign node1121 = (inp[7]) ? 4'b0000 : node1122;
													assign node1122 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node1126 = (inp[10]) ? node1128 : 4'b1000;
													assign node1128 = (inp[9]) ? 4'b0000 : 4'b1000;
											assign node1131 = (inp[2]) ? node1137 : node1132;
												assign node1132 = (inp[10]) ? node1134 : 4'b0100;
													assign node1134 = (inp[12]) ? 4'b0000 : 4'b0000;
												assign node1137 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node1140 = (inp[2]) ? node1152 : node1141;
											assign node1141 = (inp[7]) ? node1149 : node1142;
												assign node1142 = (inp[10]) ? node1146 : node1143;
													assign node1143 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node1146 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node1149 = (inp[9]) ? 4'b0001 : 4'b1001;
											assign node1152 = (inp[7]) ? node1156 : node1153;
												assign node1153 = (inp[9]) ? 4'b1000 : 4'b0000;
												assign node1156 = (inp[12]) ? 4'b0000 : node1157;
													assign node1157 = (inp[14]) ? 4'b0000 : 4'b0000;
									assign node1161 = (inp[11]) ? node1185 : node1162;
										assign node1162 = (inp[2]) ? node1176 : node1163;
											assign node1163 = (inp[14]) ? node1169 : node1164;
												assign node1164 = (inp[0]) ? node1166 : 4'b0000;
													assign node1166 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node1169 = (inp[10]) ? node1173 : node1170;
													assign node1170 = (inp[9]) ? 4'b0001 : 4'b0100;
													assign node1173 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node1176 = (inp[14]) ? node1182 : node1177;
												assign node1177 = (inp[12]) ? node1179 : 4'b0001;
													assign node1179 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node1182 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node1185 = (inp[9]) ? node1191 : node1186;
											assign node1186 = (inp[10]) ? 4'b1001 : node1187;
												assign node1187 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node1191 = (inp[7]) ? node1193 : 4'b0001;
												assign node1193 = (inp[14]) ? 4'b0001 : 4'b0101;
						assign node1196 = (inp[11]) ? node1318 : node1197;
							assign node1197 = (inp[13]) ? node1263 : node1198;
								assign node1198 = (inp[12]) ? node1238 : node1199;
									assign node1199 = (inp[4]) ? node1219 : node1200;
										assign node1200 = (inp[2]) ? node1212 : node1201;
											assign node1201 = (inp[1]) ? node1209 : node1202;
												assign node1202 = (inp[9]) ? node1206 : node1203;
													assign node1203 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node1206 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node1209 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node1212 = (inp[7]) ? node1216 : node1213;
												assign node1213 = (inp[9]) ? 4'b0000 : 4'b1000;
												assign node1216 = (inp[9]) ? 4'b1000 : 4'b0000;
										assign node1219 = (inp[10]) ? node1231 : node1220;
											assign node1220 = (inp[14]) ? node1226 : node1221;
												assign node1221 = (inp[2]) ? node1223 : 4'b1000;
													assign node1223 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node1226 = (inp[2]) ? 4'b1000 : node1227;
													assign node1227 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node1231 = (inp[2]) ? node1233 : 4'b0000;
												assign node1233 = (inp[14]) ? node1235 : 4'b0001;
													assign node1235 = (inp[1]) ? 4'b0001 : 4'b1000;
									assign node1238 = (inp[4]) ? node1248 : node1239;
										assign node1239 = (inp[1]) ? 4'b0000 : node1240;
											assign node1240 = (inp[14]) ? node1242 : 4'b0000;
												assign node1242 = (inp[10]) ? 4'b1000 : node1243;
													assign node1243 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node1248 = (inp[14]) ? node1256 : node1249;
											assign node1249 = (inp[1]) ? node1251 : 4'b1001;
												assign node1251 = (inp[9]) ? node1253 : 4'b0001;
													assign node1253 = (inp[7]) ? 4'b1000 : 4'b0001;
											assign node1256 = (inp[2]) ? node1258 : 4'b0001;
												assign node1258 = (inp[0]) ? node1260 : 4'b0000;
													assign node1260 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node1263 = (inp[4]) ? node1303 : node1264;
									assign node1264 = (inp[0]) ? node1282 : node1265;
										assign node1265 = (inp[12]) ? node1273 : node1266;
											assign node1266 = (inp[2]) ? 4'b0001 : node1267;
												assign node1267 = (inp[1]) ? 4'b1000 : node1268;
													assign node1268 = (inp[14]) ? 4'b1001 : 4'b0001;
											assign node1273 = (inp[2]) ? node1277 : node1274;
												assign node1274 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node1277 = (inp[7]) ? node1279 : 4'b0000;
													assign node1279 = (inp[9]) ? 4'b1001 : 4'b0000;
										assign node1282 = (inp[9]) ? node1292 : node1283;
											assign node1283 = (inp[12]) ? node1287 : node1284;
												assign node1284 = (inp[10]) ? 4'b1000 : 4'b0001;
												assign node1287 = (inp[10]) ? 4'b0001 : node1288;
													assign node1288 = (inp[2]) ? 4'b1000 : 4'b0001;
											assign node1292 = (inp[10]) ? node1298 : node1293;
												assign node1293 = (inp[12]) ? node1295 : 4'b1000;
													assign node1295 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node1298 = (inp[12]) ? node1300 : 4'b0000;
													assign node1300 = (inp[1]) ? 4'b0000 : 4'b1000;
									assign node1303 = (inp[10]) ? node1313 : node1304;
										assign node1304 = (inp[7]) ? 4'b0000 : node1305;
											assign node1305 = (inp[9]) ? node1309 : node1306;
												assign node1306 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1309 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node1313 = (inp[1]) ? 4'b0000 : node1314;
											assign node1314 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node1318 = (inp[1]) ? node1388 : node1319;
								assign node1319 = (inp[4]) ? node1359 : node1320;
									assign node1320 = (inp[12]) ? node1342 : node1321;
										assign node1321 = (inp[9]) ? node1331 : node1322;
											assign node1322 = (inp[13]) ? node1328 : node1323;
												assign node1323 = (inp[2]) ? node1325 : 4'b0000;
													assign node1325 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node1328 = (inp[0]) ? 4'b0001 : 4'b1000;
											assign node1331 = (inp[0]) ? node1337 : node1332;
												assign node1332 = (inp[2]) ? 4'b0001 : node1333;
													assign node1333 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node1337 = (inp[14]) ? 4'b1000 : node1338;
													assign node1338 = (inp[13]) ? 4'b0000 : 4'b1001;
										assign node1342 = (inp[14]) ? node1350 : node1343;
											assign node1343 = (inp[0]) ? node1347 : node1344;
												assign node1344 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node1347 = (inp[13]) ? 4'b0001 : 4'b1000;
											assign node1350 = (inp[2]) ? node1356 : node1351;
												assign node1351 = (inp[0]) ? 4'b1001 : node1352;
													assign node1352 = (inp[9]) ? 4'b0001 : 4'b1001;
												assign node1356 = (inp[9]) ? 4'b1000 : 4'b1001;
									assign node1359 = (inp[10]) ? node1377 : node1360;
										assign node1360 = (inp[2]) ? node1366 : node1361;
											assign node1361 = (inp[13]) ? 4'b0001 : node1362;
												assign node1362 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node1366 = (inp[12]) ? node1372 : node1367;
												assign node1367 = (inp[13]) ? 4'b0001 : node1368;
													assign node1368 = (inp[9]) ? 4'b1000 : 4'b0001;
												assign node1372 = (inp[0]) ? 4'b0000 : node1373;
													assign node1373 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node1377 = (inp[13]) ? 4'b0000 : node1378;
											assign node1378 = (inp[2]) ? node1382 : node1379;
												assign node1379 = (inp[0]) ? 4'b0001 : 4'b1000;
												assign node1382 = (inp[7]) ? node1384 : 4'b0000;
													assign node1384 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node1388 = (inp[4]) ? node1418 : node1389;
									assign node1389 = (inp[10]) ? node1401 : node1390;
										assign node1390 = (inp[9]) ? node1396 : node1391;
											assign node1391 = (inp[7]) ? node1393 : 4'b0001;
												assign node1393 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node1396 = (inp[7]) ? node1398 : 4'b1001;
												assign node1398 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node1401 = (inp[14]) ? node1413 : node1402;
											assign node1402 = (inp[2]) ? node1408 : node1403;
												assign node1403 = (inp[7]) ? node1405 : 4'b0001;
													assign node1405 = (inp[12]) ? 4'b0001 : 4'b0001;
												assign node1408 = (inp[7]) ? node1410 : 4'b1001;
													assign node1410 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node1413 = (inp[13]) ? node1415 : 4'b0001;
												assign node1415 = (inp[9]) ? 4'b0001 : 4'b1001;
									assign node1418 = (inp[13]) ? node1424 : node1419;
										assign node1419 = (inp[10]) ? 4'b0001 : node1420;
											assign node1420 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node1424 = (inp[10]) ? 4'b0000 : 4'b0001;
			assign node1427 = (inp[9]) ? node1987 : node1428;
				assign node1428 = (inp[6]) ? node1568 : node1429;
					assign node1429 = (inp[0]) ? 4'b1001 : node1430;
						assign node1430 = (inp[5]) ? node1462 : node1431;
							assign node1431 = (inp[3]) ? node1433 : 4'b1011;
								assign node1433 = (inp[2]) ? 4'b1011 : node1434;
									assign node1434 = (inp[4]) ? node1442 : node1435;
										assign node1435 = (inp[7]) ? 4'b1011 : node1436;
											assign node1436 = (inp[13]) ? node1438 : 4'b0001;
												assign node1438 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node1442 = (inp[13]) ? node1456 : node1443;
											assign node1443 = (inp[10]) ? node1451 : node1444;
												assign node1444 = (inp[7]) ? node1448 : node1445;
													assign node1445 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node1448 = (inp[1]) ? 4'b0001 : 4'b1011;
												assign node1451 = (inp[11]) ? 4'b0000 : node1452;
													assign node1452 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node1456 = (inp[10]) ? 4'b1001 : node1457;
												assign node1457 = (inp[12]) ? 4'b0000 : 4'b1000;
							assign node1462 = (inp[2]) ? node1538 : node1463;
								assign node1463 = (inp[13]) ? node1509 : node1464;
									assign node1464 = (inp[3]) ? node1490 : node1465;
										assign node1465 = (inp[7]) ? node1477 : node1466;
											assign node1466 = (inp[12]) ? node1472 : node1467;
												assign node1467 = (inp[14]) ? node1469 : 4'b0101;
													assign node1469 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node1472 = (inp[10]) ? node1474 : 4'b1100;
													assign node1474 = (inp[1]) ? 4'b0100 : 4'b0100;
											assign node1477 = (inp[4]) ? node1485 : node1478;
												assign node1478 = (inp[12]) ? node1482 : node1479;
													assign node1479 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1482 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node1485 = (inp[12]) ? node1487 : 4'b0101;
													assign node1487 = (inp[10]) ? 4'b0101 : 4'b1001;
										assign node1490 = (inp[1]) ? node1496 : node1491;
											assign node1491 = (inp[4]) ? 4'b0000 : node1492;
												assign node1492 = (inp[11]) ? 4'b0000 : 4'b0101;
											assign node1496 = (inp[10]) ? node1504 : node1497;
												assign node1497 = (inp[12]) ? node1501 : node1498;
													assign node1498 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node1501 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node1504 = (inp[14]) ? node1506 : 4'b0001;
													assign node1506 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node1509 = (inp[1]) ? node1523 : node1510;
										assign node1510 = (inp[3]) ? node1516 : node1511;
											assign node1511 = (inp[7]) ? node1513 : 4'b1100;
												assign node1513 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node1516 = (inp[14]) ? 4'b0101 : node1517;
												assign node1517 = (inp[12]) ? node1519 : 4'b1000;
													assign node1519 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node1523 = (inp[14]) ? node1529 : node1524;
											assign node1524 = (inp[12]) ? node1526 : 4'b1001;
												assign node1526 = (inp[10]) ? 4'b1001 : 4'b0101;
											assign node1529 = (inp[3]) ? node1535 : node1530;
												assign node1530 = (inp[11]) ? node1532 : 4'b0100;
													assign node1532 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node1535 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node1538 = (inp[3]) ? node1540 : 4'b1011;
									assign node1540 = (inp[14]) ? node1552 : node1541;
										assign node1541 = (inp[7]) ? node1547 : node1542;
											assign node1542 = (inp[1]) ? 4'b1001 : node1543;
												assign node1543 = (inp[4]) ? 4'b1000 : 4'b0000;
											assign node1547 = (inp[1]) ? node1549 : 4'b1011;
												assign node1549 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node1552 = (inp[7]) ? node1558 : node1553;
											assign node1553 = (inp[13]) ? node1555 : 4'b0000;
												assign node1555 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1558 = (inp[13]) ? node1562 : node1559;
												assign node1559 = (inp[12]) ? 4'b1011 : 4'b0000;
												assign node1562 = (inp[12]) ? node1564 : 4'b1000;
													assign node1564 = (inp[10]) ? 4'b1000 : 4'b0000;
					assign node1568 = (inp[0]) ? node1844 : node1569;
						assign node1569 = (inp[1]) ? node1713 : node1570;
							assign node1570 = (inp[3]) ? node1642 : node1571;
								assign node1571 = (inp[4]) ? node1611 : node1572;
									assign node1572 = (inp[7]) ? node1586 : node1573;
										assign node1573 = (inp[2]) ? node1575 : 4'b0100;
											assign node1575 = (inp[14]) ? node1581 : node1576;
												assign node1576 = (inp[10]) ? node1578 : 4'b1000;
													assign node1578 = (inp[13]) ? 4'b1000 : 4'b0100;
												assign node1581 = (inp[10]) ? node1583 : 4'b0101;
													assign node1583 = (inp[11]) ? 4'b0100 : 4'b0100;
										assign node1586 = (inp[14]) ? node1596 : node1587;
											assign node1587 = (inp[5]) ? node1593 : node1588;
												assign node1588 = (inp[2]) ? node1590 : 4'b0000;
													assign node1590 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node1593 = (inp[12]) ? 4'b0000 : 4'b1001;
											assign node1596 = (inp[5]) ? node1604 : node1597;
												assign node1597 = (inp[11]) ? node1601 : node1598;
													assign node1598 = (inp[2]) ? 4'b0001 : 4'b0001;
													assign node1601 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node1604 = (inp[13]) ? node1608 : node1605;
													assign node1605 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node1608 = (inp[10]) ? 4'b0100 : 4'b1100;
									assign node1611 = (inp[11]) ? node1627 : node1612;
										assign node1612 = (inp[10]) ? node1620 : node1613;
											assign node1613 = (inp[12]) ? 4'b0100 : node1614;
												assign node1614 = (inp[14]) ? 4'b0000 : node1615;
													assign node1615 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node1620 = (inp[7]) ? node1622 : 4'b1000;
												assign node1622 = (inp[13]) ? node1624 : 4'b1001;
													assign node1624 = (inp[2]) ? 4'b0100 : 4'b1001;
										assign node1627 = (inp[7]) ? node1633 : node1628;
											assign node1628 = (inp[14]) ? 4'b0001 : node1629;
												assign node1629 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node1633 = (inp[10]) ? node1635 : 4'b0000;
												assign node1635 = (inp[13]) ? node1639 : node1636;
													assign node1636 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node1639 = (inp[5]) ? 4'b0100 : 4'b0001;
								assign node1642 = (inp[5]) ? node1676 : node1643;
									assign node1643 = (inp[12]) ? node1661 : node1644;
										assign node1644 = (inp[4]) ? node1654 : node1645;
											assign node1645 = (inp[13]) ? node1651 : node1646;
												assign node1646 = (inp[11]) ? node1648 : 4'b0101;
													assign node1648 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1651 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node1654 = (inp[14]) ? node1656 : 4'b0001;
												assign node1656 = (inp[11]) ? node1658 : 4'b1000;
													assign node1658 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node1661 = (inp[10]) ? node1665 : node1662;
											assign node1662 = (inp[13]) ? 4'b0100 : 4'b1100;
											assign node1665 = (inp[4]) ? node1673 : node1666;
												assign node1666 = (inp[7]) ? node1670 : node1667;
													assign node1667 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node1670 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node1673 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node1676 = (inp[13]) ? node1694 : node1677;
										assign node1677 = (inp[11]) ? node1689 : node1678;
											assign node1678 = (inp[7]) ? node1684 : node1679;
												assign node1679 = (inp[10]) ? 4'b1000 : node1680;
													assign node1680 = (inp[4]) ? 4'b0000 : 4'b0000;
												assign node1684 = (inp[12]) ? node1686 : 4'b0001;
													assign node1686 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node1689 = (inp[2]) ? 4'b1000 : node1690;
												assign node1690 = (inp[12]) ? 4'b0000 : 4'b1001;
										assign node1694 = (inp[4]) ? node1706 : node1695;
											assign node1695 = (inp[11]) ? node1701 : node1696;
												assign node1696 = (inp[7]) ? node1698 : 4'b1000;
													assign node1698 = (inp[12]) ? 4'b0000 : 4'b0000;
												assign node1701 = (inp[14]) ? 4'b1001 : node1702;
													assign node1702 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node1706 = (inp[10]) ? 4'b0000 : node1707;
												assign node1707 = (inp[12]) ? 4'b0001 : node1708;
													assign node1708 = (inp[7]) ? 4'b0001 : 4'b0000;
							assign node1713 = (inp[11]) ? node1779 : node1714;
								assign node1714 = (inp[5]) ? node1752 : node1715;
									assign node1715 = (inp[14]) ? node1733 : node1716;
										assign node1716 = (inp[2]) ? node1724 : node1717;
											assign node1717 = (inp[7]) ? node1721 : node1718;
												assign node1718 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node1721 = (inp[3]) ? 4'b1000 : 4'b1001;
											assign node1724 = (inp[13]) ? node1728 : node1725;
												assign node1725 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node1728 = (inp[3]) ? node1730 : 4'b1101;
													assign node1730 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node1733 = (inp[13]) ? node1741 : node1734;
											assign node1734 = (inp[12]) ? node1736 : 4'b0100;
												assign node1736 = (inp[2]) ? node1738 : 4'b1000;
													assign node1738 = (inp[10]) ? 4'b0100 : 4'b1100;
											assign node1741 = (inp[10]) ? node1749 : node1742;
												assign node1742 = (inp[3]) ? node1746 : node1743;
													assign node1743 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node1746 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node1749 = (inp[12]) ? 4'b1100 : 4'b1000;
									assign node1752 = (inp[4]) ? node1762 : node1753;
										assign node1753 = (inp[10]) ? node1757 : node1754;
											assign node1754 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node1757 = (inp[3]) ? 4'b0001 : node1758;
												assign node1758 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node1762 = (inp[10]) ? node1772 : node1763;
											assign node1763 = (inp[3]) ? node1769 : node1764;
												assign node1764 = (inp[12]) ? 4'b0001 : node1765;
													assign node1765 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node1769 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node1772 = (inp[7]) ? 4'b0000 : node1773;
												assign node1773 = (inp[13]) ? 4'b0000 : node1774;
													assign node1774 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node1779 = (inp[3]) ? node1813 : node1780;
									assign node1780 = (inp[7]) ? node1800 : node1781;
										assign node1781 = (inp[10]) ? node1793 : node1782;
											assign node1782 = (inp[5]) ? node1788 : node1783;
												assign node1783 = (inp[13]) ? node1785 : 4'b1001;
													assign node1785 = (inp[14]) ? 4'b0101 : 4'b0001;
												assign node1788 = (inp[13]) ? 4'b1001 : node1789;
													assign node1789 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node1793 = (inp[2]) ? node1795 : 4'b0101;
												assign node1795 = (inp[13]) ? 4'b1101 : node1796;
													assign node1796 = (inp[5]) ? 4'b1101 : 4'b0101;
										assign node1800 = (inp[10]) ? node1810 : node1801;
											assign node1801 = (inp[12]) ? node1807 : node1802;
												assign node1802 = (inp[13]) ? node1804 : 4'b0101;
													assign node1804 = (inp[14]) ? 4'b1001 : 4'b0101;
												assign node1807 = (inp[5]) ? 4'b0001 : 4'b1001;
											assign node1810 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node1813 = (inp[4]) ? node1827 : node1814;
										assign node1814 = (inp[7]) ? node1822 : node1815;
											assign node1815 = (inp[2]) ? 4'b0001 : node1816;
												assign node1816 = (inp[5]) ? node1818 : 4'b0101;
													assign node1818 = (inp[12]) ? 4'b0001 : 4'b0001;
											assign node1822 = (inp[5]) ? node1824 : 4'b1101;
												assign node1824 = (inp[2]) ? 4'b0001 : 4'b1001;
										assign node1827 = (inp[12]) ? node1837 : node1828;
											assign node1828 = (inp[10]) ? node1834 : node1829;
												assign node1829 = (inp[2]) ? node1831 : 4'b0001;
													assign node1831 = (inp[5]) ? 4'b1001 : 4'b0001;
												assign node1834 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node1837 = (inp[10]) ? node1841 : node1838;
												assign node1838 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node1841 = (inp[13]) ? 4'b1001 : 4'b0001;
						assign node1844 = (inp[2]) ? node1956 : node1845;
							assign node1845 = (inp[5]) ? node1881 : node1846;
								assign node1846 = (inp[3]) ? node1848 : 4'b1001;
									assign node1848 = (inp[1]) ? node1866 : node1849;
										assign node1849 = (inp[7]) ? node1861 : node1850;
											assign node1850 = (inp[10]) ? node1858 : node1851;
												assign node1851 = (inp[13]) ? node1855 : node1852;
													assign node1852 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node1855 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node1858 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node1861 = (inp[4]) ? node1863 : 4'b1001;
												assign node1863 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node1866 = (inp[13]) ? node1876 : node1867;
											assign node1867 = (inp[7]) ? node1871 : node1868;
												assign node1868 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node1871 = (inp[4]) ? node1873 : 4'b1001;
													assign node1873 = (inp[10]) ? 4'b0001 : 4'b0001;
											assign node1876 = (inp[7]) ? node1878 : 4'b1001;
												assign node1878 = (inp[10]) ? 4'b1001 : 4'b1000;
								assign node1881 = (inp[3]) ? node1923 : node1882;
									assign node1882 = (inp[4]) ? node1902 : node1883;
										assign node1883 = (inp[7]) ? node1897 : node1884;
											assign node1884 = (inp[1]) ? node1890 : node1885;
												assign node1885 = (inp[13]) ? 4'b0101 : node1886;
													assign node1886 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node1890 = (inp[13]) ? node1894 : node1891;
													assign node1891 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node1894 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node1897 = (inp[12]) ? 4'b0000 : node1898;
												assign node1898 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node1902 = (inp[7]) ? node1912 : node1903;
											assign node1903 = (inp[11]) ? node1909 : node1904;
												assign node1904 = (inp[10]) ? node1906 : 4'b0000;
													assign node1906 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node1909 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node1912 = (inp[12]) ? node1916 : node1913;
												assign node1913 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node1916 = (inp[11]) ? node1920 : node1917;
													assign node1917 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node1920 = (inp[1]) ? 4'b0001 : 4'b0100;
									assign node1923 = (inp[4]) ? node1941 : node1924;
										assign node1924 = (inp[13]) ? node1934 : node1925;
											assign node1925 = (inp[11]) ? node1929 : node1926;
												assign node1926 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node1929 = (inp[7]) ? 4'b1001 : node1930;
													assign node1930 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node1934 = (inp[10]) ? 4'b1001 : node1935;
												assign node1935 = (inp[12]) ? 4'b1001 : node1936;
													assign node1936 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node1941 = (inp[13]) ? node1949 : node1942;
											assign node1942 = (inp[12]) ? 4'b1000 : node1943;
												assign node1943 = (inp[7]) ? 4'b0001 : node1944;
													assign node1944 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node1949 = (inp[10]) ? 4'b0000 : node1950;
												assign node1950 = (inp[14]) ? node1952 : 4'b0001;
													assign node1952 = (inp[12]) ? 4'b0000 : 4'b0000;
							assign node1956 = (inp[5]) ? node1958 : 4'b1001;
								assign node1958 = (inp[3]) ? node1960 : 4'b1001;
									assign node1960 = (inp[4]) ? node1972 : node1961;
										assign node1961 = (inp[7]) ? 4'b1001 : node1962;
											assign node1962 = (inp[12]) ? node1968 : node1963;
												assign node1963 = (inp[11]) ? 4'b0000 : node1964;
													assign node1964 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node1968 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node1972 = (inp[13]) ? node1982 : node1973;
											assign node1973 = (inp[7]) ? node1977 : node1974;
												assign node1974 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node1977 = (inp[12]) ? 4'b0000 : node1978;
													assign node1978 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1982 = (inp[10]) ? 4'b0000 : node1983;
												assign node1983 = (inp[14]) ? 4'b0000 : 4'b0001;
				assign node1987 = (inp[0]) ? node2395 : node1988;
					assign node1988 = (inp[6]) ? node2102 : node1989;
						assign node1989 = (inp[2]) ? node2073 : node1990;
							assign node1990 = (inp[5]) ? node2018 : node1991;
								assign node1991 = (inp[3]) ? node1993 : 4'b0011;
									assign node1993 = (inp[7]) ? node2009 : node1994;
										assign node1994 = (inp[4]) ? node2000 : node1995;
											assign node1995 = (inp[13]) ? node1997 : 4'b0011;
												assign node1997 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node2000 = (inp[10]) ? node2006 : node2001;
												assign node2001 = (inp[12]) ? 4'b0000 : node2002;
													assign node2002 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node2006 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node2009 = (inp[13]) ? node2011 : 4'b0011;
											assign node2011 = (inp[11]) ? node2015 : node2012;
												assign node2012 = (inp[1]) ? 4'b0001 : 4'b0011;
												assign node2015 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node2018 = (inp[11]) ? node2042 : node2019;
									assign node2019 = (inp[14]) ? node2025 : node2020;
										assign node2020 = (inp[1]) ? node2022 : 4'b1000;
											assign node2022 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node2025 = (inp[1]) ? node2033 : node2026;
											assign node2026 = (inp[13]) ? 4'b1001 : node2027;
												assign node2027 = (inp[10]) ? 4'b0101 : node2028;
													assign node2028 = (inp[12]) ? 4'b0001 : 4'b0001;
											assign node2033 = (inp[13]) ? node2039 : node2034;
												assign node2034 = (inp[12]) ? 4'b1100 : node2035;
													assign node2035 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node2039 = (inp[3]) ? 4'b0000 : 4'b1000;
									assign node2042 = (inp[1]) ? node2064 : node2043;
										assign node2043 = (inp[14]) ? node2053 : node2044;
											assign node2044 = (inp[7]) ? 4'b1100 : node2045;
												assign node2045 = (inp[12]) ? node2049 : node2046;
													assign node2046 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node2049 = (inp[13]) ? 4'b1000 : 4'b1000;
											assign node2053 = (inp[13]) ? node2059 : node2054;
												assign node2054 = (inp[10]) ? 4'b1100 : node2055;
													assign node2055 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node2059 = (inp[3]) ? 4'b0000 : node2060;
													assign node2060 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node2064 = (inp[3]) ? 4'b0001 : node2065;
											assign node2065 = (inp[4]) ? 4'b0101 : node2066;
												assign node2066 = (inp[7]) ? 4'b0001 : node2067;
													assign node2067 = (inp[10]) ? 4'b0101 : 4'b1001;
							assign node2073 = (inp[3]) ? node2075 : 4'b0011;
								assign node2075 = (inp[5]) ? node2077 : 4'b0011;
									assign node2077 = (inp[7]) ? node2093 : node2078;
										assign node2078 = (inp[4]) ? node2088 : node2079;
											assign node2079 = (inp[10]) ? node2083 : node2080;
												assign node2080 = (inp[1]) ? 4'b0001 : 4'b0011;
												assign node2083 = (inp[1]) ? 4'b0001 : node2084;
													assign node2084 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node2088 = (inp[14]) ? 4'b1000 : node2089;
												assign node2089 = (inp[1]) ? 4'b0001 : 4'b1000;
										assign node2093 = (inp[13]) ? node2095 : 4'b0011;
											assign node2095 = (inp[14]) ? 4'b0011 : node2096;
												assign node2096 = (inp[12]) ? 4'b0011 : node2097;
													assign node2097 = (inp[10]) ? 4'b0000 : 4'b0001;
						assign node2102 = (inp[5]) ? node2242 : node2103;
							assign node2103 = (inp[11]) ? node2181 : node2104;
								assign node2104 = (inp[13]) ? node2142 : node2105;
									assign node2105 = (inp[12]) ? node2123 : node2106;
										assign node2106 = (inp[3]) ? node2118 : node2107;
											assign node2107 = (inp[7]) ? node2113 : node2108;
												assign node2108 = (inp[1]) ? 4'b1101 : node2109;
													assign node2109 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node2113 = (inp[10]) ? node2115 : 4'b0001;
													assign node2115 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node2118 = (inp[4]) ? 4'b1100 : node2119;
												assign node2119 = (inp[14]) ? 4'b1101 : 4'b1000;
										assign node2123 = (inp[2]) ? node2127 : node2124;
											assign node2124 = (inp[3]) ? 4'b1000 : 4'b0001;
											assign node2127 = (inp[10]) ? node2135 : node2128;
												assign node2128 = (inp[14]) ? node2132 : node2129;
													assign node2129 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node2132 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node2135 = (inp[1]) ? node2139 : node2136;
													assign node2136 = (inp[14]) ? 4'b0001 : 4'b1100;
													assign node2139 = (inp[14]) ? 4'b1100 : 4'b1101;
									assign node2142 = (inp[4]) ? node2162 : node2143;
										assign node2143 = (inp[12]) ? node2155 : node2144;
											assign node2144 = (inp[10]) ? node2152 : node2145;
												assign node2145 = (inp[1]) ? node2149 : node2146;
													assign node2146 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node2149 = (inp[2]) ? 4'b0101 : 4'b0000;
												assign node2152 = (inp[3]) ? 4'b0100 : 4'b0101;
											assign node2155 = (inp[14]) ? node2157 : 4'b0000;
												assign node2157 = (inp[10]) ? node2159 : 4'b1100;
													assign node2159 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node2162 = (inp[10]) ? node2174 : node2163;
											assign node2163 = (inp[1]) ? node2169 : node2164;
												assign node2164 = (inp[2]) ? 4'b1001 : node2165;
													assign node2165 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node2169 = (inp[14]) ? node2171 : 4'b1001;
													assign node2171 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node2174 = (inp[1]) ? 4'b0000 : node2175;
												assign node2175 = (inp[14]) ? node2177 : 4'b1001;
													assign node2177 = (inp[12]) ? 4'b1001 : 4'b0000;
								assign node2181 = (inp[1]) ? node2219 : node2182;
									assign node2182 = (inp[3]) ? node2200 : node2183;
										assign node2183 = (inp[13]) ? node2191 : node2184;
											assign node2184 = (inp[12]) ? 4'b0000 : node2185;
												assign node2185 = (inp[10]) ? 4'b1000 : node2186;
													assign node2186 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node2191 = (inp[12]) ? node2197 : node2192;
												assign node2192 = (inp[4]) ? node2194 : 4'b0100;
													assign node2194 = (inp[7]) ? 4'b0100 : 4'b1001;
												assign node2197 = (inp[10]) ? 4'b0100 : 4'b1000;
										assign node2200 = (inp[4]) ? node2210 : node2201;
											assign node2201 = (inp[2]) ? node2203 : 4'b1101;
												assign node2203 = (inp[13]) ? node2207 : node2204;
													assign node2204 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2207 = (inp[14]) ? 4'b0000 : 4'b1100;
											assign node2210 = (inp[2]) ? node2216 : node2211;
												assign node2211 = (inp[10]) ? node2213 : 4'b1101;
													assign node2213 = (inp[12]) ? 4'b1101 : 4'b0000;
												assign node2216 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node2219 = (inp[10]) ? node2231 : node2220;
										assign node2220 = (inp[4]) ? node2224 : node2221;
											assign node2221 = (inp[3]) ? 4'b0001 : 4'b1001;
											assign node2224 = (inp[12]) ? node2228 : node2225;
												assign node2225 = (inp[14]) ? 4'b1001 : 4'b1101;
												assign node2228 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node2231 = (inp[13]) ? 4'b0101 : node2232;
											assign node2232 = (inp[12]) ? node2238 : node2233;
												assign node2233 = (inp[2]) ? node2235 : 4'b0101;
													assign node2235 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node2238 = (inp[3]) ? 4'b0001 : 4'b1001;
							assign node2242 = (inp[1]) ? node2318 : node2243;
								assign node2243 = (inp[2]) ? node2275 : node2244;
									assign node2244 = (inp[11]) ? node2260 : node2245;
										assign node2245 = (inp[14]) ? node2253 : node2246;
											assign node2246 = (inp[7]) ? node2250 : node2247;
												assign node2247 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node2250 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node2253 = (inp[3]) ? node2255 : 4'b0001;
												assign node2255 = (inp[4]) ? 4'b0000 : node2256;
													assign node2256 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node2260 = (inp[4]) ? node2268 : node2261;
											assign node2261 = (inp[3]) ? node2265 : node2262;
												assign node2262 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node2265 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node2268 = (inp[3]) ? 4'b0000 : node2269;
												assign node2269 = (inp[10]) ? node2271 : 4'b0000;
													assign node2271 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node2275 = (inp[3]) ? node2297 : node2276;
										assign node2276 = (inp[12]) ? node2290 : node2277;
											assign node2277 = (inp[10]) ? node2283 : node2278;
												assign node2278 = (inp[14]) ? node2280 : 4'b1000;
													assign node2280 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node2283 = (inp[11]) ? node2287 : node2284;
													assign node2284 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node2287 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node2290 = (inp[7]) ? node2292 : 4'b0001;
												assign node2292 = (inp[13]) ? node2294 : 4'b0000;
													assign node2294 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node2297 = (inp[14]) ? node2303 : node2298;
											assign node2298 = (inp[13]) ? node2300 : 4'b0000;
												assign node2300 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node2303 = (inp[4]) ? node2311 : node2304;
												assign node2304 = (inp[11]) ? node2308 : node2305;
													assign node2305 = (inp[13]) ? 4'b1000 : 4'b0001;
													assign node2308 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node2311 = (inp[13]) ? node2315 : node2312;
													assign node2312 = (inp[12]) ? 4'b0000 : 4'b1001;
													assign node2315 = (inp[7]) ? 4'b0000 : 4'b0000;
								assign node2318 = (inp[11]) ? node2362 : node2319;
									assign node2319 = (inp[3]) ? node2343 : node2320;
										assign node2320 = (inp[4]) ? node2334 : node2321;
											assign node2321 = (inp[10]) ? node2327 : node2322;
												assign node2322 = (inp[2]) ? 4'b1000 : node2323;
													assign node2323 = (inp[7]) ? 4'b1100 : 4'b0100;
												assign node2327 = (inp[14]) ? node2331 : node2328;
													assign node2328 = (inp[2]) ? 4'b0100 : 4'b1100;
													assign node2331 = (inp[2]) ? 4'b0100 : 4'b0001;
											assign node2334 = (inp[7]) ? node2338 : node2335;
												assign node2335 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node2338 = (inp[10]) ? node2340 : 4'b1100;
													assign node2340 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node2343 = (inp[4]) ? node2355 : node2344;
											assign node2344 = (inp[12]) ? node2348 : node2345;
												assign node2345 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node2348 = (inp[13]) ? node2352 : node2349;
													assign node2349 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2352 = (inp[2]) ? 4'b1001 : 4'b0001;
											assign node2355 = (inp[13]) ? 4'b0000 : node2356;
												assign node2356 = (inp[7]) ? node2358 : 4'b0001;
													assign node2358 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node2362 = (inp[3]) ? node2382 : node2363;
										assign node2363 = (inp[2]) ? node2371 : node2364;
											assign node2364 = (inp[13]) ? node2368 : node2365;
												assign node2365 = (inp[4]) ? 4'b0001 : 4'b1001;
												assign node2368 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node2371 = (inp[7]) ? node2377 : node2372;
												assign node2372 = (inp[14]) ? 4'b1001 : node2373;
													assign node2373 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node2377 = (inp[10]) ? 4'b1001 : node2378;
													assign node2378 = (inp[4]) ? 4'b0001 : 4'b1001;
										assign node2382 = (inp[4]) ? node2390 : node2383;
											assign node2383 = (inp[2]) ? node2385 : 4'b0001;
												assign node2385 = (inp[14]) ? 4'b0001 : node2386;
													assign node2386 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2390 = (inp[13]) ? node2392 : 4'b0001;
												assign node2392 = (inp[10]) ? 4'b0000 : 4'b0001;
					assign node2395 = (inp[6]) ? node2397 : 4'b0001;
						assign node2397 = (inp[2]) ? node2499 : node2398;
							assign node2398 = (inp[5]) ? node2422 : node2399;
								assign node2399 = (inp[3]) ? node2401 : 4'b0001;
									assign node2401 = (inp[7]) ? 4'b0001 : node2402;
										assign node2402 = (inp[4]) ? node2410 : node2403;
											assign node2403 = (inp[13]) ? node2405 : 4'b0001;
												assign node2405 = (inp[10]) ? 4'b0000 : node2406;
													assign node2406 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node2410 = (inp[1]) ? node2416 : node2411;
												assign node2411 = (inp[14]) ? 4'b1001 : node2412;
													assign node2412 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node2416 = (inp[10]) ? 4'b1001 : node2417;
													assign node2417 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node2422 = (inp[1]) ? node2462 : node2423;
									assign node2423 = (inp[7]) ? node2443 : node2424;
										assign node2424 = (inp[3]) ? node2436 : node2425;
											assign node2425 = (inp[10]) ? node2431 : node2426;
												assign node2426 = (inp[12]) ? 4'b0100 : node2427;
													assign node2427 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node2431 = (inp[13]) ? 4'b0101 : node2432;
													assign node2432 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node2436 = (inp[10]) ? 4'b0000 : node2437;
												assign node2437 = (inp[11]) ? node2439 : 4'b1001;
													assign node2439 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node2443 = (inp[3]) ? node2455 : node2444;
											assign node2444 = (inp[14]) ? node2450 : node2445;
												assign node2445 = (inp[13]) ? 4'b0000 : node2446;
													assign node2446 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2450 = (inp[11]) ? node2452 : 4'b0001;
													assign node2452 = (inp[10]) ? 4'b0001 : 4'b1000;
											assign node2455 = (inp[11]) ? 4'b0000 : node2456;
												assign node2456 = (inp[10]) ? 4'b0000 : node2457;
													assign node2457 = (inp[14]) ? 4'b0000 : 4'b0000;
									assign node2462 = (inp[11]) ? node2484 : node2463;
										assign node2463 = (inp[4]) ? node2475 : node2464;
											assign node2464 = (inp[10]) ? node2470 : node2465;
												assign node2465 = (inp[7]) ? 4'b1000 : node2466;
													assign node2466 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node2470 = (inp[13]) ? node2472 : 4'b1001;
													assign node2472 = (inp[3]) ? 4'b0001 : 4'b0000;
											assign node2475 = (inp[3]) ? node2479 : node2476;
												assign node2476 = (inp[10]) ? 4'b0000 : 4'b1100;
												assign node2479 = (inp[12]) ? node2481 : 4'b0000;
													assign node2481 = (inp[13]) ? 4'b0000 : 4'b0000;
										assign node2484 = (inp[13]) ? node2490 : node2485;
											assign node2485 = (inp[12]) ? node2487 : 4'b1001;
												assign node2487 = (inp[4]) ? 4'b0001 : 4'b1001;
											assign node2490 = (inp[12]) ? node2496 : node2491;
												assign node2491 = (inp[3]) ? node2493 : 4'b0001;
													assign node2493 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node2496 = (inp[3]) ? 4'b0001 : 4'b1001;
							assign node2499 = (inp[5]) ? node2501 : 4'b0001;
								assign node2501 = (inp[3]) ? node2503 : 4'b0001;
									assign node2503 = (inp[4]) ? node2511 : node2504;
										assign node2504 = (inp[13]) ? node2506 : 4'b0001;
											assign node2506 = (inp[14]) ? 4'b0001 : node2507;
												assign node2507 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node2511 = (inp[13]) ? node2519 : node2512;
											assign node2512 = (inp[12]) ? 4'b0000 : node2513;
												assign node2513 = (inp[10]) ? 4'b0001 : node2514;
													assign node2514 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node2519 = (inp[10]) ? 4'b0000 : node2520;
												assign node2520 = (inp[12]) ? 4'b0001 : node2521;
													assign node2521 = (inp[11]) ? 4'b0000 : 4'b0001;
		assign node2526 = (inp[9]) ? node3786 : node2527;
			assign node2527 = (inp[6]) ? node2865 : node2528;
				assign node2528 = (inp[15]) ? node2728 : node2529;
					assign node2529 = (inp[0]) ? 4'b1100 : node2530;
						assign node2530 = (inp[2]) ? node2666 : node2531;
							assign node2531 = (inp[1]) ? node2603 : node2532;
								assign node2532 = (inp[13]) ? node2568 : node2533;
									assign node2533 = (inp[3]) ? node2547 : node2534;
										assign node2534 = (inp[5]) ? node2538 : node2535;
											assign node2535 = (inp[4]) ? 4'b1001 : 4'b1110;
											assign node2538 = (inp[11]) ? 4'b1101 : node2539;
												assign node2539 = (inp[4]) ? node2543 : node2540;
													assign node2540 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node2543 = (inp[12]) ? 4'b1101 : 4'b0001;
										assign node2547 = (inp[7]) ? node2559 : node2548;
											assign node2548 = (inp[4]) ? node2554 : node2549;
												assign node2549 = (inp[12]) ? 4'b1001 : node2550;
													assign node2550 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node2554 = (inp[10]) ? node2556 : 4'b1101;
													assign node2556 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node2559 = (inp[10]) ? node2565 : node2560;
												assign node2560 = (inp[12]) ? 4'b1001 : node2561;
													assign node2561 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node2565 = (inp[4]) ? 4'b1001 : 4'b0001;
									assign node2568 = (inp[12]) ? node2588 : node2569;
										assign node2569 = (inp[10]) ? node2579 : node2570;
											assign node2570 = (inp[7]) ? node2574 : node2571;
												assign node2571 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node2574 = (inp[4]) ? node2576 : 4'b1110;
													assign node2576 = (inp[11]) ? 4'b0101 : 4'b0000;
											assign node2579 = (inp[11]) ? 4'b1001 : node2580;
												assign node2580 = (inp[14]) ? node2584 : node2581;
													assign node2581 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node2584 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node2588 = (inp[14]) ? node2594 : node2589;
											assign node2589 = (inp[3]) ? node2591 : 4'b0001;
												assign node2591 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node2594 = (inp[11]) ? node2600 : node2595;
												assign node2595 = (inp[3]) ? 4'b0100 : node2596;
													assign node2596 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node2600 = (inp[3]) ? 4'b0101 : 4'b0001;
								assign node2603 = (inp[14]) ? node2639 : node2604;
									assign node2604 = (inp[13]) ? node2622 : node2605;
										assign node2605 = (inp[11]) ? node2615 : node2606;
											assign node2606 = (inp[4]) ? 4'b0100 : node2607;
												assign node2607 = (inp[12]) ? node2611 : node2608;
													assign node2608 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node2611 = (inp[5]) ? 4'b0100 : 4'b0000;
											assign node2615 = (inp[10]) ? node2617 : 4'b0100;
												assign node2617 = (inp[4]) ? node2619 : 4'b0000;
													assign node2619 = (inp[3]) ? 4'b0100 : 4'b0000;
										assign node2622 = (inp[12]) ? node2628 : node2623;
											assign node2623 = (inp[4]) ? node2625 : 4'b1000;
												assign node2625 = (inp[3]) ? 4'b1100 : 4'b1000;
											assign node2628 = (inp[10]) ? node2634 : node2629;
												assign node2629 = (inp[11]) ? 4'b0100 : node2630;
													assign node2630 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node2634 = (inp[3]) ? node2636 : 4'b1110;
													assign node2636 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node2639 = (inp[11]) ? node2655 : node2640;
										assign node2640 = (inp[13]) ? node2648 : node2641;
											assign node2641 = (inp[12]) ? node2643 : 4'b0101;
												assign node2643 = (inp[3]) ? node2645 : 4'b1110;
													assign node2645 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node2648 = (inp[10]) ? node2652 : node2649;
												assign node2649 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node2652 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2655 = (inp[3]) ? node2661 : node2656;
											assign node2656 = (inp[5]) ? node2658 : 4'b0000;
												assign node2658 = (inp[10]) ? 4'b1000 : 4'b0100;
											assign node2661 = (inp[13]) ? node2663 : 4'b0100;
												assign node2663 = (inp[7]) ? 4'b1000 : 4'b0100;
							assign node2666 = (inp[5]) ? node2668 : 4'b1110;
								assign node2668 = (inp[3]) ? node2692 : node2669;
									assign node2669 = (inp[7]) ? node2685 : node2670;
										assign node2670 = (inp[13]) ? node2676 : node2671;
											assign node2671 = (inp[11]) ? node2673 : 4'b1110;
												assign node2673 = (inp[1]) ? 4'b0000 : 4'b1001;
											assign node2676 = (inp[4]) ? node2678 : 4'b0001;
												assign node2678 = (inp[1]) ? node2682 : node2679;
													assign node2679 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2682 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node2685 = (inp[4]) ? node2687 : 4'b1110;
											assign node2687 = (inp[14]) ? node2689 : 4'b0000;
												assign node2689 = (inp[12]) ? 4'b1110 : 4'b1000;
									assign node2692 = (inp[1]) ? node2708 : node2693;
										assign node2693 = (inp[13]) ? node2705 : node2694;
											assign node2694 = (inp[12]) ? node2700 : node2695;
												assign node2695 = (inp[14]) ? 4'b1101 : node2696;
													assign node2696 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node2700 = (inp[4]) ? node2702 : 4'b1001;
													assign node2702 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node2705 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node2708 = (inp[11]) ? node2722 : node2709;
											assign node2709 = (inp[14]) ? node2717 : node2710;
												assign node2710 = (inp[7]) ? node2714 : node2711;
													assign node2711 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node2714 = (inp[4]) ? 4'b0100 : 4'b1000;
												assign node2717 = (inp[4]) ? node2719 : 4'b1001;
													assign node2719 = (inp[7]) ? 4'b0101 : 4'b1101;
											assign node2722 = (inp[4]) ? 4'b0100 : node2723;
												assign node2723 = (inp[7]) ? 4'b0000 : 4'b0100;
					assign node2728 = (inp[0]) ? 4'b1000 : node2729;
						assign node2729 = (inp[2]) ? node2839 : node2730;
							assign node2730 = (inp[5]) ? node2760 : node2731;
								assign node2731 = (inp[3]) ? node2733 : 4'b1010;
									assign node2733 = (inp[7]) ? node2751 : node2734;
										assign node2734 = (inp[11]) ? node2740 : node2735;
											assign node2735 = (inp[10]) ? node2737 : 4'b0000;
												assign node2737 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node2740 = (inp[1]) ? node2746 : node2741;
												assign node2741 = (inp[4]) ? node2743 : 4'b0001;
													assign node2743 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node2746 = (inp[12]) ? 4'b0000 : node2747;
													assign node2747 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node2751 = (inp[4]) ? node2753 : 4'b1010;
											assign node2753 = (inp[14]) ? node2757 : node2754;
												assign node2754 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node2757 = (inp[13]) ? 4'b1000 : 4'b1010;
								assign node2760 = (inp[12]) ? node2804 : node2761;
									assign node2761 = (inp[13]) ? node2779 : node2762;
										assign node2762 = (inp[10]) ? node2772 : node2763;
											assign node2763 = (inp[14]) ? node2765 : 4'b1001;
												assign node2765 = (inp[4]) ? node2769 : node2766;
													assign node2766 = (inp[11]) ? 4'b1101 : 4'b1000;
													assign node2769 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node2772 = (inp[1]) ? node2774 : 4'b0100;
												assign node2774 = (inp[7]) ? node2776 : 4'b0101;
													assign node2776 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node2779 = (inp[1]) ? node2795 : node2780;
											assign node2780 = (inp[14]) ? node2788 : node2781;
												assign node2781 = (inp[10]) ? node2785 : node2782;
													assign node2782 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node2785 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node2788 = (inp[10]) ? node2792 : node2789;
													assign node2789 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node2792 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node2795 = (inp[14]) ? node2801 : node2796;
												assign node2796 = (inp[11]) ? 4'b1100 : node2797;
													assign node2797 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node2801 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node2804 = (inp[13]) ? node2822 : node2805;
										assign node2805 = (inp[1]) ? node2815 : node2806;
											assign node2806 = (inp[4]) ? node2810 : node2807;
												assign node2807 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node2810 = (inp[11]) ? node2812 : 4'b1101;
													assign node2812 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node2815 = (inp[11]) ? node2819 : node2816;
												assign node2816 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node2819 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node2822 = (inp[3]) ? node2830 : node2823;
											assign node2823 = (inp[1]) ? node2825 : 4'b0101;
												assign node2825 = (inp[14]) ? 4'b0101 : node2826;
													assign node2826 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node2830 = (inp[7]) ? node2836 : node2831;
												assign node2831 = (inp[14]) ? 4'b0001 : node2832;
													assign node2832 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node2836 = (inp[10]) ? 4'b0101 : 4'b0001;
							assign node2839 = (inp[3]) ? node2841 : 4'b1010;
								assign node2841 = (inp[5]) ? node2843 : 4'b1010;
									assign node2843 = (inp[4]) ? node2847 : node2844;
										assign node2844 = (inp[7]) ? 4'b1010 : 4'b0001;
										assign node2847 = (inp[13]) ? node2855 : node2848;
											assign node2848 = (inp[12]) ? node2852 : node2849;
												assign node2849 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node2852 = (inp[7]) ? 4'b1010 : 4'b1001;
											assign node2855 = (inp[12]) ? node2861 : node2856;
												assign node2856 = (inp[10]) ? node2858 : 4'b0001;
													assign node2858 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node2861 = (inp[11]) ? 4'b0001 : 4'b0000;
				assign node2865 = (inp[5]) ? node3269 : node2866;
					assign node2866 = (inp[0]) ? node3162 : node2867;
						assign node2867 = (inp[11]) ? node3025 : node2868;
							assign node2868 = (inp[3]) ? node2952 : node2869;
								assign node2869 = (inp[15]) ? node2911 : node2870;
									assign node2870 = (inp[13]) ? node2890 : node2871;
										assign node2871 = (inp[10]) ? node2877 : node2872;
											assign node2872 = (inp[12]) ? node2874 : 4'b1100;
												assign node2874 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node2877 = (inp[12]) ? node2885 : node2878;
												assign node2878 = (inp[2]) ? node2882 : node2879;
													assign node2879 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node2882 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node2885 = (inp[14]) ? node2887 : 4'b0100;
													assign node2887 = (inp[2]) ? 4'b1100 : 4'b0001;
										assign node2890 = (inp[12]) ? node2898 : node2891;
											assign node2891 = (inp[14]) ? 4'b1101 : node2892;
												assign node2892 = (inp[7]) ? node2894 : 4'b0001;
													assign node2894 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node2898 = (inp[2]) ? node2904 : node2899;
												assign node2899 = (inp[4]) ? 4'b0101 : node2900;
													assign node2900 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node2904 = (inp[4]) ? node2908 : node2905;
													assign node2905 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2908 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node2911 = (inp[7]) ? node2931 : node2912;
										assign node2912 = (inp[2]) ? node2918 : node2913;
											assign node2913 = (inp[4]) ? node2915 : 4'b1100;
												assign node2915 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node2918 = (inp[12]) ? node2924 : node2919;
												assign node2919 = (inp[1]) ? node2921 : 4'b0100;
													assign node2921 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node2924 = (inp[13]) ? node2928 : node2925;
													assign node2925 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2928 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node2931 = (inp[1]) ? node2939 : node2932;
											assign node2932 = (inp[14]) ? node2934 : 4'b1001;
												assign node2934 = (inp[13]) ? 4'b0000 : node2935;
													assign node2935 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node2939 = (inp[14]) ? node2947 : node2940;
												assign node2940 = (inp[4]) ? node2944 : node2941;
													assign node2941 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node2944 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node2947 = (inp[10]) ? 4'b0001 : node2948;
													assign node2948 = (inp[13]) ? 4'b0001 : 4'b1001;
								assign node2952 = (inp[10]) ? node2982 : node2953;
									assign node2953 = (inp[12]) ? node2971 : node2954;
										assign node2954 = (inp[1]) ? node2964 : node2955;
											assign node2955 = (inp[4]) ? node2961 : node2956;
												assign node2956 = (inp[15]) ? 4'b1101 : node2957;
													assign node2957 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node2961 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node2964 = (inp[2]) ? 4'b0001 : node2965;
												assign node2965 = (inp[13]) ? node2967 : 4'b0001;
													assign node2967 = (inp[15]) ? 4'b1001 : 4'b0001;
										assign node2971 = (inp[7]) ? node2977 : node2972;
											assign node2972 = (inp[2]) ? node2974 : 4'b1101;
												assign node2974 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node2977 = (inp[13]) ? 4'b0000 : node2978;
												assign node2978 = (inp[2]) ? 4'b1100 : 4'b1001;
									assign node2982 = (inp[12]) ? node3008 : node2983;
										assign node2983 = (inp[1]) ? node2999 : node2984;
											assign node2984 = (inp[2]) ? node2992 : node2985;
												assign node2985 = (inp[14]) ? node2989 : node2986;
													assign node2986 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node2989 = (inp[15]) ? 4'b0001 : 4'b1001;
												assign node2992 = (inp[7]) ? node2996 : node2993;
													assign node2993 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node2996 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node2999 = (inp[13]) ? node3005 : node3000;
												assign node3000 = (inp[4]) ? 4'b0000 : node3001;
													assign node3001 = (inp[2]) ? 4'b0000 : 4'b1001;
												assign node3005 = (inp[14]) ? 4'b1001 : 4'b1101;
										assign node3008 = (inp[15]) ? node3018 : node3009;
											assign node3009 = (inp[13]) ? node3015 : node3010;
												assign node3010 = (inp[14]) ? node3012 : 4'b1001;
													assign node3012 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node3015 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node3018 = (inp[2]) ? node3020 : 4'b0101;
												assign node3020 = (inp[7]) ? node3022 : 4'b0001;
													assign node3022 = (inp[14]) ? 4'b0101 : 4'b0100;
							assign node3025 = (inp[1]) ? node3101 : node3026;
								assign node3026 = (inp[2]) ? node3060 : node3027;
									assign node3027 = (inp[7]) ? node3049 : node3028;
										assign node3028 = (inp[14]) ? node3040 : node3029;
											assign node3029 = (inp[3]) ? node3033 : node3030;
												assign node3030 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node3033 = (inp[13]) ? node3037 : node3034;
													assign node3034 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node3037 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node3040 = (inp[10]) ? node3046 : node3041;
												assign node3041 = (inp[13]) ? 4'b0000 : node3042;
													assign node3042 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node3046 = (inp[12]) ? 4'b0100 : 4'b1000;
										assign node3049 = (inp[4]) ? node3057 : node3050;
											assign node3050 = (inp[3]) ? node3052 : 4'b1000;
												assign node3052 = (inp[12]) ? 4'b0000 : node3053;
													assign node3053 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node3057 = (inp[13]) ? 4'b0000 : 4'b1001;
									assign node3060 = (inp[3]) ? node3080 : node3061;
										assign node3061 = (inp[7]) ? node3071 : node3062;
											assign node3062 = (inp[15]) ? node3068 : node3063;
												assign node3063 = (inp[12]) ? 4'b0001 : node3064;
													assign node3064 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node3068 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node3071 = (inp[15]) ? node3077 : node3072;
												assign node3072 = (inp[14]) ? 4'b0101 : node3073;
													assign node3073 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node3077 = (inp[13]) ? 4'b0101 : 4'b1001;
										assign node3080 = (inp[15]) ? node3094 : node3081;
											assign node3081 = (inp[12]) ? node3089 : node3082;
												assign node3082 = (inp[4]) ? node3086 : node3083;
													assign node3083 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3086 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node3089 = (inp[13]) ? 4'b0001 : node3090;
													assign node3090 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node3094 = (inp[4]) ? 4'b0000 : node3095;
												assign node3095 = (inp[12]) ? 4'b1101 : node3096;
													assign node3096 = (inp[13]) ? 4'b0101 : 4'b0101;
								assign node3101 = (inp[10]) ? node3127 : node3102;
									assign node3102 = (inp[13]) ? node3110 : node3103;
										assign node3103 = (inp[3]) ? node3107 : node3104;
											assign node3104 = (inp[14]) ? 4'b0100 : 4'b0000;
											assign node3107 = (inp[15]) ? 4'b0000 : 4'b1000;
										assign node3110 = (inp[12]) ? node3116 : node3111;
											assign node3111 = (inp[15]) ? node3113 : 4'b0000;
												assign node3113 = (inp[4]) ? 4'b0000 : 4'b1100;
											assign node3116 = (inp[2]) ? node3122 : node3117;
												assign node3117 = (inp[15]) ? node3119 : 4'b1100;
													assign node3119 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node3122 = (inp[3]) ? node3124 : 4'b0100;
													assign node3124 = (inp[4]) ? 4'b0000 : 4'b0000;
									assign node3127 = (inp[13]) ? node3149 : node3128;
										assign node3128 = (inp[7]) ? node3140 : node3129;
											assign node3129 = (inp[14]) ? node3133 : node3130;
												assign node3130 = (inp[3]) ? 4'b1100 : 4'b0100;
												assign node3133 = (inp[3]) ? node3137 : node3134;
													assign node3134 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node3137 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node3140 = (inp[4]) ? node3146 : node3141;
												assign node3141 = (inp[3]) ? node3143 : 4'b0100;
													assign node3143 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node3146 = (inp[12]) ? 4'b1000 : 4'b0100;
										assign node3149 = (inp[2]) ? node3155 : node3150;
											assign node3150 = (inp[3]) ? 4'b1100 : node3151;
												assign node3151 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node3155 = (inp[3]) ? 4'b1000 : node3156;
												assign node3156 = (inp[4]) ? 4'b1100 : node3157;
													assign node3157 = (inp[14]) ? 4'b1100 : 4'b1000;
						assign node3162 = (inp[15]) ? node3228 : node3163;
							assign node3163 = (inp[2]) ? 4'b1100 : node3164;
								assign node3164 = (inp[1]) ? node3198 : node3165;
									assign node3165 = (inp[13]) ? node3187 : node3166;
										assign node3166 = (inp[12]) ? node3176 : node3167;
											assign node3167 = (inp[10]) ? node3173 : node3168;
												assign node3168 = (inp[3]) ? 4'b1001 : node3169;
													assign node3169 = (inp[4]) ? 4'b1001 : 4'b1100;
												assign node3173 = (inp[14]) ? 4'b0001 : 4'b0101;
											assign node3176 = (inp[7]) ? node3184 : node3177;
												assign node3177 = (inp[10]) ? node3181 : node3178;
													assign node3178 = (inp[11]) ? 4'b1001 : 4'b1100;
													assign node3181 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node3184 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node3187 = (inp[4]) ? node3193 : node3188;
											assign node3188 = (inp[7]) ? 4'b0000 : node3189;
												assign node3189 = (inp[3]) ? 4'b0100 : 4'b0000;
											assign node3193 = (inp[7]) ? 4'b1100 : node3194;
												assign node3194 = (inp[3]) ? 4'b0101 : 4'b0001;
									assign node3198 = (inp[14]) ? node3216 : node3199;
										assign node3199 = (inp[12]) ? node3203 : node3200;
											assign node3200 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node3203 = (inp[7]) ? node3211 : node3204;
												assign node3204 = (inp[3]) ? node3208 : node3205;
													assign node3205 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node3208 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node3211 = (inp[4]) ? 4'b0100 : node3212;
													assign node3212 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node3216 = (inp[11]) ? node3222 : node3217;
											assign node3217 = (inp[13]) ? node3219 : 4'b1001;
												assign node3219 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node3222 = (inp[7]) ? node3224 : 4'b0100;
												assign node3224 = (inp[13]) ? 4'b1000 : 4'b0000;
							assign node3228 = (inp[3]) ? node3230 : 4'b1000;
								assign node3230 = (inp[2]) ? 4'b1000 : node3231;
									assign node3231 = (inp[1]) ? node3249 : node3232;
										assign node3232 = (inp[13]) ? node3242 : node3233;
											assign node3233 = (inp[4]) ? node3235 : 4'b1000;
												assign node3235 = (inp[12]) ? node3239 : node3236;
													assign node3236 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node3239 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node3242 = (inp[11]) ? 4'b0001 : node3243;
												assign node3243 = (inp[12]) ? 4'b0001 : node3244;
													assign node3244 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node3249 = (inp[4]) ? node3259 : node3250;
											assign node3250 = (inp[10]) ? node3256 : node3251;
												assign node3251 = (inp[13]) ? node3253 : 4'b1000;
													assign node3253 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node3256 = (inp[12]) ? 4'b1000 : 4'b1001;
											assign node3259 = (inp[13]) ? 4'b1000 : node3260;
												assign node3260 = (inp[7]) ? node3264 : node3261;
													assign node3261 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node3264 = (inp[11]) ? 4'b0000 : 4'b0000;
					assign node3269 = (inp[3]) ? node3535 : node3270;
						assign node3270 = (inp[2]) ? node3428 : node3271;
							assign node3271 = (inp[11]) ? node3355 : node3272;
								assign node3272 = (inp[0]) ? node3316 : node3273;
									assign node3273 = (inp[4]) ? node3299 : node3274;
										assign node3274 = (inp[10]) ? node3286 : node3275;
											assign node3275 = (inp[12]) ? node3281 : node3276;
												assign node3276 = (inp[13]) ? 4'b1000 : node3277;
													assign node3277 = (inp[1]) ? 4'b0100 : 4'b0100;
												assign node3281 = (inp[14]) ? 4'b0101 : node3282;
													assign node3282 = (inp[1]) ? 4'b0101 : 4'b1000;
											assign node3286 = (inp[12]) ? node3292 : node3287;
												assign node3287 = (inp[1]) ? node3289 : 4'b0000;
													assign node3289 = (inp[13]) ? 4'b1000 : 4'b0101;
												assign node3292 = (inp[15]) ? node3296 : node3293;
													assign node3293 = (inp[1]) ? 4'b0000 : 4'b1100;
													assign node3296 = (inp[1]) ? 4'b1000 : 4'b1000;
										assign node3299 = (inp[10]) ? node3307 : node3300;
											assign node3300 = (inp[1]) ? node3304 : node3301;
												assign node3301 = (inp[13]) ? 4'b0101 : 4'b0000;
												assign node3304 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node3307 = (inp[7]) ? node3313 : node3308;
												assign node3308 = (inp[14]) ? 4'b0001 : node3309;
													assign node3309 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node3313 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node3316 = (inp[13]) ? node3334 : node3317;
										assign node3317 = (inp[10]) ? node3321 : node3318;
											assign node3318 = (inp[14]) ? 4'b1001 : 4'b1101;
											assign node3321 = (inp[14]) ? node3327 : node3322;
												assign node3322 = (inp[7]) ? 4'b0000 : node3323;
													assign node3323 = (inp[12]) ? 4'b0001 : 4'b0001;
												assign node3327 = (inp[4]) ? node3331 : node3328;
													assign node3328 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node3331 = (inp[1]) ? 4'b0001 : 4'b0101;
										assign node3334 = (inp[15]) ? node3346 : node3335;
											assign node3335 = (inp[7]) ? node3341 : node3336;
												assign node3336 = (inp[1]) ? node3338 : 4'b1001;
													assign node3338 = (inp[10]) ? 4'b0001 : 4'b0001;
												assign node3341 = (inp[4]) ? node3343 : 4'b0100;
													assign node3343 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node3346 = (inp[1]) ? node3352 : node3347;
												assign node3347 = (inp[14]) ? node3349 : 4'b0101;
													assign node3349 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node3352 = (inp[4]) ? 4'b0001 : 4'b1100;
								assign node3355 = (inp[1]) ? node3389 : node3356;
									assign node3356 = (inp[7]) ? node3368 : node3357;
										assign node3357 = (inp[14]) ? node3365 : node3358;
											assign node3358 = (inp[4]) ? node3360 : 4'b0000;
												assign node3360 = (inp[10]) ? 4'b0000 : node3361;
													assign node3361 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node3365 = (inp[0]) ? 4'b0000 : 4'b0100;
										assign node3368 = (inp[14]) ? node3382 : node3369;
											assign node3369 = (inp[15]) ? node3377 : node3370;
												assign node3370 = (inp[12]) ? node3374 : node3371;
													assign node3371 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node3374 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node3377 = (inp[13]) ? node3379 : 4'b1001;
													assign node3379 = (inp[12]) ? 4'b0101 : 4'b1001;
											assign node3382 = (inp[10]) ? node3386 : node3383;
												assign node3383 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node3386 = (inp[13]) ? 4'b0001 : 4'b0100;
									assign node3389 = (inp[13]) ? node3413 : node3390;
										assign node3390 = (inp[15]) ? node3400 : node3391;
											assign node3391 = (inp[10]) ? 4'b1000 : node3392;
												assign node3392 = (inp[7]) ? node3396 : node3393;
													assign node3393 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node3396 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node3400 = (inp[10]) ? node3408 : node3401;
												assign node3401 = (inp[0]) ? node3405 : node3402;
													assign node3402 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node3405 = (inp[4]) ? 4'b0000 : 4'b0000;
												assign node3408 = (inp[12]) ? 4'b0100 : node3409;
													assign node3409 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node3413 = (inp[10]) ? node3421 : node3414;
											assign node3414 = (inp[12]) ? node3416 : 4'b0000;
												assign node3416 = (inp[7]) ? 4'b0000 : node3417;
													assign node3417 = (inp[15]) ? 4'b0000 : 4'b1000;
											assign node3421 = (inp[14]) ? 4'b1000 : node3422;
												assign node3422 = (inp[0]) ? node3424 : 4'b1000;
													assign node3424 = (inp[7]) ? 4'b1000 : 4'b1100;
							assign node3428 = (inp[0]) ? node3500 : node3429;
								assign node3429 = (inp[4]) ? node3463 : node3430;
									assign node3430 = (inp[1]) ? node3450 : node3431;
										assign node3431 = (inp[10]) ? node3437 : node3432;
											assign node3432 = (inp[11]) ? 4'b0100 : node3433;
												assign node3433 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node3437 = (inp[7]) ? node3443 : node3438;
												assign node3438 = (inp[13]) ? node3440 : 4'b1001;
													assign node3440 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node3443 = (inp[11]) ? node3447 : node3444;
													assign node3444 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node3447 = (inp[12]) ? 4'b0000 : 4'b1100;
										assign node3450 = (inp[10]) ? node3452 : 4'b0100;
											assign node3452 = (inp[11]) ? node3460 : node3453;
												assign node3453 = (inp[14]) ? node3457 : node3454;
													assign node3454 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node3457 = (inp[12]) ? 4'b0000 : 4'b1100;
												assign node3460 = (inp[14]) ? 4'b1100 : 4'b1000;
									assign node3463 = (inp[7]) ? node3483 : node3464;
										assign node3464 = (inp[1]) ? node3474 : node3465;
											assign node3465 = (inp[11]) ? node3471 : node3466;
												assign node3466 = (inp[12]) ? 4'b1000 : node3467;
													assign node3467 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node3471 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node3474 = (inp[11]) ? node3478 : node3475;
												assign node3475 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node3478 = (inp[14]) ? 4'b1000 : node3479;
													assign node3479 = (inp[13]) ? 4'b1000 : 4'b0100;
										assign node3483 = (inp[13]) ? node3493 : node3484;
											assign node3484 = (inp[15]) ? node3490 : node3485;
												assign node3485 = (inp[14]) ? 4'b0101 : node3486;
													assign node3486 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node3490 = (inp[14]) ? 4'b0000 : 4'b1001;
											assign node3493 = (inp[14]) ? node3495 : 4'b0000;
												assign node3495 = (inp[12]) ? node3497 : 4'b1001;
													assign node3497 = (inp[1]) ? 4'b0000 : 4'b1000;
								assign node3500 = (inp[15]) ? 4'b1000 : node3501;
									assign node3501 = (inp[7]) ? node3521 : node3502;
										assign node3502 = (inp[1]) ? node3510 : node3503;
											assign node3503 = (inp[4]) ? 4'b1001 : node3504;
												assign node3504 = (inp[13]) ? node3506 : 4'b1100;
													assign node3506 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3510 = (inp[11]) ? node3516 : node3511;
												assign node3511 = (inp[14]) ? node3513 : 4'b0000;
													assign node3513 = (inp[13]) ? 4'b0001 : 4'b0001;
												assign node3516 = (inp[10]) ? node3518 : 4'b0000;
													assign node3518 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node3521 = (inp[4]) ? node3523 : 4'b1100;
											assign node3523 = (inp[1]) ? node3529 : node3524;
												assign node3524 = (inp[12]) ? 4'b1100 : node3525;
													assign node3525 = (inp[10]) ? 4'b0000 : 4'b1100;
												assign node3529 = (inp[11]) ? node3531 : 4'b0001;
													assign node3531 = (inp[13]) ? 4'b1000 : 4'b0000;
						assign node3535 = (inp[4]) ? node3685 : node3536;
							assign node3536 = (inp[1]) ? node3616 : node3537;
								assign node3537 = (inp[0]) ? node3579 : node3538;
									assign node3538 = (inp[12]) ? node3558 : node3539;
										assign node3539 = (inp[11]) ? node3551 : node3540;
											assign node3540 = (inp[7]) ? node3546 : node3541;
												assign node3541 = (inp[15]) ? node3543 : 4'b0001;
													assign node3543 = (inp[13]) ? 4'b1000 : 4'b0001;
												assign node3546 = (inp[13]) ? 4'b0001 : node3547;
													assign node3547 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node3551 = (inp[15]) ? 4'b0001 : node3552;
												assign node3552 = (inp[2]) ? node3554 : 4'b1001;
													assign node3554 = (inp[10]) ? 4'b0001 : 4'b0001;
										assign node3558 = (inp[14]) ? node3566 : node3559;
											assign node3559 = (inp[13]) ? node3561 : 4'b0001;
												assign node3561 = (inp[10]) ? 4'b1001 : node3562;
													assign node3562 = (inp[15]) ? 4'b1001 : 4'b0000;
											assign node3566 = (inp[10]) ? node3572 : node3567;
												assign node3567 = (inp[15]) ? node3569 : 4'b1000;
													assign node3569 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node3572 = (inp[7]) ? node3576 : node3573;
													assign node3573 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node3576 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node3579 = (inp[13]) ? node3597 : node3580;
										assign node3580 = (inp[15]) ? node3590 : node3581;
											assign node3581 = (inp[2]) ? node3587 : node3582;
												assign node3582 = (inp[11]) ? node3584 : 4'b1000;
													assign node3584 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node3587 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node3590 = (inp[2]) ? 4'b1000 : node3591;
												assign node3591 = (inp[12]) ? 4'b1001 : node3592;
													assign node3592 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node3597 = (inp[11]) ? node3609 : node3598;
											assign node3598 = (inp[10]) ? node3602 : node3599;
												assign node3599 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node3602 = (inp[7]) ? node3606 : node3603;
													assign node3603 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node3606 = (inp[12]) ? 4'b1001 : 4'b1000;
											assign node3609 = (inp[2]) ? node3611 : 4'b0000;
												assign node3611 = (inp[10]) ? 4'b0001 : node3612;
													assign node3612 = (inp[15]) ? 4'b0001 : 4'b1000;
								assign node3616 = (inp[11]) ? node3660 : node3617;
									assign node3617 = (inp[7]) ? node3639 : node3618;
										assign node3618 = (inp[2]) ? node3630 : node3619;
											assign node3619 = (inp[14]) ? node3625 : node3620;
												assign node3620 = (inp[15]) ? node3622 : 4'b0000;
													assign node3622 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node3625 = (inp[0]) ? 4'b0000 : node3626;
													assign node3626 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node3630 = (inp[15]) ? 4'b0001 : node3631;
												assign node3631 = (inp[10]) ? node3635 : node3632;
													assign node3632 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node3635 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node3639 = (inp[0]) ? node3647 : node3640;
											assign node3640 = (inp[12]) ? node3642 : 4'b1001;
												assign node3642 = (inp[10]) ? 4'b1001 : node3643;
													assign node3643 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node3647 = (inp[13]) ? node3653 : node3648;
												assign node3648 = (inp[2]) ? node3650 : 4'b0001;
													assign node3650 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node3653 = (inp[15]) ? node3657 : node3654;
													assign node3654 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3657 = (inp[10]) ? 4'b1000 : 4'b1000;
									assign node3660 = (inp[10]) ? node3676 : node3661;
										assign node3661 = (inp[7]) ? node3671 : node3662;
											assign node3662 = (inp[0]) ? node3668 : node3663;
												assign node3663 = (inp[15]) ? 4'b0000 : node3664;
													assign node3664 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node3668 = (inp[15]) ? 4'b1000 : 4'b0000;
											assign node3671 = (inp[15]) ? node3673 : 4'b0000;
												assign node3673 = (inp[0]) ? 4'b1000 : 4'b0000;
										assign node3676 = (inp[13]) ? 4'b1000 : node3677;
											assign node3677 = (inp[7]) ? 4'b1000 : node3678;
												assign node3678 = (inp[2]) ? 4'b0000 : node3679;
													assign node3679 = (inp[15]) ? 4'b0000 : 4'b1000;
							assign node3685 = (inp[13]) ? node3745 : node3686;
								assign node3686 = (inp[10]) ? node3712 : node3687;
									assign node3687 = (inp[11]) ? node3695 : node3688;
										assign node3688 = (inp[14]) ? node3690 : 4'b1000;
											assign node3690 = (inp[2]) ? 4'b0000 : node3691;
												assign node3691 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node3695 = (inp[1]) ? node3707 : node3696;
											assign node3696 = (inp[0]) ? node3700 : node3697;
												assign node3697 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node3700 = (inp[12]) ? node3704 : node3701;
													assign node3701 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3704 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node3707 = (inp[15]) ? 4'b0000 : node3708;
												assign node3708 = (inp[14]) ? 4'b1000 : 4'b0000;
									assign node3712 = (inp[11]) ? node3732 : node3713;
										assign node3713 = (inp[14]) ? node3723 : node3714;
											assign node3714 = (inp[1]) ? node3716 : 4'b0001;
												assign node3716 = (inp[15]) ? node3720 : node3717;
													assign node3717 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node3720 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node3723 = (inp[15]) ? node3727 : node3724;
												assign node3724 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node3727 = (inp[0]) ? node3729 : 4'b0000;
													assign node3729 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node3732 = (inp[1]) ? 4'b0000 : node3733;
											assign node3733 = (inp[2]) ? node3737 : node3734;
												assign node3734 = (inp[15]) ? 4'b0000 : 4'b1000;
												assign node3737 = (inp[14]) ? node3741 : node3738;
													assign node3738 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node3741 = (inp[15]) ? 4'b1000 : 4'b0000;
								assign node3745 = (inp[11]) ? node3775 : node3746;
									assign node3746 = (inp[10]) ? node3766 : node3747;
										assign node3747 = (inp[2]) ? node3757 : node3748;
											assign node3748 = (inp[12]) ? node3752 : node3749;
												assign node3749 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node3752 = (inp[7]) ? 4'b0001 : node3753;
													assign node3753 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node3757 = (inp[14]) ? node3759 : 4'b0000;
												assign node3759 = (inp[12]) ? node3763 : node3760;
													assign node3760 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node3763 = (inp[0]) ? 4'b0000 : 4'b0000;
										assign node3766 = (inp[1]) ? 4'b0000 : node3767;
											assign node3767 = (inp[14]) ? node3769 : 4'b0000;
												assign node3769 = (inp[7]) ? node3771 : 4'b0000;
													assign node3771 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node3775 = (inp[12]) ? 4'b0000 : node3776;
										assign node3776 = (inp[1]) ? 4'b0000 : node3777;
											assign node3777 = (inp[7]) ? node3779 : 4'b0000;
												assign node3779 = (inp[0]) ? 4'b0001 : node3780;
													assign node3780 = (inp[2]) ? 4'b0000 : 4'b0000;
			assign node3786 = (inp[15]) ? node4464 : node3787;
				assign node3787 = (inp[0]) ? node4279 : node3788;
					assign node3788 = (inp[6]) ? node3998 : node3789;
						assign node3789 = (inp[2]) ? node3931 : node3790;
							assign node3790 = (inp[3]) ? node3850 : node3791;
								assign node3791 = (inp[5]) ? node3805 : node3792;
									assign node3792 = (inp[7]) ? 4'b0110 : node3793;
										assign node3793 = (inp[4]) ? node3797 : node3794;
											assign node3794 = (inp[13]) ? 4'b0000 : 4'b0110;
											assign node3797 = (inp[13]) ? node3799 : 4'b0001;
												assign node3799 = (inp[12]) ? node3801 : 4'b0000;
													assign node3801 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node3805 = (inp[7]) ? node3827 : node3806;
										assign node3806 = (inp[4]) ? node3820 : node3807;
											assign node3807 = (inp[12]) ? node3813 : node3808;
												assign node3808 = (inp[10]) ? node3810 : 4'b0101;
													assign node3810 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node3813 = (inp[14]) ? node3817 : node3814;
													assign node3814 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node3817 = (inp[10]) ? 4'b1100 : 4'b1100;
											assign node3820 = (inp[11]) ? node3822 : 4'b1001;
												assign node3822 = (inp[1]) ? node3824 : 4'b1001;
													assign node3824 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node3827 = (inp[1]) ? node3839 : node3828;
											assign node3828 = (inp[14]) ? node3834 : node3829;
												assign node3829 = (inp[13]) ? node3831 : 4'b0101;
													assign node3831 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node3834 = (inp[13]) ? 4'b0001 : node3835;
													assign node3835 = (inp[4]) ? 4'b0100 : 4'b1100;
											assign node3839 = (inp[13]) ? node3843 : node3840;
												assign node3840 = (inp[11]) ? 4'b1100 : 4'b0101;
												assign node3843 = (inp[10]) ? node3847 : node3844;
													assign node3844 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node3847 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node3850 = (inp[4]) ? node3888 : node3851;
									assign node3851 = (inp[1]) ? node3869 : node3852;
										assign node3852 = (inp[13]) ? node3862 : node3853;
											assign node3853 = (inp[14]) ? node3859 : node3854;
												assign node3854 = (inp[10]) ? node3856 : 4'b0001;
													assign node3856 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3859 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node3862 = (inp[14]) ? node3866 : node3863;
												assign node3863 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node3866 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node3869 = (inp[11]) ? node3879 : node3870;
											assign node3870 = (inp[14]) ? node3874 : node3871;
												assign node3871 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3874 = (inp[7]) ? node3876 : 4'b0001;
													assign node3876 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node3879 = (inp[7]) ? node3885 : node3880;
												assign node3880 = (inp[5]) ? 4'b1000 : node3881;
													assign node3881 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node3885 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node3888 = (inp[7]) ? node3904 : node3889;
										assign node3889 = (inp[1]) ? node3897 : node3890;
											assign node3890 = (inp[14]) ? node3892 : 4'b0101;
												assign node3892 = (inp[13]) ? 4'b1101 : node3893;
													assign node3893 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node3897 = (inp[12]) ? node3899 : 4'b0100;
												assign node3899 = (inp[13]) ? 4'b1100 : node3900;
													assign node3900 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node3904 = (inp[1]) ? node3920 : node3905;
											assign node3905 = (inp[14]) ? node3913 : node3906;
												assign node3906 = (inp[5]) ? node3910 : node3907;
													assign node3907 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node3910 = (inp[10]) ? 4'b1001 : 4'b1001;
												assign node3913 = (inp[11]) ? node3917 : node3914;
													assign node3914 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node3917 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node3920 = (inp[13]) ? node3926 : node3921;
												assign node3921 = (inp[10]) ? 4'b1000 : node3922;
													assign node3922 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node3926 = (inp[12]) ? 4'b1000 : node3927;
													assign node3927 = (inp[14]) ? 4'b0000 : 4'b0100;
							assign node3931 = (inp[5]) ? node3933 : 4'b0110;
								assign node3933 = (inp[3]) ? node3961 : node3934;
									assign node3934 = (inp[7]) ? node3956 : node3935;
										assign node3935 = (inp[4]) ? node3945 : node3936;
											assign node3936 = (inp[13]) ? node3938 : 4'b0110;
												assign node3938 = (inp[10]) ? node3942 : node3939;
													assign node3939 = (inp[14]) ? 4'b0110 : 4'b0000;
													assign node3942 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node3945 = (inp[12]) ? node3951 : node3946;
												assign node3946 = (inp[10]) ? 4'b0000 : node3947;
													assign node3947 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node3951 = (inp[13]) ? node3953 : 4'b0001;
													assign node3953 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node3956 = (inp[11]) ? node3958 : 4'b0110;
											assign node3958 = (inp[12]) ? 4'b0000 : 4'b0110;
									assign node3961 = (inp[1]) ? node3981 : node3962;
										assign node3962 = (inp[14]) ? node3972 : node3963;
											assign node3963 = (inp[4]) ? node3969 : node3964;
												assign node3964 = (inp[7]) ? 4'b0001 : node3965;
													assign node3965 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node3969 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node3972 = (inp[11]) ? node3978 : node3973;
												assign node3973 = (inp[7]) ? 4'b0000 : node3974;
													assign node3974 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node3978 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node3981 = (inp[11]) ? node3991 : node3982;
											assign node3982 = (inp[14]) ? node3988 : node3983;
												assign node3983 = (inp[7]) ? 4'b1000 : node3984;
													assign node3984 = (inp[4]) ? 4'b1100 : 4'b0000;
												assign node3988 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node3991 = (inp[4]) ? node3995 : node3992;
												assign node3992 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node3995 = (inp[14]) ? 4'b0100 : 4'b1100;
						assign node3998 = (inp[3]) ? node4138 : node3999;
							assign node3999 = (inp[4]) ? node4077 : node4000;
								assign node4000 = (inp[13]) ? node4038 : node4001;
									assign node4001 = (inp[1]) ? node4017 : node4002;
										assign node4002 = (inp[12]) ? node4010 : node4003;
											assign node4003 = (inp[10]) ? node4007 : node4004;
												assign node4004 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node4007 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node4010 = (inp[2]) ? node4012 : 4'b0101;
												assign node4012 = (inp[14]) ? node4014 : 4'b0101;
													assign node4014 = (inp[5]) ? 4'b0100 : 4'b0100;
										assign node4017 = (inp[11]) ? node4031 : node4018;
											assign node4018 = (inp[12]) ? node4026 : node4019;
												assign node4019 = (inp[7]) ? node4023 : node4020;
													assign node4020 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node4023 = (inp[5]) ? 4'b1101 : 4'b0101;
												assign node4026 = (inp[14]) ? 4'b0101 : node4027;
													assign node4027 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node4031 = (inp[5]) ? node4033 : 4'b1100;
												assign node4033 = (inp[12]) ? node4035 : 4'b1000;
													assign node4035 = (inp[7]) ? 4'b0100 : 4'b0000;
									assign node4038 = (inp[1]) ? node4052 : node4039;
										assign node4039 = (inp[5]) ? node4043 : node4040;
											assign node4040 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node4043 = (inp[7]) ? node4049 : node4044;
												assign node4044 = (inp[11]) ? 4'b1100 : node4045;
													assign node4045 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node4049 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node4052 = (inp[11]) ? node4066 : node4053;
											assign node4053 = (inp[14]) ? node4061 : node4054;
												assign node4054 = (inp[5]) ? node4058 : node4055;
													assign node4055 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node4058 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node4061 = (inp[5]) ? node4063 : 4'b0001;
													assign node4063 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node4066 = (inp[10]) ? node4072 : node4067;
												assign node4067 = (inp[12]) ? 4'b0000 : node4068;
													assign node4068 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node4072 = (inp[2]) ? node4074 : 4'b0000;
													assign node4074 = (inp[12]) ? 4'b0100 : 4'b0000;
								assign node4077 = (inp[11]) ? node4105 : node4078;
									assign node4078 = (inp[5]) ? node4090 : node4079;
										assign node4079 = (inp[12]) ? node4083 : node4080;
											assign node4080 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node4083 = (inp[2]) ? node4085 : 4'b0001;
												assign node4085 = (inp[7]) ? 4'b1100 : node4086;
													assign node4086 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node4090 = (inp[10]) ? node4096 : node4091;
											assign node4091 = (inp[13]) ? node4093 : 4'b0000;
												assign node4093 = (inp[2]) ? 4'b1000 : 4'b0001;
											assign node4096 = (inp[7]) ? node4100 : node4097;
												assign node4097 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4100 = (inp[12]) ? node4102 : 4'b0101;
													assign node4102 = (inp[1]) ? 4'b0001 : 4'b1000;
									assign node4105 = (inp[1]) ? node4125 : node4106;
										assign node4106 = (inp[7]) ? node4112 : node4107;
											assign node4107 = (inp[13]) ? 4'b1000 : node4108;
												assign node4108 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node4112 = (inp[2]) ? node4118 : node4113;
												assign node4113 = (inp[12]) ? node4115 : 4'b1000;
													assign node4115 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node4118 = (inp[10]) ? node4122 : node4119;
													assign node4119 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node4122 = (inp[5]) ? 4'b0101 : 4'b0001;
										assign node4125 = (inp[10]) ? node4135 : node4126;
											assign node4126 = (inp[13]) ? node4130 : node4127;
												assign node4127 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node4130 = (inp[2]) ? node4132 : 4'b1000;
													assign node4132 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node4135 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node4138 = (inp[5]) ? node4216 : node4139;
								assign node4139 = (inp[11]) ? node4179 : node4140;
									assign node4140 = (inp[10]) ? node4158 : node4141;
										assign node4141 = (inp[1]) ? node4151 : node4142;
											assign node4142 = (inp[13]) ? node4148 : node4143;
												assign node4143 = (inp[7]) ? 4'b0001 : node4144;
													assign node4144 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node4148 = (inp[2]) ? 4'b1000 : 4'b0101;
											assign node4151 = (inp[2]) ? 4'b0001 : node4152;
												assign node4152 = (inp[12]) ? node4154 : 4'b1001;
													assign node4154 = (inp[14]) ? 4'b0100 : 4'b0001;
										assign node4158 = (inp[2]) ? node4170 : node4159;
											assign node4159 = (inp[13]) ? node4165 : node4160;
												assign node4160 = (inp[4]) ? 4'b1000 : node4161;
													assign node4161 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node4165 = (inp[1]) ? node4167 : 4'b0001;
													assign node4167 = (inp[4]) ? 4'b0100 : 4'b0001;
											assign node4170 = (inp[12]) ? node4176 : node4171;
												assign node4171 = (inp[4]) ? node4173 : 4'b1001;
													assign node4173 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node4176 = (inp[4]) ? 4'b1001 : 4'b1000;
									assign node4179 = (inp[1]) ? node4203 : node4180;
										assign node4180 = (inp[7]) ? node4194 : node4181;
											assign node4181 = (inp[14]) ? node4187 : node4182;
												assign node4182 = (inp[10]) ? 4'b0100 : node4183;
													assign node4183 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node4187 = (inp[4]) ? node4191 : node4188;
													assign node4188 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node4191 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node4194 = (inp[14]) ? node4198 : node4195;
												assign node4195 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node4198 = (inp[4]) ? 4'b0001 : node4199;
													assign node4199 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node4203 = (inp[10]) ? node4211 : node4204;
											assign node4204 = (inp[13]) ? 4'b1000 : node4205;
												assign node4205 = (inp[12]) ? 4'b0000 : node4206;
													assign node4206 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node4211 = (inp[13]) ? node4213 : 4'b1000;
												assign node4213 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node4216 = (inp[4]) ? node4262 : node4217;
									assign node4217 = (inp[2]) ? node4243 : node4218;
										assign node4218 = (inp[12]) ? node4230 : node4219;
											assign node4219 = (inp[10]) ? node4225 : node4220;
												assign node4220 = (inp[13]) ? node4222 : 4'b0001;
													assign node4222 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node4225 = (inp[11]) ? 4'b1000 : node4226;
													assign node4226 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node4230 = (inp[11]) ? node4238 : node4231;
												assign node4231 = (inp[7]) ? node4235 : node4232;
													assign node4232 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node4235 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node4238 = (inp[10]) ? node4240 : 4'b0000;
													assign node4240 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node4243 = (inp[12]) ? node4253 : node4244;
											assign node4244 = (inp[7]) ? 4'b1001 : node4245;
												assign node4245 = (inp[11]) ? node4249 : node4246;
													assign node4246 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node4249 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node4253 = (inp[1]) ? node4259 : node4254;
												assign node4254 = (inp[10]) ? node4256 : 4'b1001;
													assign node4256 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node4259 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node4262 = (inp[13]) ? node4270 : node4263;
										assign node4263 = (inp[10]) ? node4267 : node4264;
											assign node4264 = (inp[11]) ? 4'b1000 : 4'b0000;
											assign node4267 = (inp[14]) ? 4'b0001 : 4'b1000;
										assign node4270 = (inp[7]) ? 4'b0000 : node4271;
											assign node4271 = (inp[10]) ? 4'b0000 : node4272;
												assign node4272 = (inp[14]) ? node4274 : 4'b0001;
													assign node4274 = (inp[1]) ? 4'b0000 : 4'b0000;
					assign node4279 = (inp[6]) ? node4281 : 4'b0100;
						assign node4281 = (inp[5]) ? node4347 : node4282;
							assign node4282 = (inp[2]) ? 4'b0100 : node4283;
								assign node4283 = (inp[3]) ? node4313 : node4284;
									assign node4284 = (inp[7]) ? node4306 : node4285;
										assign node4285 = (inp[4]) ? node4295 : node4286;
											assign node4286 = (inp[12]) ? node4290 : node4287;
												assign node4287 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node4290 = (inp[1]) ? node4292 : 4'b0100;
													assign node4292 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node4295 = (inp[14]) ? node4301 : node4296;
												assign node4296 = (inp[1]) ? node4298 : 4'b0001;
													assign node4298 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node4301 = (inp[1]) ? 4'b1001 : node4302;
													assign node4302 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node4306 = (inp[13]) ? node4308 : 4'b0100;
											assign node4308 = (inp[4]) ? node4310 : 4'b0100;
												assign node4310 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node4313 = (inp[7]) ? node4325 : node4314;
										assign node4314 = (inp[4]) ? node4316 : 4'b1001;
											assign node4316 = (inp[11]) ? node4322 : node4317;
												assign node4317 = (inp[1]) ? 4'b1101 : node4318;
													assign node4318 = (inp[14]) ? 4'b0100 : 4'b1101;
												assign node4322 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node4325 = (inp[1]) ? node4337 : node4326;
											assign node4326 = (inp[11]) ? node4332 : node4327;
												assign node4327 = (inp[14]) ? node4329 : 4'b1001;
													assign node4329 = (inp[4]) ? 4'b1000 : 4'b0000;
												assign node4332 = (inp[14]) ? node4334 : 4'b0101;
													assign node4334 = (inp[13]) ? 4'b0001 : 4'b0001;
											assign node4337 = (inp[13]) ? node4341 : node4338;
												assign node4338 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4341 = (inp[11]) ? node4343 : 4'b1001;
													assign node4343 = (inp[4]) ? 4'b0100 : 4'b0000;
							assign node4347 = (inp[3]) ? node4395 : node4348;
								assign node4348 = (inp[7]) ? node4374 : node4349;
									assign node4349 = (inp[4]) ? node4365 : node4350;
										assign node4350 = (inp[2]) ? node4360 : node4351;
											assign node4351 = (inp[11]) ? node4357 : node4352;
												assign node4352 = (inp[10]) ? 4'b1001 : node4353;
													assign node4353 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4357 = (inp[12]) ? 4'b0000 : 4'b0101;
											assign node4360 = (inp[11]) ? 4'b0100 : node4361;
												assign node4361 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node4365 = (inp[1]) ? node4371 : node4366;
											assign node4366 = (inp[11]) ? 4'b1001 : node4367;
												assign node4367 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node4371 = (inp[11]) ? 4'b1000 : 4'b0001;
									assign node4374 = (inp[2]) ? node4388 : node4375;
										assign node4375 = (inp[4]) ? node4381 : node4376;
											assign node4376 = (inp[1]) ? node4378 : 4'b0100;
												assign node4378 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node4381 = (inp[11]) ? node4385 : node4382;
												assign node4382 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node4385 = (inp[1]) ? 4'b0000 : 4'b1000;
										assign node4388 = (inp[4]) ? node4390 : 4'b0100;
											assign node4390 = (inp[11]) ? node4392 : 4'b0100;
												assign node4392 = (inp[10]) ? 4'b0001 : 4'b0100;
								assign node4395 = (inp[1]) ? node4437 : node4396;
									assign node4396 = (inp[13]) ? node4424 : node4397;
										assign node4397 = (inp[12]) ? node4411 : node4398;
											assign node4398 = (inp[4]) ? node4406 : node4399;
												assign node4399 = (inp[10]) ? node4403 : node4400;
													assign node4400 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node4403 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node4406 = (inp[11]) ? node4408 : 4'b0001;
													assign node4408 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node4411 = (inp[4]) ? node4419 : node4412;
												assign node4412 = (inp[14]) ? node4416 : node4413;
													assign node4413 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node4416 = (inp[7]) ? 4'b0001 : 4'b0001;
												assign node4419 = (inp[14]) ? 4'b0000 : node4420;
													assign node4420 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node4424 = (inp[12]) ? node4426 : 4'b0000;
											assign node4426 = (inp[14]) ? node4432 : node4427;
												assign node4427 = (inp[10]) ? 4'b1000 : node4428;
													assign node4428 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node4432 = (inp[4]) ? node4434 : 4'b0001;
													assign node4434 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node4437 = (inp[11]) ? node4457 : node4438;
										assign node4438 = (inp[12]) ? node4448 : node4439;
											assign node4439 = (inp[10]) ? node4445 : node4440;
												assign node4440 = (inp[4]) ? 4'b1001 : node4441;
													assign node4441 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node4445 = (inp[2]) ? 4'b0001 : 4'b1001;
											assign node4448 = (inp[4]) ? node4454 : node4449;
												assign node4449 = (inp[7]) ? 4'b0000 : node4450;
													assign node4450 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node4454 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node4457 = (inp[10]) ? 4'b0000 : node4458;
											assign node4458 = (inp[13]) ? node4460 : 4'b0000;
												assign node4460 = (inp[12]) ? 4'b1000 : 4'b0000;
				assign node4464 = (inp[0]) ? node4868 : node4465;
					assign node4465 = (inp[6]) ? node4595 : node4466;
						assign node4466 = (inp[2]) ? node4576 : node4467;
							assign node4467 = (inp[5]) ? node4501 : node4468;
								assign node4468 = (inp[3]) ? node4470 : 4'b0010;
									assign node4470 = (inp[7]) ? node4492 : node4471;
										assign node4471 = (inp[4]) ? node4481 : node4472;
											assign node4472 = (inp[10]) ? node4478 : node4473;
												assign node4473 = (inp[12]) ? 4'b0010 : node4474;
													assign node4474 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node4478 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node4481 = (inp[12]) ? node4487 : node4482;
												assign node4482 = (inp[13]) ? node4484 : 4'b1000;
													assign node4484 = (inp[1]) ? 4'b0000 : 4'b0000;
												assign node4487 = (inp[10]) ? node4489 : 4'b1001;
													assign node4489 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node4492 = (inp[4]) ? node4494 : 4'b0010;
											assign node4494 = (inp[1]) ? node4496 : 4'b0010;
												assign node4496 = (inp[13]) ? node4498 : 4'b0010;
													assign node4498 = (inp[14]) ? 4'b0001 : 4'b0000;
								assign node4501 = (inp[1]) ? node4531 : node4502;
									assign node4502 = (inp[13]) ? node4518 : node4503;
										assign node4503 = (inp[10]) ? node4509 : node4504;
											assign node4504 = (inp[3]) ? node4506 : 4'b0001;
												assign node4506 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node4509 = (inp[14]) ? node4515 : node4510;
												assign node4510 = (inp[3]) ? node4512 : 4'b1001;
													assign node4512 = (inp[7]) ? 4'b1101 : 4'b0101;
												assign node4515 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node4518 = (inp[11]) ? node4524 : node4519;
											assign node4519 = (inp[10]) ? 4'b0100 : node4520;
												assign node4520 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node4524 = (inp[10]) ? node4526 : 4'b1101;
												assign node4526 = (inp[7]) ? node4528 : 4'b1001;
													assign node4528 = (inp[3]) ? 4'b1101 : 4'b1001;
									assign node4531 = (inp[14]) ? node4553 : node4532;
										assign node4532 = (inp[13]) ? node4540 : node4533;
											assign node4533 = (inp[7]) ? 4'b0000 : node4534;
												assign node4534 = (inp[10]) ? node4536 : 4'b1000;
													assign node4536 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node4540 = (inp[12]) ? node4546 : node4541;
												assign node4541 = (inp[3]) ? node4543 : 4'b0100;
													assign node4543 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node4546 = (inp[10]) ? node4550 : node4547;
													assign node4547 = (inp[11]) ? 4'b1100 : 4'b1000;
													assign node4550 = (inp[3]) ? 4'b0000 : 4'b0000;
										assign node4553 = (inp[11]) ? node4565 : node4554;
											assign node4554 = (inp[13]) ? node4558 : node4555;
												assign node4555 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node4558 = (inp[10]) ? node4562 : node4559;
													assign node4559 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4562 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node4565 = (inp[10]) ? node4571 : node4566;
												assign node4566 = (inp[7]) ? 4'b1100 : node4567;
													assign node4567 = (inp[3]) ? 4'b0000 : 4'b1000;
												assign node4571 = (inp[13]) ? node4573 : 4'b1100;
													assign node4573 = (inp[4]) ? 4'b0100 : 4'b0000;
							assign node4576 = (inp[4]) ? node4578 : 4'b0010;
								assign node4578 = (inp[3]) ? node4580 : 4'b0010;
									assign node4580 = (inp[5]) ? node4582 : 4'b0010;
										assign node4582 = (inp[7]) ? node4588 : node4583;
											assign node4583 = (inp[1]) ? node4585 : 4'b1001;
												assign node4585 = (inp[14]) ? 4'b1001 : 4'b0000;
											assign node4588 = (inp[13]) ? node4590 : 4'b0010;
												assign node4590 = (inp[1]) ? node4592 : 4'b0010;
													assign node4592 = (inp[11]) ? 4'b0000 : 4'b0000;
						assign node4595 = (inp[11]) ? node4759 : node4596;
							assign node4596 = (inp[3]) ? node4678 : node4597;
								assign node4597 = (inp[14]) ? node4639 : node4598;
									assign node4598 = (inp[1]) ? node4620 : node4599;
										assign node4599 = (inp[5]) ? node4611 : node4600;
											assign node4600 = (inp[12]) ? node4606 : node4601;
												assign node4601 = (inp[4]) ? node4603 : 4'b0101;
													assign node4603 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node4606 = (inp[13]) ? node4608 : 4'b0001;
													assign node4608 = (inp[2]) ? 4'b1001 : 4'b1001;
											assign node4611 = (inp[2]) ? node4615 : node4612;
												assign node4612 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4615 = (inp[7]) ? 4'b0101 : node4616;
													assign node4616 = (inp[4]) ? 4'b0000 : 4'b1001;
										assign node4620 = (inp[4]) ? node4630 : node4621;
											assign node4621 = (inp[5]) ? node4623 : 4'b0000;
												assign node4623 = (inp[13]) ? node4627 : node4624;
													assign node4624 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node4627 = (inp[12]) ? 4'b0101 : 4'b0000;
											assign node4630 = (inp[12]) ? node4636 : node4631;
												assign node4631 = (inp[2]) ? node4633 : 4'b0100;
													assign node4633 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node4636 = (inp[13]) ? 4'b1000 : 4'b1100;
									assign node4639 = (inp[1]) ? node4661 : node4640;
										assign node4640 = (inp[5]) ? node4654 : node4641;
											assign node4641 = (inp[13]) ? node4649 : node4642;
												assign node4642 = (inp[7]) ? node4646 : node4643;
													assign node4643 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node4646 = (inp[12]) ? 4'b0000 : 4'b0000;
												assign node4649 = (inp[10]) ? node4651 : 4'b1000;
													assign node4651 = (inp[4]) ? 4'b1001 : 4'b0100;
											assign node4654 = (inp[4]) ? node4656 : 4'b1001;
												assign node4656 = (inp[2]) ? node4658 : 4'b0000;
													assign node4658 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node4661 = (inp[2]) ? node4669 : node4662;
											assign node4662 = (inp[10]) ? node4664 : 4'b0001;
												assign node4664 = (inp[5]) ? node4666 : 4'b1001;
													assign node4666 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node4669 = (inp[10]) ? node4675 : node4670;
												assign node4670 = (inp[7]) ? node4672 : 4'b0001;
													assign node4672 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node4675 = (inp[4]) ? 4'b0000 : 4'b1101;
								assign node4678 = (inp[5]) ? node4720 : node4679;
									assign node4679 = (inp[7]) ? node4699 : node4680;
										assign node4680 = (inp[13]) ? node4692 : node4681;
											assign node4681 = (inp[4]) ? node4687 : node4682;
												assign node4682 = (inp[14]) ? node4684 : 4'b1100;
													assign node4684 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node4687 = (inp[1]) ? node4689 : 4'b1001;
													assign node4689 = (inp[14]) ? 4'b0001 : 4'b0101;
											assign node4692 = (inp[10]) ? node4694 : 4'b0001;
												assign node4694 = (inp[1]) ? node4696 : 4'b1000;
													assign node4696 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node4699 = (inp[2]) ? node4707 : node4700;
											assign node4700 = (inp[4]) ? 4'b1101 : node4701;
												assign node4701 = (inp[13]) ? node4703 : 4'b1001;
													assign node4703 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node4707 = (inp[13]) ? node4713 : node4708;
												assign node4708 = (inp[10]) ? 4'b1100 : node4709;
													assign node4709 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node4713 = (inp[10]) ? node4717 : node4714;
													assign node4714 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node4717 = (inp[12]) ? 4'b0100 : 4'b0001;
									assign node4720 = (inp[4]) ? node4736 : node4721;
										assign node4721 = (inp[10]) ? node4731 : node4722;
											assign node4722 = (inp[13]) ? 4'b0001 : node4723;
												assign node4723 = (inp[2]) ? node4727 : node4724;
													assign node4724 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node4727 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node4731 = (inp[2]) ? 4'b0001 : node4732;
												assign node4732 = (inp[1]) ? 4'b1000 : 4'b0001;
										assign node4736 = (inp[7]) ? node4746 : node4737;
											assign node4737 = (inp[1]) ? node4743 : node4738;
												assign node4738 = (inp[12]) ? node4740 : 4'b0001;
													assign node4740 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node4743 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node4746 = (inp[10]) ? node4752 : node4747;
												assign node4747 = (inp[13]) ? node4749 : 4'b1000;
													assign node4749 = (inp[12]) ? 4'b0000 : 4'b0000;
												assign node4752 = (inp[13]) ? node4756 : node4753;
													assign node4753 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4756 = (inp[1]) ? 4'b0000 : 4'b0000;
							assign node4759 = (inp[1]) ? node4821 : node4760;
								assign node4760 = (inp[3]) ? node4790 : node4761;
									assign node4761 = (inp[4]) ? node4779 : node4762;
										assign node4762 = (inp[5]) ? node4770 : node4763;
											assign node4763 = (inp[13]) ? node4765 : 4'b0001;
												assign node4765 = (inp[10]) ? node4767 : 4'b1001;
													assign node4767 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node4770 = (inp[2]) ? node4776 : node4771;
												assign node4771 = (inp[10]) ? 4'b1000 : node4772;
													assign node4772 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node4776 = (inp[10]) ? 4'b0100 : 4'b1000;
										assign node4779 = (inp[7]) ? node4787 : node4780;
											assign node4780 = (inp[12]) ? node4784 : node4781;
												assign node4781 = (inp[14]) ? 4'b0101 : 4'b1101;
												assign node4784 = (inp[5]) ? 4'b0001 : 4'b0101;
											assign node4787 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node4790 = (inp[5]) ? node4810 : node4791;
										assign node4791 = (inp[2]) ? node4799 : node4792;
											assign node4792 = (inp[7]) ? 4'b0100 : node4793;
												assign node4793 = (inp[10]) ? node4795 : 4'b1100;
													assign node4795 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node4799 = (inp[4]) ? node4805 : node4800;
												assign node4800 = (inp[13]) ? 4'b0001 : node4801;
													assign node4801 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node4805 = (inp[10]) ? 4'b0000 : node4806;
													assign node4806 = (inp[7]) ? 4'b1101 : 4'b0000;
										assign node4810 = (inp[14]) ? node4814 : node4811;
											assign node4811 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node4814 = (inp[12]) ? 4'b0000 : node4815;
												assign node4815 = (inp[4]) ? 4'b0000 : node4816;
													assign node4816 = (inp[2]) ? 4'b0001 : 4'b1001;
								assign node4821 = (inp[5]) ? node4847 : node4822;
									assign node4822 = (inp[14]) ? node4830 : node4823;
										assign node4823 = (inp[4]) ? 4'b0000 : node4824;
											assign node4824 = (inp[3]) ? 4'b0100 : node4825;
												assign node4825 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node4830 = (inp[10]) ? node4836 : node4831;
											assign node4831 = (inp[12]) ? 4'b0100 : node4832;
												assign node4832 = (inp[13]) ? 4'b1000 : 4'b1100;
											assign node4836 = (inp[12]) ? node4842 : node4837;
												assign node4837 = (inp[2]) ? 4'b0100 : node4838;
													assign node4838 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node4842 = (inp[3]) ? node4844 : 4'b1000;
													assign node4844 = (inp[2]) ? 4'b0000 : 4'b0000;
									assign node4847 = (inp[4]) ? node4863 : node4848;
										assign node4848 = (inp[14]) ? node4860 : node4849;
											assign node4849 = (inp[3]) ? node4855 : node4850;
												assign node4850 = (inp[2]) ? 4'b1000 : node4851;
													assign node4851 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node4855 = (inp[12]) ? 4'b0000 : node4856;
													assign node4856 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node4860 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node4863 = (inp[12]) ? node4865 : 4'b0000;
											assign node4865 = (inp[7]) ? 4'b0000 : 4'b1000;
					assign node4868 = (inp[6]) ? node4870 : 4'b0000;
						assign node4870 = (inp[2]) ? node4954 : node4871;
							assign node4871 = (inp[5]) ? node4897 : node4872;
								assign node4872 = (inp[3]) ? node4874 : 4'b0000;
									assign node4874 = (inp[7]) ? 4'b0000 : node4875;
										assign node4875 = (inp[4]) ? node4883 : node4876;
											assign node4876 = (inp[12]) ? 4'b0000 : node4877;
												assign node4877 = (inp[14]) ? node4879 : 4'b0000;
													assign node4879 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node4883 = (inp[10]) ? node4891 : node4884;
												assign node4884 = (inp[1]) ? node4888 : node4885;
													assign node4885 = (inp[13]) ? 4'b1000 : 4'b0001;
													assign node4888 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node4891 = (inp[12]) ? node4893 : 4'b0001;
													assign node4893 = (inp[13]) ? 4'b1001 : 4'b0001;
								assign node4897 = (inp[3]) ? node4927 : node4898;
									assign node4898 = (inp[7]) ? node4912 : node4899;
										assign node4899 = (inp[1]) ? node4909 : node4900;
											assign node4900 = (inp[14]) ? node4906 : node4901;
												assign node4901 = (inp[4]) ? 4'b1001 : node4902;
													assign node4902 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node4906 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node4909 = (inp[11]) ? 4'b0000 : 4'b0101;
										assign node4912 = (inp[10]) ? node4920 : node4913;
											assign node4913 = (inp[11]) ? node4917 : node4914;
												assign node4914 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node4917 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node4920 = (inp[4]) ? 4'b0000 : node4921;
												assign node4921 = (inp[12]) ? node4923 : 4'b1001;
													assign node4923 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node4927 = (inp[10]) ? node4941 : node4928;
										assign node4928 = (inp[4]) ? node4932 : node4929;
											assign node4929 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node4932 = (inp[1]) ? 4'b0000 : node4933;
												assign node4933 = (inp[13]) ? node4937 : node4934;
													assign node4934 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node4937 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node4941 = (inp[13]) ? node4949 : node4942;
											assign node4942 = (inp[1]) ? node4944 : 4'b1000;
												assign node4944 = (inp[4]) ? 4'b0000 : node4945;
													assign node4945 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node4949 = (inp[7]) ? node4951 : 4'b0000;
												assign node4951 = (inp[4]) ? 4'b0000 : 4'b1000;
							assign node4954 = (inp[4]) ? node4956 : 4'b0000;
								assign node4956 = (inp[5]) ? node4958 : 4'b0000;
									assign node4958 = (inp[3]) ? node4960 : 4'b0000;
										assign node4960 = (inp[7]) ? node4968 : node4961;
											assign node4961 = (inp[12]) ? node4963 : 4'b0001;
												assign node4963 = (inp[11]) ? node4965 : 4'b0000;
													assign node4965 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node4968 = (inp[13]) ? node4970 : 4'b0000;
												assign node4970 = (inp[1]) ? 4'b0000 : 4'b0001;

endmodule