module dtc_split875_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node8;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node15;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node23;
	wire [14-1:0] node26;
	wire [14-1:0] node27;
	wire [14-1:0] node30;
	wire [14-1:0] node33;
	wire [14-1:0] node34;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node39;
	wire [14-1:0] node42;
	wire [14-1:0] node43;
	wire [14-1:0] node46;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node54;
	wire [14-1:0] node57;
	wire [14-1:0] node58;
	wire [14-1:0] node61;
	wire [14-1:0] node64;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node71;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node78;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node86;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node93;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node102;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node109;
	wire [14-1:0] node112;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node117;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node124;

	assign outp = (inp[8]) ? node64 : node1;
		assign node1 = (inp[3]) ? node33 : node2;
			assign node2 = (inp[13]) ? node18 : node3;
				assign node3 = (inp[9]) ? node11 : node4;
					assign node4 = (inp[6]) ? node8 : node5;
						assign node5 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
						assign node8 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
					assign node11 = (inp[2]) ? node15 : node12;
						assign node12 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node15 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
				assign node18 = (inp[9]) ? node26 : node19;
					assign node19 = (inp[1]) ? node23 : node20;
						assign node20 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node23 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
					assign node26 = (inp[10]) ? node30 : node27;
						assign node27 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node30 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
			assign node33 = (inp[5]) ? node49 : node34;
				assign node34 = (inp[13]) ? node42 : node35;
					assign node35 = (inp[12]) ? node39 : node36;
						assign node36 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node39 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
					assign node42 = (inp[0]) ? node46 : node43;
						assign node43 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node46 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
				assign node49 = (inp[6]) ? node57 : node50;
					assign node50 = (inp[12]) ? node54 : node51;
						assign node51 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node54 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node57 = (inp[4]) ? node61 : node58;
						assign node58 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node61 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
		assign node64 = (inp[12]) ? node96 : node65;
			assign node65 = (inp[2]) ? node81 : node66;
				assign node66 = (inp[9]) ? node74 : node67;
					assign node67 = (inp[13]) ? node71 : node68;
						assign node68 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node71 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
					assign node74 = (inp[7]) ? node78 : node75;
						assign node75 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node78 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
				assign node81 = (inp[4]) ? node89 : node82;
					assign node82 = (inp[5]) ? node86 : node83;
						assign node83 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node86 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node89 = (inp[9]) ? node93 : node90;
						assign node90 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node93 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
			assign node96 = (inp[6]) ? node112 : node97;
				assign node97 = (inp[3]) ? node105 : node98;
					assign node98 = (inp[7]) ? node102 : node99;
						assign node99 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node102 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node105 = (inp[4]) ? node109 : node106;
						assign node106 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node109 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
				assign node112 = (inp[13]) ? node120 : node113;
					assign node113 = (inp[10]) ? node117 : node114;
						assign node114 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node117 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node120 = (inp[4]) ? node124 : node121;
						assign node121 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node124 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;

endmodule