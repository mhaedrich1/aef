module dtc_split66_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node13;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node69;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node107;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node122;
	wire [1-1:0] node124;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node131;
	wire [1-1:0] node134;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node145;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node162;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node171;
	wire [1-1:0] node173;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node187;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node194;
	wire [1-1:0] node197;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node211;
	wire [1-1:0] node212;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node226;
	wire [1-1:0] node230;
	wire [1-1:0] node232;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node249;
	wire [1-1:0] node251;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node259;
	wire [1-1:0] node262;
	wire [1-1:0] node264;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node269;
	wire [1-1:0] node272;
	wire [1-1:0] node273;
	wire [1-1:0] node277;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node283;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node292;
	wire [1-1:0] node294;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node308;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node332;
	wire [1-1:0] node334;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node342;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node355;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node365;
	wire [1-1:0] node366;
	wire [1-1:0] node370;
	wire [1-1:0] node372;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node390;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node400;
	wire [1-1:0] node403;
	wire [1-1:0] node405;
	wire [1-1:0] node406;
	wire [1-1:0] node408;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node421;
	wire [1-1:0] node425;
	wire [1-1:0] node427;
	wire [1-1:0] node428;
	wire [1-1:0] node430;
	wire [1-1:0] node434;
	wire [1-1:0] node436;
	wire [1-1:0] node438;
	wire [1-1:0] node440;
	wire [1-1:0] node441;
	wire [1-1:0] node444;
	wire [1-1:0] node447;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node454;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node462;
	wire [1-1:0] node463;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node474;
	wire [1-1:0] node476;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node484;
	wire [1-1:0] node485;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node499;
	wire [1-1:0] node501;
	wire [1-1:0] node505;
	wire [1-1:0] node506;
	wire [1-1:0] node507;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node519;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node528;
	wire [1-1:0] node531;
	wire [1-1:0] node533;
	wire [1-1:0] node535;
	wire [1-1:0] node539;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node548;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node555;
	wire [1-1:0] node558;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node564;
	wire [1-1:0] node565;
	wire [1-1:0] node567;
	wire [1-1:0] node570;
	wire [1-1:0] node571;
	wire [1-1:0] node575;
	wire [1-1:0] node577;
	wire [1-1:0] node580;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node585;
	wire [1-1:0] node588;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node594;
	wire [1-1:0] node597;
	wire [1-1:0] node599;
	wire [1-1:0] node600;
	wire [1-1:0] node601;
	wire [1-1:0] node603;
	wire [1-1:0] node606;
	wire [1-1:0] node607;
	wire [1-1:0] node609;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node618;
	wire [1-1:0] node619;
	wire [1-1:0] node620;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node630;
	wire [1-1:0] node632;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node646;
	wire [1-1:0] node650;
	wire [1-1:0] node652;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node663;
	wire [1-1:0] node664;
	wire [1-1:0] node665;
	wire [1-1:0] node669;
	wire [1-1:0] node671;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node706;
	wire [1-1:0] node707;
	wire [1-1:0] node708;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node718;
	wire [1-1:0] node719;
	wire [1-1:0] node720;
	wire [1-1:0] node721;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node731;
	wire [1-1:0] node733;
	wire [1-1:0] node736;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node747;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node755;
	wire [1-1:0] node756;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node761;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node770;
	wire [1-1:0] node771;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node779;
	wire [1-1:0] node780;
	wire [1-1:0] node781;
	wire [1-1:0] node783;
	wire [1-1:0] node786;
	wire [1-1:0] node787;
	wire [1-1:0] node789;
	wire [1-1:0] node792;
	wire [1-1:0] node793;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node807;
	wire [1-1:0] node809;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node817;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node825;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node831;
	wire [1-1:0] node832;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node843;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node851;
	wire [1-1:0] node852;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node861;
	wire [1-1:0] node862;
	wire [1-1:0] node863;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node867;
	wire [1-1:0] node869;
	wire [1-1:0] node872;
	wire [1-1:0] node873;
	wire [1-1:0] node875;
	wire [1-1:0] node878;
	wire [1-1:0] node880;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node886;
	wire [1-1:0] node887;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node894;
	wire [1-1:0] node895;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node905;
	wire [1-1:0] node906;
	wire [1-1:0] node907;
	wire [1-1:0] node908;
	wire [1-1:0] node912;
	wire [1-1:0] node914;
	wire [1-1:0] node917;
	wire [1-1:0] node918;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node925;
	wire [1-1:0] node926;
	wire [1-1:0] node927;
	wire [1-1:0] node929;
	wire [1-1:0] node932;
	wire [1-1:0] node935;
	wire [1-1:0] node937;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node947;
	wire [1-1:0] node948;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node955;
	wire [1-1:0] node956;
	wire [1-1:0] node959;
	wire [1-1:0] node962;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node968;
	wire [1-1:0] node972;
	wire [1-1:0] node973;
	wire [1-1:0] node974;
	wire [1-1:0] node975;
	wire [1-1:0] node978;
	wire [1-1:0] node980;
	wire [1-1:0] node983;
	wire [1-1:0] node984;
	wire [1-1:0] node985;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node991;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node1001;
	wire [1-1:0] node1002;
	wire [1-1:0] node1006;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1011;
	wire [1-1:0] node1015;
	wire [1-1:0] node1017;
	wire [1-1:0] node1019;
	wire [1-1:0] node1023;
	wire [1-1:0] node1024;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1028;
	wire [1-1:0] node1029;
	wire [1-1:0] node1031;
	wire [1-1:0] node1034;
	wire [1-1:0] node1036;
	wire [1-1:0] node1039;
	wire [1-1:0] node1041;
	wire [1-1:0] node1045;
	wire [1-1:0] node1046;
	wire [1-1:0] node1047;
	wire [1-1:0] node1048;
	wire [1-1:0] node1049;
	wire [1-1:0] node1053;
	wire [1-1:0] node1055;
	wire [1-1:0] node1058;
	wire [1-1:0] node1059;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1066;
	wire [1-1:0] node1071;
	wire [1-1:0] node1072;
	wire [1-1:0] node1073;
	wire [1-1:0] node1074;
	wire [1-1:0] node1078;
	wire [1-1:0] node1080;
	wire [1-1:0] node1083;
	wire [1-1:0] node1085;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1091;
	wire [1-1:0] node1093;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1099;
	wire [1-1:0] node1100;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1105;
	wire [1-1:0] node1109;
	wire [1-1:0] node1112;
	wire [1-1:0] node1114;
	wire [1-1:0] node1118;
	wire [1-1:0] node1119;
	wire [1-1:0] node1120;
	wire [1-1:0] node1122;
	wire [1-1:0] node1125;
	wire [1-1:0] node1126;
	wire [1-1:0] node1128;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1136;
	wire [1-1:0] node1138;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1144;
	wire [1-1:0] node1145;
	wire [1-1:0] node1147;
	wire [1-1:0] node1150;
	wire [1-1:0] node1151;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1161;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1170;
	wire [1-1:0] node1172;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1178;
	wire [1-1:0] node1179;
	wire [1-1:0] node1180;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1187;
	wire [1-1:0] node1188;
	wire [1-1:0] node1192;
	wire [1-1:0] node1193;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1200;
	wire [1-1:0] node1201;
	wire [1-1:0] node1203;
	wire [1-1:0] node1206;
	wire [1-1:0] node1207;
	wire [1-1:0] node1209;
	wire [1-1:0] node1212;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1219;
	wire [1-1:0] node1222;
	wire [1-1:0] node1223;
	wire [1-1:0] node1225;
	wire [1-1:0] node1228;
	wire [1-1:0] node1230;
	wire [1-1:0] node1233;
	wire [1-1:0] node1234;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1238;
	wire [1-1:0] node1240;
	wire [1-1:0] node1243;
	wire [1-1:0] node1246;
	wire [1-1:0] node1247;
	wire [1-1:0] node1252;
	wire [1-1:0] node1253;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1260;
	wire [1-1:0] node1263;
	wire [1-1:0] node1265;
	wire [1-1:0] node1266;
	wire [1-1:0] node1270;
	wire [1-1:0] node1271;
	wire [1-1:0] node1272;
	wire [1-1:0] node1274;
	wire [1-1:0] node1280;
	wire [1-1:0] node1281;
	wire [1-1:0] node1282;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1289;
	wire [1-1:0] node1291;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1303;
	wire [1-1:0] node1304;
	wire [1-1:0] node1308;
	wire [1-1:0] node1309;
	wire [1-1:0] node1311;
	wire [1-1:0] node1312;
	wire [1-1:0] node1314;
	wire [1-1:0] node1315;
	wire [1-1:0] node1321;
	wire [1-1:0] node1322;
	wire [1-1:0] node1323;
	wire [1-1:0] node1324;
	wire [1-1:0] node1325;
	wire [1-1:0] node1327;
	wire [1-1:0] node1328;
	wire [1-1:0] node1329;
	wire [1-1:0] node1331;
	wire [1-1:0] node1334;
	wire [1-1:0] node1336;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1347;
	wire [1-1:0] node1348;
	wire [1-1:0] node1350;
	wire [1-1:0] node1353;
	wire [1-1:0] node1354;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1363;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1368;
	wire [1-1:0] node1372;
	wire [1-1:0] node1374;
	wire [1-1:0] node1377;
	wire [1-1:0] node1379;
	wire [1-1:0] node1382;
	wire [1-1:0] node1383;
	wire [1-1:0] node1385;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1388;
	wire [1-1:0] node1392;
	wire [1-1:0] node1393;
	wire [1-1:0] node1397;
	wire [1-1:0] node1399;
	wire [1-1:0] node1403;
	wire [1-1:0] node1404;
	wire [1-1:0] node1405;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1411;
	wire [1-1:0] node1414;
	wire [1-1:0] node1415;
	wire [1-1:0] node1417;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1430;
	wire [1-1:0] node1432;
	wire [1-1:0] node1435;
	wire [1-1:0] node1436;
	wire [1-1:0] node1440;
	wire [1-1:0] node1442;
	wire [1-1:0] node1445;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1450;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1457;
	wire [1-1:0] node1460;
	wire [1-1:0] node1462;
	wire [1-1:0] node1463;
	wire [1-1:0] node1464;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1470;
	wire [1-1:0] node1471;
	wire [1-1:0] node1475;
	wire [1-1:0] node1477;
	wire [1-1:0] node1481;
	wire [1-1:0] node1482;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1486;
	wire [1-1:0] node1488;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1494;
	wire [1-1:0] node1497;
	wire [1-1:0] node1499;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1505;
	wire [1-1:0] node1506;
	wire [1-1:0] node1507;
	wire [1-1:0] node1509;
	wire [1-1:0] node1512;
	wire [1-1:0] node1514;
	wire [1-1:0] node1517;
	wire [1-1:0] node1518;
	wire [1-1:0] node1522;
	wire [1-1:0] node1524;
	wire [1-1:0] node1525;
	wire [1-1:0] node1527;
	wire [1-1:0] node1530;
	wire [1-1:0] node1532;
	wire [1-1:0] node1533;
	wire [1-1:0] node1537;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1541;
	wire [1-1:0] node1542;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1558;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1562;
	wire [1-1:0] node1563;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1569;
	wire [1-1:0] node1570;
	wire [1-1:0] node1574;
	wire [1-1:0] node1576;
	wire [1-1:0] node1580;
	wire [1-1:0] node1581;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1586;
	wire [1-1:0] node1589;
	wire [1-1:0] node1590;
	wire [1-1:0] node1591;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1603;
	wire [1-1:0] node1605;
	wire [1-1:0] node1608;
	wire [1-1:0] node1610;
	wire [1-1:0] node1613;
	wire [1-1:0] node1614;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1621;
	wire [1-1:0] node1622;
	wire [1-1:0] node1623;
	wire [1-1:0] node1624;
	wire [1-1:0] node1628;
	wire [1-1:0] node1629;
	wire [1-1:0] node1633;
	wire [1-1:0] node1635;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1641;
	wire [1-1:0] node1642;
	wire [1-1:0] node1643;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1653;
	wire [1-1:0] node1654;
	wire [1-1:0] node1658;
	wire [1-1:0] node1660;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1667;
	wire [1-1:0] node1668;
	wire [1-1:0] node1670;
	wire [1-1:0] node1673;
	wire [1-1:0] node1675;
	wire [1-1:0] node1678;
	wire [1-1:0] node1679;
	wire [1-1:0] node1683;
	wire [1-1:0] node1685;
	wire [1-1:0] node1686;
	wire [1-1:0] node1687;
	wire [1-1:0] node1691;
	wire [1-1:0] node1692;
	wire [1-1:0] node1694;
	wire [1-1:0] node1697;
	wire [1-1:0] node1699;
	wire [1-1:0] node1702;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1706;
	wire [1-1:0] node1708;
	wire [1-1:0] node1711;
	wire [1-1:0] node1712;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1725;
	wire [1-1:0] node1726;
	wire [1-1:0] node1728;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1731;
	wire [1-1:0] node1735;
	wire [1-1:0] node1737;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1746;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1756;
	wire [1-1:0] node1757;
	wire [1-1:0] node1761;
	wire [1-1:0] node1762;
	wire [1-1:0] node1763;
	wire [1-1:0] node1764;
	wire [1-1:0] node1768;
	wire [1-1:0] node1769;
	wire [1-1:0] node1773;
	wire [1-1:0] node1775;
	wire [1-1:0] node1776;
	wire [1-1:0] node1777;
	wire [1-1:0] node1781;
	wire [1-1:0] node1784;
	wire [1-1:0] node1785;
	wire [1-1:0] node1787;
	wire [1-1:0] node1788;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1794;
	wire [1-1:0] node1795;
	wire [1-1:0] node1799;
	wire [1-1:0] node1800;
	wire [1-1:0] node1805;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1809;
	wire [1-1:0] node1810;
	wire [1-1:0] node1811;
	wire [1-1:0] node1815;
	wire [1-1:0] node1816;
	wire [1-1:0] node1818;
	wire [1-1:0] node1821;
	wire [1-1:0] node1823;
	wire [1-1:0] node1827;
	wire [1-1:0] node1828;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1831;
	wire [1-1:0] node1832;
	wire [1-1:0] node1834;
	wire [1-1:0] node1837;
	wire [1-1:0] node1839;
	wire [1-1:0] node1842;
	wire [1-1:0] node1843;
	wire [1-1:0] node1848;
	wire [1-1:0] node1849;
	wire [1-1:0] node1851;
	wire [1-1:0] node1854;
	wire [1-1:0] node1855;
	wire [1-1:0] node1856;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1865;
	wire [1-1:0] node1867;
	wire [1-1:0] node1868;
	wire [1-1:0] node1869;
	wire [1-1:0] node1870;
	wire [1-1:0] node1873;
	wire [1-1:0] node1875;
	wire [1-1:0] node1878;
	wire [1-1:0] node1880;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1886;
	wire [1-1:0] node1887;
	wire [1-1:0] node1888;
	wire [1-1:0] node1889;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1893;
	wire [1-1:0] node1894;
	wire [1-1:0] node1898;
	wire [1-1:0] node1901;
	wire [1-1:0] node1903;
	wire [1-1:0] node1907;
	wire [1-1:0] node1908;
	wire [1-1:0] node1909;
	wire [1-1:0] node1910;
	wire [1-1:0] node1912;
	wire [1-1:0] node1914;
	wire [1-1:0] node1917;
	wire [1-1:0] node1918;
	wire [1-1:0] node1923;
	wire [1-1:0] node1924;
	wire [1-1:0] node1926;
	wire [1-1:0] node1929;
	wire [1-1:0] node1930;
	wire [1-1:0] node1931;
	wire [1-1:0] node1935;
	wire [1-1:0] node1936;
	wire [1-1:0] node1940;
	wire [1-1:0] node1941;
	wire [1-1:0] node1943;
	wire [1-1:0] node1944;
	wire [1-1:0] node1945;
	wire [1-1:0] node1946;
	wire [1-1:0] node1950;
	wire [1-1:0] node1951;
	wire [1-1:0] node1955;
	wire [1-1:0] node1957;
	wire [1-1:0] node1961;
	wire [1-1:0] node1962;
	wire [1-1:0] node1963;
	wire [1-1:0] node1965;
	wire [1-1:0] node1966;
	wire [1-1:0] node1967;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1974;
	wire [1-1:0] node1976;
	wire [1-1:0] node1979;
	wire [1-1:0] node1980;
	wire [1-1:0] node1985;
	wire [1-1:0] node1986;
	wire [1-1:0] node1987;
	wire [1-1:0] node1988;
	wire [1-1:0] node1989;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1997;
	wire [1-1:0] node1998;
	wire [1-1:0] node2002;
	wire [1-1:0] node2004;
	wire [1-1:0] node2005;
	wire [1-1:0] node2007;
	wire [1-1:0] node2010;
	wire [1-1:0] node2011;
	wire [1-1:0] node2013;
	wire [1-1:0] node2016;
	wire [1-1:0] node2017;
	wire [1-1:0] node2021;
	wire [1-1:0] node2023;
	wire [1-1:0] node2024;
	wire [1-1:0] node2025;
	wire [1-1:0] node2027;
	wire [1-1:0] node2030;
	wire [1-1:0] node2031;
	wire [1-1:0] node2033;
	wire [1-1:0] node2036;
	wire [1-1:0] node2038;
	wire [1-1:0] node2042;
	wire [1-1:0] node2043;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2047;
	wire [1-1:0] node2048;
	wire [1-1:0] node2050;
	wire [1-1:0] node2053;
	wire [1-1:0] node2055;
	wire [1-1:0] node2058;
	wire [1-1:0] node2059;
	wire [1-1:0] node2064;
	wire [1-1:0] node2065;
	wire [1-1:0] node2066;
	wire [1-1:0] node2067;
	wire [1-1:0] node2068;
	wire [1-1:0] node2069;
	wire [1-1:0] node2073;
	wire [1-1:0] node2074;
	wire [1-1:0] node2078;
	wire [1-1:0] node2080;
	wire [1-1:0] node2083;
	wire [1-1:0] node2085;
	wire [1-1:0] node2086;
	wire [1-1:0] node2087;
	wire [1-1:0] node2091;
	wire [1-1:0] node2092;
	wire [1-1:0] node2094;
	wire [1-1:0] node2097;
	wire [1-1:0] node2099;
	wire [1-1:0] node2102;
	wire [1-1:0] node2104;
	wire [1-1:0] node2105;
	wire [1-1:0] node2106;
	wire [1-1:0] node2108;
	wire [1-1:0] node2111;
	wire [1-1:0] node2112;
	wire [1-1:0] node2114;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2123;
	wire [1-1:0] node2124;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2128;
	wire [1-1:0] node2129;
	wire [1-1:0] node2130;
	wire [1-1:0] node2132;
	wire [1-1:0] node2135;
	wire [1-1:0] node2137;
	wire [1-1:0] node2140;
	wire [1-1:0] node2141;
	wire [1-1:0] node2146;
	wire [1-1:0] node2147;
	wire [1-1:0] node2148;
	wire [1-1:0] node2149;
	wire [1-1:0] node2151;
	wire [1-1:0] node2154;
	wire [1-1:0] node2155;
	wire [1-1:0] node2156;
	wire [1-1:0] node2160;
	wire [1-1:0] node2161;
	wire [1-1:0] node2165;
	wire [1-1:0] node2167;
	wire [1-1:0] node2168;
	wire [1-1:0] node2169;
	wire [1-1:0] node2170;
	wire [1-1:0] node2174;
	wire [1-1:0] node2175;
	wire [1-1:0] node2179;
	wire [1-1:0] node2180;
	wire [1-1:0] node2184;
	wire [1-1:0] node2186;
	wire [1-1:0] node2187;
	wire [1-1:0] node2188;
	wire [1-1:0] node2189;
	wire [1-1:0] node2191;
	wire [1-1:0] node2194;
	wire [1-1:0] node2195;
	wire [1-1:0] node2199;
	wire [1-1:0] node2201;
	wire [1-1:0] node2205;
	wire [1-1:0] node2206;
	wire [1-1:0] node2207;
	wire [1-1:0] node2208;
	wire [1-1:0] node2210;
	wire [1-1:0] node2211;
	wire [1-1:0] node2212;
	wire [1-1:0] node2213;
	wire [1-1:0] node2215;
	wire [1-1:0] node2218;
	wire [1-1:0] node2220;
	wire [1-1:0] node2223;
	wire [1-1:0] node2225;
	wire [1-1:0] node2229;
	wire [1-1:0] node2230;
	wire [1-1:0] node2231;
	wire [1-1:0] node2232;
	wire [1-1:0] node2233;
	wire [1-1:0] node2237;
	wire [1-1:0] node2238;
	wire [1-1:0] node2239;
	wire [1-1:0] node2243;
	wire [1-1:0] node2244;
	wire [1-1:0] node2249;
	wire [1-1:0] node2250;
	wire [1-1:0] node2251;
	wire [1-1:0] node2253;
	wire [1-1:0] node2256;
	wire [1-1:0] node2258;
	wire [1-1:0] node2261;
	wire [1-1:0] node2262;
	wire [1-1:0] node2266;
	wire [1-1:0] node2267;
	wire [1-1:0] node2269;
	wire [1-1:0] node2270;
	wire [1-1:0] node2271;
	wire [1-1:0] node2272;
	wire [1-1:0] node2276;
	wire [1-1:0] node2278;
	wire [1-1:0] node2281;
	wire [1-1:0] node2282;
	wire [1-1:0] node2287;
	wire [1-1:0] node2288;
	wire [1-1:0] node2289;
	wire [1-1:0] node2290;
	wire [1-1:0] node2292;
	wire [1-1:0] node2293;
	wire [1-1:0] node2295;
	wire [1-1:0] node2298;
	wire [1-1:0] node2299;
	wire [1-1:0] node2301;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2310;
	wire [1-1:0] node2311;
	wire [1-1:0] node2312;
	wire [1-1:0] node2313;
	wire [1-1:0] node2314;
	wire [1-1:0] node2318;
	wire [1-1:0] node2319;
	wire [1-1:0] node2320;
	wire [1-1:0] node2321;
	wire [1-1:0] node2324;
	wire [1-1:0] node2327;
	wire [1-1:0] node2329;
	wire [1-1:0] node2332;
	wire [1-1:0] node2336;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2339;
	wire [1-1:0] node2343;
	wire [1-1:0] node2344;
	wire [1-1:0] node2348;
	wire [1-1:0] node2349;
	wire [1-1:0] node2353;
	wire [1-1:0] node2354;
	wire [1-1:0] node2356;
	wire [1-1:0] node2357;
	wire [1-1:0] node2358;
	wire [1-1:0] node2359;
	wire [1-1:0] node2363;
	wire [1-1:0] node2365;
	wire [1-1:0] node2368;
	wire [1-1:0] node2370;
	wire [1-1:0] node2374;
	wire [1-1:0] node2375;
	wire [1-1:0] node2376;
	wire [1-1:0] node2377;
	wire [1-1:0] node2379;
	wire [1-1:0] node2380;
	wire [1-1:0] node2381;
	wire [1-1:0] node2385;
	wire [1-1:0] node2386;
	wire [1-1:0] node2387;
	wire [1-1:0] node2391;
	wire [1-1:0] node2393;
	wire [1-1:0] node2397;
	wire [1-1:0] node2398;
	wire [1-1:0] node2399;
	wire [1-1:0] node2400;
	wire [1-1:0] node2401;
	wire [1-1:0] node2402;
	wire [1-1:0] node2406;
	wire [1-1:0] node2408;
	wire [1-1:0] node2411;
	wire [1-1:0] node2413;
	wire [1-1:0] node2416;
	wire [1-1:0] node2418;
	wire [1-1:0] node2419;
	wire [1-1:0] node2420;
	wire [1-1:0] node2424;
	wire [1-1:0] node2425;
	wire [1-1:0] node2427;
	wire [1-1:0] node2430;
	wire [1-1:0] node2431;
	wire [1-1:0] node2435;
	wire [1-1:0] node2437;
	wire [1-1:0] node2438;
	wire [1-1:0] node2439;
	wire [1-1:0] node2440;
	wire [1-1:0] node2441;
	wire [1-1:0] node2445;
	wire [1-1:0] node2447;
	wire [1-1:0] node2450;
	wire [1-1:0] node2452;
	wire [1-1:0] node2456;
	wire [1-1:0] node2457;
	wire [1-1:0] node2458;
	wire [1-1:0] node2459;
	wire [1-1:0] node2460;
	wire [1-1:0] node2461;
	wire [1-1:0] node2463;
	wire [1-1:0] node2464;
	wire [1-1:0] node2465;
	wire [1-1:0] node2467;
	wire [1-1:0] node2470;
	wire [1-1:0] node2471;
	wire [1-1:0] node2473;
	wire [1-1:0] node2476;
	wire [1-1:0] node2477;
	wire [1-1:0] node2482;
	wire [1-1:0] node2483;
	wire [1-1:0] node2484;
	wire [1-1:0] node2485;
	wire [1-1:0] node2486;
	wire [1-1:0] node2487;
	wire [1-1:0] node2488;
	wire [1-1:0] node2490;
	wire [1-1:0] node2494;
	wire [1-1:0] node2495;
	wire [1-1:0] node2499;
	wire [1-1:0] node2501;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;
	wire [1-1:0] node2507;
	wire [1-1:0] node2509;
	wire [1-1:0] node2512;
	wire [1-1:0] node2514;
	wire [1-1:0] node2517;
	wire [1-1:0] node2519;
	wire [1-1:0] node2522;
	wire [1-1:0] node2523;
	wire [1-1:0] node2525;
	wire [1-1:0] node2526;
	wire [1-1:0] node2528;
	wire [1-1:0] node2531;
	wire [1-1:0] node2532;
	wire [1-1:0] node2533;
	wire [1-1:0] node2537;
	wire [1-1:0] node2539;
	wire [1-1:0] node2543;
	wire [1-1:0] node2544;
	wire [1-1:0] node2546;
	wire [1-1:0] node2547;
	wire [1-1:0] node2548;
	wire [1-1:0] node2549;
	wire [1-1:0] node2551;
	wire [1-1:0] node2554;
	wire [1-1:0] node2555;
	wire [1-1:0] node2559;
	wire [1-1:0] node2560;
	wire [1-1:0] node2565;
	wire [1-1:0] node2566;
	wire [1-1:0] node2567;
	wire [1-1:0] node2568;
	wire [1-1:0] node2569;
	wire [1-1:0] node2570;
	wire [1-1:0] node2574;
	wire [1-1:0] node2575;
	wire [1-1:0] node2576;
	wire [1-1:0] node2580;
	wire [1-1:0] node2581;
	wire [1-1:0] node2586;
	wire [1-1:0] node2587;
	wire [1-1:0] node2589;
	wire [1-1:0] node2592;
	wire [1-1:0] node2593;
	wire [1-1:0] node2595;
	wire [1-1:0] node2598;
	wire [1-1:0] node2600;
	wire [1-1:0] node2603;
	wire [1-1:0] node2604;
	wire [1-1:0] node2606;
	wire [1-1:0] node2607;
	wire [1-1:0] node2608;
	wire [1-1:0] node2610;
	wire [1-1:0] node2613;
	wire [1-1:0] node2615;
	wire [1-1:0] node2618;
	wire [1-1:0] node2620;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2626;
	wire [1-1:0] node2627;
	wire [1-1:0] node2629;
	wire [1-1:0] node2630;
	wire [1-1:0] node2631;
	wire [1-1:0] node2632;
	wire [1-1:0] node2636;
	wire [1-1:0] node2638;
	wire [1-1:0] node2641;
	wire [1-1:0] node2642;
	wire [1-1:0] node2647;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2654;
	wire [1-1:0] node2655;
	wire [1-1:0] node2656;
	wire [1-1:0] node2660;
	wire [1-1:0] node2661;
	wire [1-1:0] node2665;
	wire [1-1:0] node2667;
	wire [1-1:0] node2668;
	wire [1-1:0] node2669;
	wire [1-1:0] node2670;
	wire [1-1:0] node2674;
	wire [1-1:0] node2676;
	wire [1-1:0] node2679;
	wire [1-1:0] node2681;
	wire [1-1:0] node2684;
	wire [1-1:0] node2685;
	wire [1-1:0] node2687;
	wire [1-1:0] node2688;
	wire [1-1:0] node2689;
	wire [1-1:0] node2693;
	wire [1-1:0] node2694;
	wire [1-1:0] node2695;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2705;
	wire [1-1:0] node2706;
	wire [1-1:0] node2707;
	wire [1-1:0] node2708;
	wire [1-1:0] node2709;
	wire [1-1:0] node2711;
	wire [1-1:0] node2712;
	wire [1-1:0] node2713;
	wire [1-1:0] node2714;
	wire [1-1:0] node2715;
	wire [1-1:0] node2716;
	wire [1-1:0] node2719;
	wire [1-1:0] node2723;
	wire [1-1:0] node2724;
	wire [1-1:0] node2727;
	wire [1-1:0] node2729;
	wire [1-1:0] node2732;
	wire [1-1:0] node2734;
	wire [1-1:0] node2738;
	wire [1-1:0] node2739;
	wire [1-1:0] node2740;
	wire [1-1:0] node2741;
	wire [1-1:0] node2742;
	wire [1-1:0] node2743;
	wire [1-1:0] node2747;
	wire [1-1:0] node2748;
	wire [1-1:0] node2752;
	wire [1-1:0] node2754;
	wire [1-1:0] node2758;
	wire [1-1:0] node2759;
	wire [1-1:0] node2760;
	wire [1-1:0] node2762;
	wire [1-1:0] node2765;
	wire [1-1:0] node2766;
	wire [1-1:0] node2770;
	wire [1-1:0] node2772;
	wire [1-1:0] node2775;
	wire [1-1:0] node2777;
	wire [1-1:0] node2778;
	wire [1-1:0] node2779;
	wire [1-1:0] node2780;
	wire [1-1:0] node2781;
	wire [1-1:0] node2785;
	wire [1-1:0] node2787;
	wire [1-1:0] node2790;
	wire [1-1:0] node2791;
	wire [1-1:0] node2796;
	wire [1-1:0] node2797;
	wire [1-1:0] node2798;
	wire [1-1:0] node2799;
	wire [1-1:0] node2801;
	wire [1-1:0] node2802;
	wire [1-1:0] node2803;
	wire [1-1:0] node2804;
	wire [1-1:0] node2805;
	wire [1-1:0] node2810;
	wire [1-1:0] node2811;
	wire [1-1:0] node2816;
	wire [1-1:0] node2817;
	wire [1-1:0] node2818;
	wire [1-1:0] node2819;
	wire [1-1:0] node2821;
	wire [1-1:0] node2824;
	wire [1-1:0] node2825;
	wire [1-1:0] node2829;
	wire [1-1:0] node2831;
	wire [1-1:0] node2834;
	wire [1-1:0] node2836;
	wire [1-1:0] node2837;
	wire [1-1:0] node2838;
	wire [1-1:0] node2842;
	wire [1-1:0] node2843;
	wire [1-1:0] node2845;
	wire [1-1:0] node2848;
	wire [1-1:0] node2850;
	wire [1-1:0] node2853;
	wire [1-1:0] node2855;
	wire [1-1:0] node2856;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2859;
	wire [1-1:0] node2863;
	wire [1-1:0] node2865;
	wire [1-1:0] node2868;
	wire [1-1:0] node2870;
	wire [1-1:0] node2874;
	wire [1-1:0] node2875;
	wire [1-1:0] node2877;
	wire [1-1:0] node2878;
	wire [1-1:0] node2879;
	wire [1-1:0] node2880;
	wire [1-1:0] node2881;
	wire [1-1:0] node2885;
	wire [1-1:0] node2886;
	wire [1-1:0] node2890;
	wire [1-1:0] node2892;
	wire [1-1:0] node2896;
	wire [1-1:0] node2897;
	wire [1-1:0] node2898;
	wire [1-1:0] node2899;
	wire [1-1:0] node2900;
	wire [1-1:0] node2901;
	wire [1-1:0] node2905;
	wire [1-1:0] node2906;
	wire [1-1:0] node2908;
	wire [1-1:0] node2911;
	wire [1-1:0] node2912;
	wire [1-1:0] node2917;
	wire [1-1:0] node2918;
	wire [1-1:0] node2919;
	wire [1-1:0] node2921;
	wire [1-1:0] node2924;
	wire [1-1:0] node2925;
	wire [1-1:0] node2929;
	wire [1-1:0] node2930;
	wire [1-1:0] node2934;
	wire [1-1:0] node2935;
	wire [1-1:0] node2937;
	wire [1-1:0] node2938;
	wire [1-1:0] node2939;
	wire [1-1:0] node2941;
	wire [1-1:0] node2944;
	wire [1-1:0] node2945;
	wire [1-1:0] node2949;
	wire [1-1:0] node2951;
	wire [1-1:0] node2955;
	wire [1-1:0] node2956;
	wire [1-1:0] node2957;
	wire [1-1:0] node2958;
	wire [1-1:0] node2960;
	wire [1-1:0] node2961;
	wire [1-1:0] node2962;
	wire [1-1:0] node2963;
	wire [1-1:0] node2967;
	wire [1-1:0] node2968;
	wire [1-1:0] node2969;
	wire [1-1:0] node2973;
	wire [1-1:0] node2975;
	wire [1-1:0] node2979;
	wire [1-1:0] node2980;
	wire [1-1:0] node2981;
	wire [1-1:0] node2982;
	wire [1-1:0] node2983;
	wire [1-1:0] node2984;
	wire [1-1:0] node2986;
	wire [1-1:0] node2989;
	wire [1-1:0] node2991;
	wire [1-1:0] node2994;
	wire [1-1:0] node2995;
	wire [1-1:0] node3000;
	wire [1-1:0] node3001;
	wire [1-1:0] node3002;
	wire [1-1:0] node3004;
	wire [1-1:0] node3007;
	wire [1-1:0] node3009;
	wire [1-1:0] node3012;
	wire [1-1:0] node3013;
	wire [1-1:0] node3017;
	wire [1-1:0] node3018;
	wire [1-1:0] node3020;
	wire [1-1:0] node3021;
	wire [1-1:0] node3022;
	wire [1-1:0] node3026;
	wire [1-1:0] node3027;
	wire [1-1:0] node3028;
	wire [1-1:0] node3032;
	wire [1-1:0] node3033;
	wire [1-1:0] node3038;
	wire [1-1:0] node3039;
	wire [1-1:0] node3040;
	wire [1-1:0] node3042;
	wire [1-1:0] node3043;
	wire [1-1:0] node3044;
	wire [1-1:0] node3046;
	wire [1-1:0] node3049;
	wire [1-1:0] node3050;
	wire [1-1:0] node3052;
	wire [1-1:0] node3055;
	wire [1-1:0] node3057;
	wire [1-1:0] node3061;
	wire [1-1:0] node3062;
	wire [1-1:0] node3063;
	wire [1-1:0] node3064;
	wire [1-1:0] node3065;
	wire [1-1:0] node3066;
	wire [1-1:0] node3070;
	wire [1-1:0] node3071;
	wire [1-1:0] node3075;
	wire [1-1:0] node3077;
	wire [1-1:0] node3081;
	wire [1-1:0] node3082;
	wire [1-1:0] node3083;
	wire [1-1:0] node3087;
	wire [1-1:0] node3088;
	wire [1-1:0] node3090;
	wire [1-1:0] node3093;
	wire [1-1:0] node3095;
	wire [1-1:0] node3098;
	wire [1-1:0] node3099;
	wire [1-1:0] node3101;
	wire [1-1:0] node3102;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3108;
	wire [1-1:0] node3109;
	wire [1-1:0] node3111;
	wire [1-1:0] node3115;
	wire [1-1:0] node3117;
	wire [1-1:0] node3121;
	wire [1-1:0] node3122;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3126;
	wire [1-1:0] node3127;
	wire [1-1:0] node3128;
	wire [1-1:0] node3129;
	wire [1-1:0] node3133;
	wire [1-1:0] node3134;
	wire [1-1:0] node3138;
	wire [1-1:0] node3139;
	wire [1-1:0] node3144;
	wire [1-1:0] node3145;
	wire [1-1:0] node3146;
	wire [1-1:0] node3147;
	wire [1-1:0] node3149;
	wire [1-1:0] node3152;
	wire [1-1:0] node3153;
	wire [1-1:0] node3155;
	wire [1-1:0] node3158;
	wire [1-1:0] node3162;
	wire [1-1:0] node3163;
	wire [1-1:0] node3164;
	wire [1-1:0] node3165;
	wire [1-1:0] node3169;
	wire [1-1:0] node3170;
	wire [1-1:0] node3174;
	wire [1-1:0] node3176;
	wire [1-1:0] node3179;
	wire [1-1:0] node3180;
	wire [1-1:0] node3182;
	wire [1-1:0] node3183;
	wire [1-1:0] node3184;
	wire [1-1:0] node3188;
	wire [1-1:0] node3189;
	wire [1-1:0] node3191;
	wire [1-1:0] node3194;
	wire [1-1:0] node3195;
	wire [1-1:0] node3200;
	wire [1-1:0] node3201;
	wire [1-1:0] node3202;
	wire [1-1:0] node3204;
	wire [1-1:0] node3205;
	wire [1-1:0] node3206;
	wire [1-1:0] node3208;
	wire [1-1:0] node3211;
	wire [1-1:0] node3212;
	wire [1-1:0] node3214;
	wire [1-1:0] node3217;
	wire [1-1:0] node3219;
	wire [1-1:0] node3223;
	wire [1-1:0] node3224;
	wire [1-1:0] node3225;
	wire [1-1:0] node3226;
	wire [1-1:0] node3227;
	wire [1-1:0] node3231;
	wire [1-1:0] node3232;
	wire [1-1:0] node3233;
	wire [1-1:0] node3237;
	wire [1-1:0] node3239;
	wire [1-1:0] node3243;
	wire [1-1:0] node3244;
	wire [1-1:0] node3245;
	wire [1-1:0] node3246;
	wire [1-1:0] node3250;
	wire [1-1:0] node3251;
	wire [1-1:0] node3255;
	wire [1-1:0] node3256;
	wire [1-1:0] node3260;
	wire [1-1:0] node3262;
	wire [1-1:0] node3263;
	wire [1-1:0] node3264;
	wire [1-1:0] node3265;
	wire [1-1:0] node3266;
	wire [1-1:0] node3270;
	wire [1-1:0] node3271;
	wire [1-1:0] node3275;
	wire [1-1:0] node3277;

	assign outp = (inp[5]) ? node2374 : node1;
		assign node1 = (inp[6]) ? node857 : node2;
			assign node2 = (inp[12]) ? node84 : node3;
				assign node3 = (inp[0]) ? node25 : node4;
					assign node4 = (inp[1]) ? node6 : 1'b1;
						assign node6 = (inp[8]) ? 1'b1 : node7;
							assign node7 = (inp[14]) ? node13 : node8;
								assign node8 = (inp[13]) ? node10 : 1'b0;
									assign node10 = (inp[11]) ? 1'b0 : 1'b1;
								assign node13 = (inp[2]) ? node19 : node14;
									assign node14 = (inp[11]) ? 1'b1 : node15;
										assign node15 = (inp[13]) ? 1'b0 : 1'b1;
									assign node19 = (inp[11]) ? 1'b0 : node20;
										assign node20 = (inp[13]) ? 1'b1 : 1'b0;
					assign node25 = (inp[4]) ? node63 : node26;
						assign node26 = (inp[1]) ? node44 : node27;
							assign node27 = (inp[14]) ? node33 : node28;
								assign node28 = (inp[11]) ? 1'b0 : node29;
									assign node29 = (inp[13]) ? 1'b1 : 1'b0;
								assign node33 = (inp[2]) ? node39 : node34;
									assign node34 = (inp[11]) ? 1'b1 : node35;
										assign node35 = (inp[13]) ? 1'b0 : 1'b1;
									assign node39 = (inp[11]) ? 1'b0 : node40;
										assign node40 = (inp[13]) ? 1'b1 : 1'b0;
							assign node44 = (inp[8]) ? node46 : 1'b1;
								assign node46 = (inp[11]) ? node58 : node47;
									assign node47 = (inp[13]) ? node53 : node48;
										assign node48 = (inp[14]) ? node50 : 1'b0;
											assign node50 = (inp[2]) ? 1'b0 : 1'b1;
										assign node53 = (inp[14]) ? node55 : 1'b1;
											assign node55 = (inp[2]) ? 1'b1 : 1'b0;
									assign node58 = (inp[2]) ? 1'b0 : node59;
										assign node59 = (inp[14]) ? 1'b1 : 1'b0;
						assign node63 = (inp[1]) ? node65 : 1'b1;
							assign node65 = (inp[8]) ? 1'b1 : node66;
								assign node66 = (inp[13]) ? node72 : node67;
									assign node67 = (inp[14]) ? node69 : 1'b0;
										assign node69 = (inp[2]) ? 1'b0 : 1'b1;
									assign node72 = (inp[11]) ? node78 : node73;
										assign node73 = (inp[2]) ? 1'b1 : node74;
											assign node74 = (inp[14]) ? 1'b0 : 1'b1;
										assign node78 = (inp[2]) ? 1'b0 : node79;
											assign node79 = (inp[14]) ? 1'b1 : 1'b0;
				assign node84 = (inp[15]) ? node776 : node85;
					assign node85 = (inp[10]) ? node539 : node86;
						assign node86 = (inp[9]) ? node298 : node87;
							assign node87 = (inp[7]) ? node217 : node88;
								assign node88 = (inp[3]) ? node162 : node89;
									assign node89 = (inp[1]) ? node111 : node90;
										assign node90 = (inp[4]) ? 1'b0 : node91;
											assign node91 = (inp[0]) ? node93 : 1'b0;
												assign node93 = (inp[14]) ? node99 : node94;
													assign node94 = (inp[11]) ? 1'b1 : node95;
														assign node95 = (inp[13]) ? 1'b0 : 1'b1;
													assign node99 = (inp[13]) ? node101 : 1'b0;
														assign node101 = (inp[8]) ? node103 : 1'b1;
															assign node103 = (inp[11]) ? node107 : node104;
																assign node104 = (inp[2]) ? 1'b0 : 1'b1;
																assign node107 = (inp[2]) ? 1'b1 : 1'b0;
										assign node111 = (inp[8]) ? node145 : node112;
											assign node112 = (inp[4]) ? node128 : node113;
												assign node113 = (inp[0]) ? 1'b0 : node114;
													assign node114 = (inp[11]) ? node122 : node115;
														assign node115 = (inp[2]) ? 1'b0 : node116;
															assign node116 = (inp[13]) ? 1'b1 : node117;
																assign node117 = (inp[14]) ? 1'b0 : 1'b1;
														assign node122 = (inp[14]) ? node124 : 1'b1;
															assign node124 = (inp[13]) ? 1'b1 : 1'b0;
												assign node128 = (inp[13]) ? node134 : node129;
													assign node129 = (inp[14]) ? node131 : 1'b1;
														assign node131 = (inp[2]) ? 1'b1 : 1'b0;
													assign node134 = (inp[11]) ? node140 : node135;
														assign node135 = (inp[2]) ? 1'b0 : node136;
															assign node136 = (inp[14]) ? 1'b1 : 1'b0;
														assign node140 = (inp[2]) ? 1'b1 : node141;
															assign node141 = (inp[14]) ? 1'b0 : 1'b1;
											assign node145 = (inp[0]) ? node147 : 1'b0;
												assign node147 = (inp[4]) ? 1'b0 : node148;
													assign node148 = (inp[11]) ? node156 : node149;
														assign node149 = (inp[13]) ? 1'b0 : node150;
															assign node150 = (inp[14]) ? node152 : 1'b1;
																assign node152 = (inp[2]) ? 1'b1 : 1'b0;
														assign node156 = (inp[14]) ? node158 : 1'b1;
															assign node158 = (inp[2]) ? 1'b1 : 1'b0;
									assign node162 = (inp[0]) ? node182 : node163;
										assign node163 = (inp[1]) ? node165 : 1'b1;
											assign node165 = (inp[8]) ? 1'b1 : node166;
												assign node166 = (inp[11]) ? node176 : node167;
													assign node167 = (inp[13]) ? node171 : node168;
														assign node168 = (inp[14]) ? 1'b1 : 1'b0;
														assign node171 = (inp[14]) ? node173 : 1'b1;
															assign node173 = (inp[2]) ? 1'b1 : 1'b0;
													assign node176 = (inp[2]) ? 1'b0 : node177;
														assign node177 = (inp[14]) ? 1'b1 : 1'b0;
										assign node182 = (inp[4]) ? node206 : node183;
											assign node183 = (inp[1]) ? node197 : node184;
												assign node184 = (inp[14]) ? node190 : node185;
													assign node185 = (inp[13]) ? node187 : 1'b0;
														assign node187 = (inp[11]) ? 1'b0 : 1'b1;
													assign node190 = (inp[2]) ? node194 : node191;
														assign node191 = (inp[11]) ? 1'b1 : 1'b0;
														assign node194 = (inp[11]) ? 1'b0 : 1'b1;
												assign node197 = (inp[8]) ? node199 : 1'b1;
													assign node199 = (inp[11]) ? node201 : 1'b1;
														assign node201 = (inp[2]) ? 1'b0 : node202;
															assign node202 = (inp[14]) ? 1'b1 : 1'b0;
											assign node206 = (inp[8]) ? 1'b1 : node207;
												assign node207 = (inp[1]) ? node209 : 1'b1;
													assign node209 = (inp[14]) ? node211 : 1'b0;
														assign node211 = (inp[11]) ? 1'b0 : node212;
															assign node212 = (inp[2]) ? 1'b1 : 1'b0;
								assign node217 = (inp[8]) ? node277 : node218;
									assign node218 = (inp[1]) ? node236 : node219;
										assign node219 = (inp[0]) ? node221 : 1'b0;
											assign node221 = (inp[4]) ? 1'b0 : node222;
												assign node222 = (inp[11]) ? node230 : node223;
													assign node223 = (inp[13]) ? 1'b0 : node224;
														assign node224 = (inp[14]) ? node226 : 1'b1;
															assign node226 = (inp[3]) ? 1'b0 : 1'b1;
													assign node230 = (inp[14]) ? node232 : 1'b1;
														assign node232 = (inp[2]) ? 1'b1 : 1'b0;
										assign node236 = (inp[0]) ? node254 : node237;
											assign node237 = (inp[13]) ? node243 : node238;
												assign node238 = (inp[14]) ? node240 : 1'b1;
													assign node240 = (inp[2]) ? 1'b1 : 1'b0;
												assign node243 = (inp[11]) ? node249 : node244;
													assign node244 = (inp[2]) ? 1'b0 : node245;
														assign node245 = (inp[14]) ? 1'b1 : 1'b0;
													assign node249 = (inp[14]) ? node251 : 1'b1;
														assign node251 = (inp[2]) ? 1'b1 : 1'b0;
											assign node254 = (inp[4]) ? node256 : 1'b0;
												assign node256 = (inp[13]) ? node262 : node257;
													assign node257 = (inp[14]) ? node259 : 1'b1;
														assign node259 = (inp[2]) ? 1'b1 : 1'b0;
													assign node262 = (inp[14]) ? node264 : 1'b0;
														assign node264 = (inp[3]) ? node272 : node265;
															assign node265 = (inp[2]) ? node269 : node266;
																assign node266 = (inp[11]) ? 1'b0 : 1'b1;
																assign node269 = (inp[11]) ? 1'b1 : 1'b0;
															assign node272 = (inp[11]) ? 1'b1 : node273;
																assign node273 = (inp[2]) ? 1'b0 : 1'b1;
									assign node277 = (inp[0]) ? node279 : 1'b0;
										assign node279 = (inp[4]) ? 1'b0 : node280;
											assign node280 = (inp[14]) ? node286 : node281;
												assign node281 = (inp[13]) ? node283 : 1'b1;
													assign node283 = (inp[11]) ? 1'b1 : 1'b0;
												assign node286 = (inp[2]) ? node292 : node287;
													assign node287 = (inp[11]) ? 1'b0 : node288;
														assign node288 = (inp[13]) ? 1'b1 : 1'b0;
													assign node292 = (inp[13]) ? node294 : 1'b1;
														assign node294 = (inp[11]) ? 1'b1 : 1'b0;
							assign node298 = (inp[3]) ? node376 : node299;
								assign node299 = (inp[4]) ? node355 : node300;
									assign node300 = (inp[0]) ? node318 : node301;
										assign node301 = (inp[1]) ? node303 : 1'b1;
											assign node303 = (inp[8]) ? 1'b1 : node304;
												assign node304 = (inp[11]) ? node312 : node305;
													assign node305 = (inp[13]) ? 1'b1 : node306;
														assign node306 = (inp[14]) ? node308 : 1'b0;
															assign node308 = (inp[2]) ? 1'b0 : 1'b1;
													assign node312 = (inp[2]) ? 1'b0 : node313;
														assign node313 = (inp[14]) ? 1'b1 : 1'b0;
										assign node318 = (inp[8]) ? node338 : node319;
											assign node319 = (inp[1]) ? 1'b1 : node320;
												assign node320 = (inp[14]) ? node326 : node321;
													assign node321 = (inp[11]) ? 1'b0 : node322;
														assign node322 = (inp[13]) ? 1'b1 : 1'b0;
													assign node326 = (inp[2]) ? node332 : node327;
														assign node327 = (inp[11]) ? 1'b1 : node328;
															assign node328 = (inp[13]) ? 1'b0 : 1'b1;
														assign node332 = (inp[13]) ? node334 : 1'b0;
															assign node334 = (inp[11]) ? 1'b0 : 1'b1;
											assign node338 = (inp[2]) ? node350 : node339;
												assign node339 = (inp[14]) ? node345 : node340;
													assign node340 = (inp[13]) ? node342 : 1'b0;
														assign node342 = (inp[11]) ? 1'b0 : 1'b1;
													assign node345 = (inp[11]) ? 1'b1 : node346;
														assign node346 = (inp[13]) ? 1'b0 : 1'b1;
												assign node350 = (inp[11]) ? 1'b0 : node351;
													assign node351 = (inp[13]) ? 1'b1 : 1'b0;
									assign node355 = (inp[1]) ? node357 : 1'b1;
										assign node357 = (inp[8]) ? 1'b1 : node358;
											assign node358 = (inp[11]) ? node370 : node359;
												assign node359 = (inp[13]) ? node365 : node360;
													assign node360 = (inp[2]) ? 1'b0 : node361;
														assign node361 = (inp[14]) ? 1'b1 : 1'b0;
													assign node365 = (inp[2]) ? 1'b1 : node366;
														assign node366 = (inp[14]) ? 1'b0 : 1'b1;
												assign node370 = (inp[14]) ? node372 : 1'b0;
													assign node372 = (inp[2]) ? 1'b0 : 1'b1;
								assign node376 = (inp[7]) ? node468 : node377;
									assign node377 = (inp[8]) ? node447 : node378;
										assign node378 = (inp[13]) ? node412 : node379;
											assign node379 = (inp[14]) ? node403 : node380;
												assign node380 = (inp[11]) ? node386 : node381;
													assign node381 = (inp[1]) ? 1'b1 : node382;
														assign node382 = (inp[0]) ? 1'b1 : 1'b0;
													assign node386 = (inp[0]) ? node390 : node387;
														assign node387 = (inp[1]) ? 1'b1 : 1'b0;
														assign node390 = (inp[2]) ? node396 : node391;
															assign node391 = (inp[1]) ? 1'b0 : node392;
																assign node392 = (inp[4]) ? 1'b0 : 1'b1;
															assign node396 = (inp[4]) ? node400 : node397;
																assign node397 = (inp[1]) ? 1'b0 : 1'b1;
																assign node400 = (inp[1]) ? 1'b1 : 1'b0;
												assign node403 = (inp[2]) ? node405 : 1'b0;
													assign node405 = (inp[1]) ? 1'b1 : node406;
														assign node406 = (inp[0]) ? node408 : 1'b0;
															assign node408 = (inp[4]) ? 1'b0 : 1'b1;
											assign node412 = (inp[2]) ? node434 : node413;
												assign node413 = (inp[0]) ? node425 : node414;
													assign node414 = (inp[1]) ? node416 : 1'b0;
														assign node416 = (inp[4]) ? 1'b1 : node417;
															assign node417 = (inp[11]) ? node421 : node418;
																assign node418 = (inp[14]) ? 1'b1 : 1'b0;
																assign node421 = (inp[14]) ? 1'b0 : 1'b1;
													assign node425 = (inp[11]) ? node427 : 1'b0;
														assign node427 = (inp[14]) ? 1'b0 : node428;
															assign node428 = (inp[1]) ? node430 : 1'b1;
																assign node430 = (inp[4]) ? 1'b1 : 1'b0;
												assign node434 = (inp[11]) ? node436 : 1'b0;
													assign node436 = (inp[14]) ? node438 : 1'b0;
														assign node438 = (inp[0]) ? node440 : 1'b0;
															assign node440 = (inp[1]) ? node444 : node441;
																assign node441 = (inp[4]) ? 1'b0 : 1'b1;
																assign node444 = (inp[4]) ? 1'b1 : 1'b0;
										assign node447 = (inp[0]) ? node449 : 1'b0;
											assign node449 = (inp[4]) ? 1'b0 : node450;
												assign node450 = (inp[11]) ? node462 : node451;
													assign node451 = (inp[13]) ? node457 : node452;
														assign node452 = (inp[14]) ? node454 : 1'b1;
															assign node454 = (inp[2]) ? 1'b1 : 1'b0;
														assign node457 = (inp[2]) ? 1'b0 : node458;
															assign node458 = (inp[14]) ? 1'b1 : 1'b0;
													assign node462 = (inp[2]) ? 1'b1 : node463;
														assign node463 = (inp[14]) ? 1'b0 : 1'b1;
									assign node468 = (inp[0]) ? node490 : node469;
										assign node469 = (inp[8]) ? 1'b1 : node470;
											assign node470 = (inp[1]) ? node472 : 1'b1;
												assign node472 = (inp[11]) ? node484 : node473;
													assign node473 = (inp[13]) ? node479 : node474;
														assign node474 = (inp[14]) ? node476 : 1'b0;
															assign node476 = (inp[2]) ? 1'b0 : 1'b1;
														assign node479 = (inp[2]) ? 1'b1 : node480;
															assign node480 = (inp[14]) ? 1'b0 : 1'b1;
													assign node484 = (inp[2]) ? 1'b0 : node485;
														assign node485 = (inp[14]) ? 1'b1 : 1'b0;
										assign node490 = (inp[4]) ? node522 : node491;
											assign node491 = (inp[8]) ? node505 : node492;
												assign node492 = (inp[1]) ? 1'b1 : node493;
													assign node493 = (inp[13]) ? node499 : node494;
														assign node494 = (inp[2]) ? 1'b0 : node495;
															assign node495 = (inp[14]) ? 1'b1 : 1'b0;
														assign node499 = (inp[11]) ? node501 : 1'b1;
															assign node501 = (inp[2]) ? 1'b0 : 1'b1;
												assign node505 = (inp[14]) ? node511 : node506;
													assign node506 = (inp[11]) ? 1'b0 : node507;
														assign node507 = (inp[13]) ? 1'b1 : 1'b0;
													assign node511 = (inp[2]) ? node517 : node512;
														assign node512 = (inp[13]) ? node514 : 1'b1;
															assign node514 = (inp[11]) ? 1'b1 : 1'b0;
														assign node517 = (inp[13]) ? node519 : 1'b0;
															assign node519 = (inp[11]) ? 1'b0 : 1'b1;
											assign node522 = (inp[8]) ? 1'b1 : node523;
												assign node523 = (inp[1]) ? node525 : 1'b1;
													assign node525 = (inp[14]) ? node531 : node526;
														assign node526 = (inp[13]) ? node528 : 1'b0;
															assign node528 = (inp[11]) ? 1'b0 : 1'b1;
														assign node531 = (inp[2]) ? node533 : 1'b1;
															assign node533 = (inp[13]) ? node535 : 1'b0;
																assign node535 = (inp[11]) ? 1'b0 : 1'b1;
						assign node539 = (inp[7]) ? node695 : node540;
							assign node540 = (inp[3]) ? node618 : node541;
								assign node541 = (inp[8]) ? node597 : node542;
									assign node542 = (inp[1]) ? node562 : node543;
										assign node543 = (inp[0]) ? node545 : 1'b0;
											assign node545 = (inp[4]) ? 1'b0 : node546;
												assign node546 = (inp[13]) ? node552 : node547;
													assign node547 = (inp[2]) ? 1'b1 : node548;
														assign node548 = (inp[14]) ? 1'b0 : 1'b1;
													assign node552 = (inp[11]) ? node558 : node553;
														assign node553 = (inp[14]) ? node555 : 1'b0;
															assign node555 = (inp[2]) ? 1'b0 : 1'b1;
														assign node558 = (inp[2]) ? 1'b1 : 1'b0;
										assign node562 = (inp[0]) ? node580 : node563;
											assign node563 = (inp[11]) ? node575 : node564;
												assign node564 = (inp[13]) ? node570 : node565;
													assign node565 = (inp[14]) ? node567 : 1'b1;
														assign node567 = (inp[2]) ? 1'b1 : 1'b0;
													assign node570 = (inp[2]) ? 1'b0 : node571;
														assign node571 = (inp[14]) ? 1'b1 : 1'b0;
												assign node575 = (inp[14]) ? node577 : 1'b1;
													assign node577 = (inp[2]) ? 1'b1 : 1'b0;
											assign node580 = (inp[4]) ? node582 : 1'b0;
												assign node582 = (inp[14]) ? node588 : node583;
													assign node583 = (inp[13]) ? node585 : 1'b1;
														assign node585 = (inp[11]) ? 1'b1 : 1'b0;
													assign node588 = (inp[2]) ? node594 : node589;
														assign node589 = (inp[11]) ? 1'b0 : node590;
															assign node590 = (inp[13]) ? 1'b1 : 1'b0;
														assign node594 = (inp[11]) ? 1'b1 : 1'b0;
									assign node597 = (inp[0]) ? node599 : 1'b0;
										assign node599 = (inp[4]) ? 1'b0 : node600;
											assign node600 = (inp[13]) ? node606 : node601;
												assign node601 = (inp[14]) ? node603 : 1'b1;
													assign node603 = (inp[2]) ? 1'b1 : 1'b0;
												assign node606 = (inp[11]) ? node612 : node607;
													assign node607 = (inp[14]) ? node609 : 1'b0;
														assign node609 = (inp[2]) ? 1'b0 : 1'b1;
													assign node612 = (inp[14]) ? node614 : 1'b1;
														assign node614 = (inp[2]) ? 1'b1 : 1'b0;
								assign node618 = (inp[8]) ? node674 : node619;
									assign node619 = (inp[1]) ? node641 : node620;
										assign node620 = (inp[0]) ? node622 : 1'b1;
											assign node622 = (inp[4]) ? 1'b1 : node623;
												assign node623 = (inp[11]) ? node635 : node624;
													assign node624 = (inp[13]) ? node630 : node625;
														assign node625 = (inp[2]) ? 1'b0 : node626;
															assign node626 = (inp[14]) ? 1'b1 : 1'b0;
														assign node630 = (inp[14]) ? node632 : 1'b1;
															assign node632 = (inp[2]) ? 1'b1 : 1'b0;
													assign node635 = (inp[2]) ? 1'b0 : node636;
														assign node636 = (inp[14]) ? 1'b1 : 1'b0;
										assign node641 = (inp[14]) ? node655 : node642;
											assign node642 = (inp[11]) ? node650 : node643;
												assign node643 = (inp[13]) ? 1'b1 : node644;
													assign node644 = (inp[0]) ? node646 : 1'b0;
														assign node646 = (inp[4]) ? 1'b0 : 1'b1;
												assign node650 = (inp[0]) ? node652 : 1'b0;
													assign node652 = (inp[4]) ? 1'b0 : 1'b1;
											assign node655 = (inp[2]) ? node663 : node656;
												assign node656 = (inp[13]) ? node658 : 1'b1;
													assign node658 = (inp[11]) ? 1'b1 : node659;
														assign node659 = (inp[0]) ? 1'b1 : 1'b0;
												assign node663 = (inp[4]) ? node669 : node664;
													assign node664 = (inp[0]) ? 1'b1 : node665;
														assign node665 = (inp[13]) ? 1'b1 : 1'b0;
													assign node669 = (inp[13]) ? node671 : 1'b0;
														assign node671 = (inp[11]) ? 1'b0 : 1'b1;
									assign node674 = (inp[4]) ? 1'b1 : node675;
										assign node675 = (inp[0]) ? node677 : 1'b1;
											assign node677 = (inp[11]) ? node689 : node678;
												assign node678 = (inp[13]) ? node684 : node679;
													assign node679 = (inp[2]) ? 1'b0 : node680;
														assign node680 = (inp[14]) ? 1'b1 : 1'b0;
													assign node684 = (inp[2]) ? 1'b1 : node685;
														assign node685 = (inp[14]) ? 1'b0 : 1'b1;
												assign node689 = (inp[2]) ? 1'b0 : node690;
													assign node690 = (inp[14]) ? 1'b1 : 1'b0;
							assign node695 = (inp[4]) ? node755 : node696;
								assign node696 = (inp[0]) ? node718 : node697;
									assign node697 = (inp[1]) ? node699 : 1'b0;
										assign node699 = (inp[8]) ? 1'b0 : node700;
											assign node700 = (inp[13]) ? node706 : node701;
												assign node701 = (inp[2]) ? 1'b1 : node702;
													assign node702 = (inp[14]) ? 1'b0 : 1'b1;
												assign node706 = (inp[11]) ? node712 : node707;
													assign node707 = (inp[2]) ? 1'b0 : node708;
														assign node708 = (inp[14]) ? 1'b1 : 1'b0;
													assign node712 = (inp[2]) ? 1'b1 : node713;
														assign node713 = (inp[14]) ? 1'b0 : 1'b1;
									assign node718 = (inp[1]) ? node736 : node719;
										assign node719 = (inp[13]) ? node725 : node720;
											assign node720 = (inp[2]) ? 1'b1 : node721;
												assign node721 = (inp[14]) ? 1'b0 : 1'b1;
											assign node725 = (inp[11]) ? node731 : node726;
												assign node726 = (inp[2]) ? 1'b0 : node727;
													assign node727 = (inp[14]) ? 1'b1 : 1'b0;
												assign node731 = (inp[14]) ? node733 : 1'b1;
													assign node733 = (inp[2]) ? 1'b1 : 1'b0;
										assign node736 = (inp[8]) ? node738 : 1'b0;
											assign node738 = (inp[13]) ? node744 : node739;
												assign node739 = (inp[14]) ? node741 : 1'b1;
													assign node741 = (inp[2]) ? 1'b1 : 1'b0;
												assign node744 = (inp[11]) ? node750 : node745;
													assign node745 = (inp[14]) ? node747 : 1'b0;
														assign node747 = (inp[2]) ? 1'b0 : 1'b1;
													assign node750 = (inp[14]) ? node752 : 1'b1;
														assign node752 = (inp[2]) ? 1'b1 : 1'b0;
								assign node755 = (inp[8]) ? 1'b0 : node756;
									assign node756 = (inp[1]) ? node758 : 1'b0;
										assign node758 = (inp[13]) ? node764 : node759;
											assign node759 = (inp[14]) ? node761 : 1'b1;
												assign node761 = (inp[2]) ? 1'b1 : 1'b0;
											assign node764 = (inp[11]) ? node770 : node765;
												assign node765 = (inp[2]) ? 1'b0 : node766;
													assign node766 = (inp[14]) ? 1'b1 : 1'b0;
												assign node770 = (inp[2]) ? 1'b1 : node771;
													assign node771 = (inp[14]) ? 1'b0 : 1'b1;
					assign node776 = (inp[1]) ? node798 : node777;
						assign node777 = (inp[0]) ? node779 : 1'b1;
							assign node779 = (inp[4]) ? 1'b1 : node780;
								assign node780 = (inp[13]) ? node786 : node781;
									assign node781 = (inp[14]) ? node783 : 1'b0;
										assign node783 = (inp[2]) ? 1'b0 : 1'b1;
									assign node786 = (inp[11]) ? node792 : node787;
										assign node787 = (inp[14]) ? node789 : 1'b1;
											assign node789 = (inp[2]) ? 1'b1 : 1'b0;
										assign node792 = (inp[2]) ? 1'b0 : node793;
											assign node793 = (inp[14]) ? 1'b1 : 1'b0;
						assign node798 = (inp[8]) ? node836 : node799;
							assign node799 = (inp[0]) ? node817 : node800;
								assign node800 = (inp[2]) ? node812 : node801;
									assign node801 = (inp[14]) ? node807 : node802;
										assign node802 = (inp[11]) ? 1'b0 : node803;
											assign node803 = (inp[13]) ? 1'b1 : 1'b0;
										assign node807 = (inp[13]) ? node809 : 1'b1;
											assign node809 = (inp[11]) ? 1'b1 : 1'b0;
									assign node812 = (inp[11]) ? 1'b0 : node813;
										assign node813 = (inp[13]) ? 1'b1 : 1'b0;
								assign node817 = (inp[4]) ? node819 : 1'b1;
									assign node819 = (inp[13]) ? node825 : node820;
										assign node820 = (inp[2]) ? 1'b0 : node821;
											assign node821 = (inp[14]) ? 1'b1 : 1'b0;
										assign node825 = (inp[11]) ? node831 : node826;
											assign node826 = (inp[2]) ? 1'b1 : node827;
												assign node827 = (inp[14]) ? 1'b0 : 1'b1;
											assign node831 = (inp[2]) ? 1'b0 : node832;
												assign node832 = (inp[14]) ? 1'b1 : 1'b0;
							assign node836 = (inp[4]) ? 1'b1 : node837;
								assign node837 = (inp[0]) ? node839 : 1'b1;
									assign node839 = (inp[11]) ? node851 : node840;
										assign node840 = (inp[13]) ? node846 : node841;
											assign node841 = (inp[14]) ? node843 : 1'b0;
												assign node843 = (inp[2]) ? 1'b0 : 1'b1;
											assign node846 = (inp[2]) ? 1'b1 : node847;
												assign node847 = (inp[14]) ? 1'b0 : 1'b1;
										assign node851 = (inp[2]) ? 1'b0 : node852;
											assign node852 = (inp[14]) ? 1'b1 : 1'b0;
			assign node857 = (inp[15]) ? node1639 : node858;
				assign node858 = (inp[12]) ? node1558 : node859;
					assign node859 = (inp[7]) ? node1321 : node860;
						assign node860 = (inp[3]) ? node1096 : node861;
							assign node861 = (inp[9]) ? node941 : node862;
								assign node862 = (inp[0]) ? node884 : node863;
									assign node863 = (inp[1]) ? node865 : 1'b0;
										assign node865 = (inp[8]) ? 1'b0 : node866;
											assign node866 = (inp[13]) ? node872 : node867;
												assign node867 = (inp[14]) ? node869 : 1'b1;
													assign node869 = (inp[2]) ? 1'b1 : 1'b0;
												assign node872 = (inp[11]) ? node878 : node873;
													assign node873 = (inp[14]) ? node875 : 1'b0;
														assign node875 = (inp[2]) ? 1'b0 : 1'b1;
													assign node878 = (inp[14]) ? node880 : 1'b1;
														assign node880 = (inp[2]) ? 1'b1 : 1'b0;
									assign node884 = (inp[4]) ? node922 : node885;
										assign node885 = (inp[8]) ? node905 : node886;
											assign node886 = (inp[1]) ? 1'b0 : node887;
												assign node887 = (inp[2]) ? node899 : node888;
													assign node888 = (inp[14]) ? node894 : node889;
														assign node889 = (inp[11]) ? 1'b1 : node890;
															assign node890 = (inp[13]) ? 1'b0 : 1'b1;
														assign node894 = (inp[11]) ? 1'b0 : node895;
															assign node895 = (inp[13]) ? 1'b1 : 1'b0;
													assign node899 = (inp[11]) ? 1'b1 : node900;
														assign node900 = (inp[13]) ? 1'b0 : 1'b1;
											assign node905 = (inp[11]) ? node917 : node906;
												assign node906 = (inp[13]) ? node912 : node907;
													assign node907 = (inp[2]) ? 1'b1 : node908;
														assign node908 = (inp[14]) ? 1'b0 : 1'b1;
													assign node912 = (inp[14]) ? node914 : 1'b0;
														assign node914 = (inp[2]) ? 1'b0 : 1'b1;
												assign node917 = (inp[2]) ? 1'b1 : node918;
													assign node918 = (inp[14]) ? 1'b0 : 1'b1;
										assign node922 = (inp[8]) ? 1'b0 : node923;
											assign node923 = (inp[1]) ? node925 : 1'b0;
												assign node925 = (inp[11]) ? node935 : node926;
													assign node926 = (inp[13]) ? node932 : node927;
														assign node927 = (inp[14]) ? node929 : 1'b1;
															assign node929 = (inp[2]) ? 1'b1 : 1'b0;
														assign node932 = (inp[14]) ? 1'b1 : 1'b0;
													assign node935 = (inp[14]) ? node937 : 1'b1;
														assign node937 = (inp[2]) ? 1'b1 : 1'b0;
								assign node941 = (inp[10]) ? node1023 : node942;
									assign node942 = (inp[1]) ? node972 : node943;
										assign node943 = (inp[4]) ? 1'b1 : node944;
											assign node944 = (inp[0]) ? node946 : 1'b1;
												assign node946 = (inp[14]) ? node952 : node947;
													assign node947 = (inp[11]) ? 1'b0 : node948;
														assign node948 = (inp[13]) ? 1'b1 : 1'b0;
													assign node952 = (inp[8]) ? node962 : node953;
														assign node953 = (inp[13]) ? node955 : 1'b0;
															assign node955 = (inp[11]) ? node959 : node956;
																assign node956 = (inp[2]) ? 1'b1 : 1'b0;
																assign node959 = (inp[2]) ? 1'b0 : 1'b1;
														assign node962 = (inp[13]) ? node964 : 1'b1;
															assign node964 = (inp[2]) ? node968 : node965;
																assign node965 = (inp[11]) ? 1'b1 : 1'b0;
																assign node968 = (inp[11]) ? 1'b0 : 1'b1;
										assign node972 = (inp[8]) ? node1006 : node973;
											assign node973 = (inp[14]) ? node983 : node974;
												assign node974 = (inp[11]) ? node978 : node975;
													assign node975 = (inp[13]) ? 1'b1 : 1'b0;
													assign node978 = (inp[0]) ? node980 : 1'b0;
														assign node980 = (inp[4]) ? 1'b0 : 1'b1;
												assign node983 = (inp[4]) ? node995 : node984;
													assign node984 = (inp[0]) ? 1'b1 : node985;
														assign node985 = (inp[13]) ? node987 : 1'b1;
															assign node987 = (inp[11]) ? node991 : node988;
																assign node988 = (inp[2]) ? 1'b1 : 1'b0;
																assign node991 = (inp[2]) ? 1'b0 : 1'b1;
													assign node995 = (inp[2]) ? node1001 : node996;
														assign node996 = (inp[11]) ? 1'b1 : node997;
															assign node997 = (inp[13]) ? 1'b0 : 1'b1;
														assign node1001 = (inp[11]) ? 1'b0 : node1002;
															assign node1002 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1006 = (inp[0]) ? node1008 : 1'b1;
												assign node1008 = (inp[4]) ? 1'b1 : node1009;
													assign node1009 = (inp[13]) ? node1015 : node1010;
														assign node1010 = (inp[2]) ? 1'b0 : node1011;
															assign node1011 = (inp[14]) ? 1'b1 : 1'b0;
														assign node1015 = (inp[11]) ? node1017 : 1'b1;
															assign node1017 = (inp[14]) ? node1019 : 1'b0;
																assign node1019 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1023 = (inp[1]) ? node1045 : node1024;
										assign node1024 = (inp[0]) ? node1026 : 1'b0;
											assign node1026 = (inp[4]) ? 1'b0 : node1027;
												assign node1027 = (inp[11]) ? node1039 : node1028;
													assign node1028 = (inp[13]) ? node1034 : node1029;
														assign node1029 = (inp[14]) ? node1031 : 1'b1;
															assign node1031 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1034 = (inp[14]) ? node1036 : 1'b0;
															assign node1036 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1039 = (inp[14]) ? node1041 : 1'b1;
														assign node1041 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1045 = (inp[11]) ? node1071 : node1046;
											assign node1046 = (inp[13]) ? node1058 : node1047;
												assign node1047 = (inp[2]) ? node1053 : node1048;
													assign node1048 = (inp[0]) ? 1'b0 : node1049;
														assign node1049 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1053 = (inp[8]) ? node1055 : 1'b1;
														assign node1055 = (inp[0]) ? 1'b1 : 1'b0;
												assign node1058 = (inp[2]) ? 1'b0 : node1059;
													assign node1059 = (inp[14]) ? node1061 : 1'b0;
														assign node1061 = (inp[4]) ? 1'b0 : node1062;
															assign node1062 = (inp[8]) ? node1066 : node1063;
																assign node1063 = (inp[0]) ? 1'b0 : 1'b1;
																assign node1066 = (inp[0]) ? 1'b1 : 1'b0;
											assign node1071 = (inp[14]) ? node1083 : node1072;
												assign node1072 = (inp[8]) ? node1078 : node1073;
													assign node1073 = (inp[4]) ? 1'b1 : node1074;
														assign node1074 = (inp[0]) ? 1'b0 : 1'b1;
													assign node1078 = (inp[0]) ? node1080 : 1'b0;
														assign node1080 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1083 = (inp[2]) ? node1085 : 1'b0;
													assign node1085 = (inp[13]) ? node1091 : node1086;
														assign node1086 = (inp[8]) ? 1'b0 : node1087;
															assign node1087 = (inp[4]) ? 1'b1 : 1'b0;
														assign node1091 = (inp[8]) ? node1093 : 1'b1;
															assign node1093 = (inp[0]) ? 1'b1 : 1'b0;
							assign node1096 = (inp[9]) ? node1176 : node1097;
								assign node1097 = (inp[4]) ? node1155 : node1098;
									assign node1098 = (inp[0]) ? node1118 : node1099;
										assign node1099 = (inp[8]) ? 1'b1 : node1100;
											assign node1100 = (inp[1]) ? node1102 : 1'b1;
												assign node1102 = (inp[2]) ? node1112 : node1103;
													assign node1103 = (inp[11]) ? node1109 : node1104;
														assign node1104 = (inp[10]) ? 1'b1 : node1105;
															assign node1105 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1109 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1112 = (inp[13]) ? node1114 : 1'b0;
														assign node1114 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1118 = (inp[1]) ? node1136 : node1119;
											assign node1119 = (inp[13]) ? node1125 : node1120;
												assign node1120 = (inp[14]) ? node1122 : 1'b0;
													assign node1122 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1125 = (inp[11]) ? node1131 : node1126;
													assign node1126 = (inp[14]) ? node1128 : 1'b1;
														assign node1128 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1131 = (inp[2]) ? 1'b0 : node1132;
														assign node1132 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1136 = (inp[8]) ? node1138 : 1'b1;
												assign node1138 = (inp[14]) ? node1144 : node1139;
													assign node1139 = (inp[11]) ? 1'b0 : node1140;
														assign node1140 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1144 = (inp[2]) ? node1150 : node1145;
														assign node1145 = (inp[13]) ? node1147 : 1'b1;
															assign node1147 = (inp[11]) ? 1'b1 : 1'b0;
														assign node1150 = (inp[11]) ? 1'b0 : node1151;
															assign node1151 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1155 = (inp[8]) ? 1'b1 : node1156;
										assign node1156 = (inp[1]) ? node1158 : 1'b1;
											assign node1158 = (inp[13]) ? node1164 : node1159;
												assign node1159 = (inp[14]) ? node1161 : 1'b0;
													assign node1161 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1164 = (inp[11]) ? node1170 : node1165;
													assign node1165 = (inp[2]) ? 1'b1 : node1166;
														assign node1166 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1170 = (inp[14]) ? node1172 : 1'b0;
														assign node1172 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1176 = (inp[10]) ? node1252 : node1177;
									assign node1177 = (inp[8]) ? node1233 : node1178;
										assign node1178 = (inp[1]) ? node1198 : node1179;
											assign node1179 = (inp[4]) ? 1'b0 : node1180;
												assign node1180 = (inp[0]) ? node1182 : 1'b0;
													assign node1182 = (inp[2]) ? node1192 : node1183;
														assign node1183 = (inp[14]) ? node1187 : node1184;
															assign node1184 = (inp[13]) ? 1'b0 : 1'b1;
															assign node1187 = (inp[11]) ? 1'b0 : node1188;
																assign node1188 = (inp[13]) ? 1'b1 : 1'b0;
														assign node1192 = (inp[11]) ? 1'b1 : node1193;
															assign node1193 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1198 = (inp[4]) ? node1216 : node1199;
												assign node1199 = (inp[0]) ? 1'b0 : node1200;
													assign node1200 = (inp[14]) ? node1206 : node1201;
														assign node1201 = (inp[13]) ? node1203 : 1'b1;
															assign node1203 = (inp[11]) ? 1'b1 : 1'b0;
														assign node1206 = (inp[2]) ? node1212 : node1207;
															assign node1207 = (inp[13]) ? node1209 : 1'b0;
																assign node1209 = (inp[11]) ? 1'b0 : 1'b1;
															assign node1212 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1216 = (inp[14]) ? node1222 : node1217;
													assign node1217 = (inp[13]) ? node1219 : 1'b1;
														assign node1219 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1222 = (inp[2]) ? node1228 : node1223;
														assign node1223 = (inp[13]) ? node1225 : 1'b0;
															assign node1225 = (inp[11]) ? 1'b0 : 1'b1;
														assign node1228 = (inp[13]) ? node1230 : 1'b1;
															assign node1230 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1233 = (inp[4]) ? 1'b0 : node1234;
											assign node1234 = (inp[0]) ? node1236 : 1'b0;
												assign node1236 = (inp[11]) ? node1246 : node1237;
													assign node1237 = (inp[13]) ? node1243 : node1238;
														assign node1238 = (inp[14]) ? node1240 : 1'b1;
															assign node1240 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1243 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1246 = (inp[2]) ? 1'b1 : node1247;
														assign node1247 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1252 = (inp[1]) ? node1280 : node1253;
										assign node1253 = (inp[0]) ? node1255 : 1'b1;
											assign node1255 = (inp[4]) ? 1'b1 : node1256;
												assign node1256 = (inp[8]) ? node1270 : node1257;
													assign node1257 = (inp[13]) ? node1263 : node1258;
														assign node1258 = (inp[14]) ? node1260 : 1'b0;
															assign node1260 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1263 = (inp[14]) ? node1265 : 1'b1;
															assign node1265 = (inp[2]) ? 1'b1 : node1266;
																assign node1266 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1270 = (inp[2]) ? 1'b0 : node1271;
														assign node1271 = (inp[11]) ? 1'b0 : node1272;
															assign node1272 = (inp[14]) ? node1274 : 1'b1;
																assign node1274 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1280 = (inp[8]) ? node1308 : node1281;
											assign node1281 = (inp[2]) ? node1295 : node1282;
												assign node1282 = (inp[14]) ? 1'b1 : node1283;
													assign node1283 = (inp[4]) ? node1289 : node1284;
														assign node1284 = (inp[0]) ? 1'b1 : node1285;
															assign node1285 = (inp[11]) ? 1'b0 : 1'b1;
														assign node1289 = (inp[13]) ? node1291 : 1'b0;
															assign node1291 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1295 = (inp[11]) ? node1303 : node1296;
													assign node1296 = (inp[13]) ? 1'b1 : node1297;
														assign node1297 = (inp[4]) ? 1'b0 : node1298;
															assign node1298 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1303 = (inp[4]) ? 1'b0 : node1304;
														assign node1304 = (inp[0]) ? 1'b1 : 1'b0;
											assign node1308 = (inp[4]) ? 1'b1 : node1309;
												assign node1309 = (inp[0]) ? node1311 : 1'b1;
													assign node1311 = (inp[2]) ? 1'b0 : node1312;
														assign node1312 = (inp[14]) ? node1314 : 1'b0;
															assign node1314 = (inp[11]) ? 1'b1 : node1315;
																assign node1315 = (inp[13]) ? 1'b0 : 1'b1;
						assign node1321 = (inp[9]) ? node1403 : node1322;
							assign node1322 = (inp[4]) ? node1382 : node1323;
								assign node1323 = (inp[0]) ? node1345 : node1324;
									assign node1324 = (inp[8]) ? 1'b0 : node1325;
										assign node1325 = (inp[1]) ? node1327 : 1'b0;
											assign node1327 = (inp[2]) ? node1339 : node1328;
												assign node1328 = (inp[14]) ? node1334 : node1329;
													assign node1329 = (inp[13]) ? node1331 : 1'b1;
														assign node1331 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1334 = (inp[13]) ? node1336 : 1'b0;
														assign node1336 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1339 = (inp[11]) ? 1'b1 : node1340;
													assign node1340 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1345 = (inp[1]) ? node1363 : node1346;
										assign node1346 = (inp[2]) ? node1358 : node1347;
											assign node1347 = (inp[14]) ? node1353 : node1348;
												assign node1348 = (inp[13]) ? node1350 : 1'b1;
													assign node1350 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1353 = (inp[11]) ? 1'b0 : node1354;
													assign node1354 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1358 = (inp[11]) ? 1'b1 : node1359;
												assign node1359 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1363 = (inp[8]) ? node1365 : 1'b0;
											assign node1365 = (inp[2]) ? node1377 : node1366;
												assign node1366 = (inp[14]) ? node1372 : node1367;
													assign node1367 = (inp[11]) ? 1'b1 : node1368;
														assign node1368 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1372 = (inp[13]) ? node1374 : 1'b0;
														assign node1374 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1377 = (inp[13]) ? node1379 : 1'b1;
													assign node1379 = (inp[11]) ? 1'b1 : 1'b0;
								assign node1382 = (inp[8]) ? 1'b0 : node1383;
									assign node1383 = (inp[1]) ? node1385 : 1'b0;
										assign node1385 = (inp[2]) ? node1397 : node1386;
											assign node1386 = (inp[14]) ? node1392 : node1387;
												assign node1387 = (inp[11]) ? 1'b1 : node1388;
													assign node1388 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1392 = (inp[11]) ? 1'b0 : node1393;
													assign node1393 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1397 = (inp[13]) ? node1399 : 1'b1;
												assign node1399 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1403 = (inp[10]) ? node1481 : node1404;
								assign node1404 = (inp[1]) ? node1426 : node1405;
									assign node1405 = (inp[0]) ? node1407 : 1'b1;
										assign node1407 = (inp[4]) ? 1'b1 : node1408;
											assign node1408 = (inp[13]) ? node1414 : node1409;
												assign node1409 = (inp[14]) ? node1411 : 1'b0;
													assign node1411 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1414 = (inp[11]) ? node1420 : node1415;
													assign node1415 = (inp[14]) ? node1417 : 1'b1;
														assign node1417 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1420 = (inp[2]) ? 1'b0 : node1421;
														assign node1421 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1426 = (inp[8]) ? node1460 : node1427;
										assign node1427 = (inp[0]) ? node1445 : node1428;
											assign node1428 = (inp[2]) ? node1440 : node1429;
												assign node1429 = (inp[14]) ? node1435 : node1430;
													assign node1430 = (inp[13]) ? node1432 : 1'b0;
														assign node1432 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1435 = (inp[11]) ? 1'b1 : node1436;
														assign node1436 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1440 = (inp[13]) ? node1442 : 1'b0;
													assign node1442 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1445 = (inp[4]) ? node1447 : 1'b1;
												assign node1447 = (inp[13]) ? node1453 : node1448;
													assign node1448 = (inp[14]) ? node1450 : 1'b0;
														assign node1450 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1453 = (inp[11]) ? node1457 : node1454;
														assign node1454 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1457 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1460 = (inp[0]) ? node1462 : 1'b1;
											assign node1462 = (inp[4]) ? 1'b1 : node1463;
												assign node1463 = (inp[2]) ? node1475 : node1464;
													assign node1464 = (inp[14]) ? node1470 : node1465;
														assign node1465 = (inp[11]) ? 1'b0 : node1466;
															assign node1466 = (inp[13]) ? 1'b1 : 1'b0;
														assign node1470 = (inp[11]) ? 1'b1 : node1471;
															assign node1471 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1475 = (inp[13]) ? node1477 : 1'b0;
														assign node1477 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1481 = (inp[1]) ? node1503 : node1482;
									assign node1482 = (inp[0]) ? node1484 : 1'b0;
										assign node1484 = (inp[4]) ? 1'b0 : node1485;
											assign node1485 = (inp[14]) ? node1491 : node1486;
												assign node1486 = (inp[13]) ? node1488 : 1'b1;
													assign node1488 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1491 = (inp[2]) ? node1497 : node1492;
													assign node1492 = (inp[13]) ? node1494 : 1'b0;
														assign node1494 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1497 = (inp[13]) ? node1499 : 1'b1;
														assign node1499 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1503 = (inp[8]) ? node1537 : node1504;
										assign node1504 = (inp[0]) ? node1522 : node1505;
											assign node1505 = (inp[11]) ? node1517 : node1506;
												assign node1506 = (inp[13]) ? node1512 : node1507;
													assign node1507 = (inp[14]) ? node1509 : 1'b1;
														assign node1509 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1512 = (inp[14]) ? node1514 : 1'b0;
														assign node1514 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1517 = (inp[2]) ? 1'b1 : node1518;
													assign node1518 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1522 = (inp[4]) ? node1524 : 1'b0;
												assign node1524 = (inp[14]) ? node1530 : node1525;
													assign node1525 = (inp[13]) ? node1527 : 1'b1;
														assign node1527 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1530 = (inp[2]) ? node1532 : 1'b0;
														assign node1532 = (inp[11]) ? 1'b1 : node1533;
															assign node1533 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1537 = (inp[0]) ? node1539 : 1'b0;
											assign node1539 = (inp[4]) ? 1'b0 : node1540;
												assign node1540 = (inp[14]) ? node1546 : node1541;
													assign node1541 = (inp[11]) ? 1'b1 : node1542;
														assign node1542 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1546 = (inp[2]) ? node1552 : node1547;
														assign node1547 = (inp[11]) ? 1'b0 : node1548;
															assign node1548 = (inp[13]) ? 1'b1 : 1'b0;
														assign node1552 = (inp[11]) ? 1'b1 : node1553;
															assign node1553 = (inp[13]) ? 1'b0 : 1'b1;
					assign node1558 = (inp[1]) ? node1580 : node1559;
						assign node1559 = (inp[4]) ? 1'b1 : node1560;
							assign node1560 = (inp[0]) ? node1562 : 1'b1;
								assign node1562 = (inp[11]) ? node1574 : node1563;
									assign node1563 = (inp[13]) ? node1569 : node1564;
										assign node1564 = (inp[2]) ? 1'b0 : node1565;
											assign node1565 = (inp[14]) ? 1'b1 : 1'b0;
										assign node1569 = (inp[2]) ? 1'b1 : node1570;
											assign node1570 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1574 = (inp[14]) ? node1576 : 1'b0;
										assign node1576 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1580 = (inp[8]) ? node1618 : node1581;
							assign node1581 = (inp[4]) ? node1601 : node1582;
								assign node1582 = (inp[0]) ? 1'b1 : node1583;
									assign node1583 = (inp[14]) ? node1589 : node1584;
										assign node1584 = (inp[13]) ? node1586 : 1'b0;
											assign node1586 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1589 = (inp[2]) ? node1595 : node1590;
											assign node1590 = (inp[11]) ? 1'b1 : node1591;
												assign node1591 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1595 = (inp[11]) ? 1'b0 : node1596;
												assign node1596 = (inp[13]) ? 1'b1 : 1'b0;
								assign node1601 = (inp[11]) ? node1613 : node1602;
									assign node1602 = (inp[13]) ? node1608 : node1603;
										assign node1603 = (inp[14]) ? node1605 : 1'b0;
											assign node1605 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1608 = (inp[14]) ? node1610 : 1'b1;
											assign node1610 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1613 = (inp[2]) ? 1'b0 : node1614;
										assign node1614 = (inp[14]) ? 1'b1 : 1'b0;
							assign node1618 = (inp[4]) ? 1'b1 : node1619;
								assign node1619 = (inp[0]) ? node1621 : 1'b1;
									assign node1621 = (inp[2]) ? node1633 : node1622;
										assign node1622 = (inp[14]) ? node1628 : node1623;
											assign node1623 = (inp[11]) ? 1'b0 : node1624;
												assign node1624 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1628 = (inp[11]) ? 1'b1 : node1629;
												assign node1629 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1633 = (inp[13]) ? node1635 : 1'b0;
											assign node1635 = (inp[11]) ? 1'b0 : 1'b1;
				assign node1639 = (inp[7]) ? node2123 : node1640;
					assign node1640 = (inp[3]) ? node1884 : node1641;
						assign node1641 = (inp[9]) ? node1723 : node1642;
							assign node1642 = (inp[0]) ? node1664 : node1643;
								assign node1643 = (inp[1]) ? node1645 : 1'b0;
									assign node1645 = (inp[8]) ? 1'b0 : node1646;
										assign node1646 = (inp[11]) ? node1658 : node1647;
											assign node1647 = (inp[13]) ? node1653 : node1648;
												assign node1648 = (inp[2]) ? 1'b1 : node1649;
													assign node1649 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1653 = (inp[2]) ? 1'b0 : node1654;
													assign node1654 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1658 = (inp[14]) ? node1660 : 1'b1;
												assign node1660 = (inp[2]) ? 1'b1 : 1'b0;
								assign node1664 = (inp[4]) ? node1702 : node1665;
									assign node1665 = (inp[1]) ? node1683 : node1666;
										assign node1666 = (inp[11]) ? node1678 : node1667;
											assign node1667 = (inp[13]) ? node1673 : node1668;
												assign node1668 = (inp[14]) ? node1670 : 1'b1;
													assign node1670 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1673 = (inp[14]) ? node1675 : 1'b0;
													assign node1675 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1678 = (inp[2]) ? 1'b1 : node1679;
												assign node1679 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1683 = (inp[8]) ? node1685 : 1'b0;
											assign node1685 = (inp[14]) ? node1691 : node1686;
												assign node1686 = (inp[11]) ? 1'b1 : node1687;
													assign node1687 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1691 = (inp[2]) ? node1697 : node1692;
													assign node1692 = (inp[13]) ? node1694 : 1'b0;
														assign node1694 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1697 = (inp[13]) ? node1699 : 1'b1;
														assign node1699 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1702 = (inp[1]) ? node1704 : 1'b0;
										assign node1704 = (inp[8]) ? 1'b0 : node1705;
											assign node1705 = (inp[14]) ? node1711 : node1706;
												assign node1706 = (inp[13]) ? node1708 : 1'b1;
													assign node1708 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1711 = (inp[2]) ? node1717 : node1712;
													assign node1712 = (inp[13]) ? node1714 : 1'b0;
														assign node1714 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1717 = (inp[11]) ? 1'b1 : node1718;
														assign node1718 = (inp[13]) ? 1'b0 : 1'b1;
							assign node1723 = (inp[10]) ? node1805 : node1724;
								assign node1724 = (inp[0]) ? node1746 : node1725;
									assign node1725 = (inp[8]) ? 1'b1 : node1726;
										assign node1726 = (inp[1]) ? node1728 : 1'b1;
											assign node1728 = (inp[2]) ? node1740 : node1729;
												assign node1729 = (inp[14]) ? node1735 : node1730;
													assign node1730 = (inp[11]) ? 1'b0 : node1731;
														assign node1731 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1735 = (inp[13]) ? node1737 : 1'b1;
														assign node1737 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1740 = (inp[11]) ? 1'b0 : node1741;
													assign node1741 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1746 = (inp[4]) ? node1784 : node1747;
										assign node1747 = (inp[13]) ? node1761 : node1748;
											assign node1748 = (inp[2]) ? node1756 : node1749;
												assign node1749 = (inp[14]) ? 1'b1 : node1750;
													assign node1750 = (inp[8]) ? 1'b0 : node1751;
														assign node1751 = (inp[1]) ? 1'b1 : 1'b0;
												assign node1756 = (inp[8]) ? 1'b0 : node1757;
													assign node1757 = (inp[1]) ? 1'b1 : 1'b0;
											assign node1761 = (inp[1]) ? node1773 : node1762;
												assign node1762 = (inp[11]) ? node1768 : node1763;
													assign node1763 = (inp[2]) ? 1'b1 : node1764;
														assign node1764 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1768 = (inp[2]) ? 1'b0 : node1769;
														assign node1769 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1773 = (inp[8]) ? node1775 : 1'b1;
													assign node1775 = (inp[11]) ? node1781 : node1776;
														assign node1776 = (inp[2]) ? 1'b1 : node1777;
															assign node1777 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1781 = (inp[14]) ? 1'b1 : 1'b0;
										assign node1784 = (inp[8]) ? 1'b1 : node1785;
											assign node1785 = (inp[1]) ? node1787 : 1'b1;
												assign node1787 = (inp[11]) ? node1799 : node1788;
													assign node1788 = (inp[13]) ? node1794 : node1789;
														assign node1789 = (inp[2]) ? 1'b0 : node1790;
															assign node1790 = (inp[14]) ? 1'b1 : 1'b0;
														assign node1794 = (inp[2]) ? 1'b1 : node1795;
															assign node1795 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1799 = (inp[2]) ? 1'b0 : node1800;
														assign node1800 = (inp[14]) ? 1'b1 : 1'b0;
								assign node1805 = (inp[1]) ? node1827 : node1806;
									assign node1806 = (inp[4]) ? 1'b0 : node1807;
										assign node1807 = (inp[0]) ? node1809 : 1'b0;
											assign node1809 = (inp[14]) ? node1815 : node1810;
												assign node1810 = (inp[11]) ? 1'b1 : node1811;
													assign node1811 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1815 = (inp[2]) ? node1821 : node1816;
													assign node1816 = (inp[13]) ? node1818 : 1'b0;
														assign node1818 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1821 = (inp[13]) ? node1823 : 1'b1;
														assign node1823 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1827 = (inp[8]) ? node1865 : node1828;
										assign node1828 = (inp[4]) ? node1848 : node1829;
											assign node1829 = (inp[0]) ? 1'b0 : node1830;
												assign node1830 = (inp[11]) ? node1842 : node1831;
													assign node1831 = (inp[13]) ? node1837 : node1832;
														assign node1832 = (inp[14]) ? node1834 : 1'b1;
															assign node1834 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1837 = (inp[14]) ? node1839 : 1'b0;
															assign node1839 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1842 = (inp[2]) ? 1'b1 : node1843;
														assign node1843 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1848 = (inp[14]) ? node1854 : node1849;
												assign node1849 = (inp[13]) ? node1851 : 1'b1;
													assign node1851 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1854 = (inp[2]) ? node1860 : node1855;
													assign node1855 = (inp[11]) ? 1'b0 : node1856;
														assign node1856 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1860 = (inp[11]) ? 1'b1 : node1861;
														assign node1861 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1865 = (inp[0]) ? node1867 : 1'b0;
											assign node1867 = (inp[4]) ? 1'b0 : node1868;
												assign node1868 = (inp[11]) ? node1878 : node1869;
													assign node1869 = (inp[13]) ? node1873 : node1870;
														assign node1870 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1873 = (inp[14]) ? node1875 : 1'b0;
															assign node1875 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1878 = (inp[14]) ? node1880 : 1'b1;
														assign node1880 = (inp[2]) ? 1'b1 : 1'b0;
						assign node1884 = (inp[10]) ? node2042 : node1885;
							assign node1885 = (inp[9]) ? node1961 : node1886;
								assign node1886 = (inp[8]) ? node1940 : node1887;
									assign node1887 = (inp[1]) ? node1907 : node1888;
										assign node1888 = (inp[4]) ? 1'b1 : node1889;
											assign node1889 = (inp[0]) ? node1891 : 1'b1;
												assign node1891 = (inp[2]) ? node1901 : node1892;
													assign node1892 = (inp[14]) ? node1898 : node1893;
														assign node1893 = (inp[11]) ? 1'b0 : node1894;
															assign node1894 = (inp[12]) ? 1'b1 : 1'b0;
														assign node1898 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1901 = (inp[13]) ? node1903 : 1'b0;
														assign node1903 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1907 = (inp[4]) ? node1923 : node1908;
											assign node1908 = (inp[0]) ? 1'b1 : node1909;
												assign node1909 = (inp[11]) ? node1917 : node1910;
													assign node1910 = (inp[13]) ? node1912 : 1'b0;
														assign node1912 = (inp[14]) ? node1914 : 1'b1;
															assign node1914 = (inp[12]) ? 1'b1 : 1'b0;
													assign node1917 = (inp[2]) ? 1'b0 : node1918;
														assign node1918 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1923 = (inp[13]) ? node1929 : node1924;
												assign node1924 = (inp[14]) ? node1926 : 1'b0;
													assign node1926 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1929 = (inp[11]) ? node1935 : node1930;
													assign node1930 = (inp[2]) ? 1'b1 : node1931;
														assign node1931 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1935 = (inp[2]) ? 1'b0 : node1936;
														assign node1936 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1940 = (inp[4]) ? 1'b1 : node1941;
										assign node1941 = (inp[0]) ? node1943 : 1'b1;
											assign node1943 = (inp[2]) ? node1955 : node1944;
												assign node1944 = (inp[14]) ? node1950 : node1945;
													assign node1945 = (inp[11]) ? 1'b0 : node1946;
														assign node1946 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1950 = (inp[11]) ? 1'b1 : node1951;
														assign node1951 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1955 = (inp[13]) ? node1957 : 1'b0;
													assign node1957 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1961 = (inp[1]) ? node1985 : node1962;
									assign node1962 = (inp[4]) ? 1'b0 : node1963;
										assign node1963 = (inp[0]) ? node1965 : 1'b0;
											assign node1965 = (inp[2]) ? node1979 : node1966;
												assign node1966 = (inp[14]) ? node1974 : node1967;
													assign node1967 = (inp[12]) ? node1969 : 1'b1;
														assign node1969 = (inp[11]) ? 1'b1 : node1970;
															assign node1970 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1974 = (inp[13]) ? node1976 : 1'b0;
														assign node1976 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1979 = (inp[11]) ? 1'b1 : node1980;
													assign node1980 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1985 = (inp[8]) ? node2021 : node1986;
										assign node1986 = (inp[0]) ? node2002 : node1987;
											assign node1987 = (inp[2]) ? node1997 : node1988;
												assign node1988 = (inp[14]) ? node1992 : node1989;
													assign node1989 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1992 = (inp[11]) ? 1'b0 : node1993;
														assign node1993 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1997 = (inp[11]) ? 1'b1 : node1998;
													assign node1998 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2002 = (inp[4]) ? node2004 : 1'b0;
												assign node2004 = (inp[14]) ? node2010 : node2005;
													assign node2005 = (inp[13]) ? node2007 : 1'b1;
														assign node2007 = (inp[11]) ? 1'b1 : 1'b0;
													assign node2010 = (inp[2]) ? node2016 : node2011;
														assign node2011 = (inp[13]) ? node2013 : 1'b0;
															assign node2013 = (inp[12]) ? 1'b1 : 1'b0;
														assign node2016 = (inp[11]) ? 1'b1 : node2017;
															assign node2017 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2021 = (inp[0]) ? node2023 : 1'b0;
											assign node2023 = (inp[4]) ? 1'b0 : node2024;
												assign node2024 = (inp[13]) ? node2030 : node2025;
													assign node2025 = (inp[14]) ? node2027 : 1'b1;
														assign node2027 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2030 = (inp[11]) ? node2036 : node2031;
														assign node2031 = (inp[14]) ? node2033 : 1'b0;
															assign node2033 = (inp[2]) ? 1'b0 : 1'b1;
														assign node2036 = (inp[12]) ? node2038 : 1'b1;
															assign node2038 = (inp[14]) ? 1'b0 : 1'b1;
							assign node2042 = (inp[1]) ? node2064 : node2043;
								assign node2043 = (inp[0]) ? node2045 : 1'b1;
									assign node2045 = (inp[4]) ? 1'b1 : node2046;
										assign node2046 = (inp[11]) ? node2058 : node2047;
											assign node2047 = (inp[13]) ? node2053 : node2048;
												assign node2048 = (inp[14]) ? node2050 : 1'b0;
													assign node2050 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2053 = (inp[14]) ? node2055 : 1'b1;
													assign node2055 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2058 = (inp[2]) ? 1'b0 : node2059;
												assign node2059 = (inp[14]) ? 1'b1 : 1'b0;
								assign node2064 = (inp[8]) ? node2102 : node2065;
									assign node2065 = (inp[0]) ? node2083 : node2066;
										assign node2066 = (inp[11]) ? node2078 : node2067;
											assign node2067 = (inp[13]) ? node2073 : node2068;
												assign node2068 = (inp[2]) ? 1'b0 : node2069;
													assign node2069 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2073 = (inp[2]) ? 1'b1 : node2074;
													assign node2074 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2078 = (inp[14]) ? node2080 : 1'b0;
												assign node2080 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2083 = (inp[4]) ? node2085 : 1'b1;
											assign node2085 = (inp[14]) ? node2091 : node2086;
												assign node2086 = (inp[11]) ? 1'b0 : node2087;
													assign node2087 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2091 = (inp[2]) ? node2097 : node2092;
													assign node2092 = (inp[13]) ? node2094 : 1'b1;
														assign node2094 = (inp[11]) ? 1'b1 : 1'b0;
													assign node2097 = (inp[13]) ? node2099 : 1'b0;
														assign node2099 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2102 = (inp[0]) ? node2104 : 1'b1;
										assign node2104 = (inp[4]) ? 1'b1 : node2105;
											assign node2105 = (inp[14]) ? node2111 : node2106;
												assign node2106 = (inp[13]) ? node2108 : 1'b0;
													assign node2108 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2111 = (inp[2]) ? node2117 : node2112;
													assign node2112 = (inp[13]) ? node2114 : 1'b1;
														assign node2114 = (inp[11]) ? 1'b1 : 1'b0;
													assign node2117 = (inp[11]) ? 1'b0 : node2118;
														assign node2118 = (inp[13]) ? 1'b1 : 1'b0;
					assign node2123 = (inp[9]) ? node2205 : node2124;
						assign node2124 = (inp[1]) ? node2146 : node2125;
							assign node2125 = (inp[4]) ? 1'b0 : node2126;
								assign node2126 = (inp[0]) ? node2128 : 1'b0;
									assign node2128 = (inp[11]) ? node2140 : node2129;
										assign node2129 = (inp[13]) ? node2135 : node2130;
											assign node2130 = (inp[14]) ? node2132 : 1'b1;
												assign node2132 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2135 = (inp[14]) ? node2137 : 1'b0;
												assign node2137 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2140 = (inp[2]) ? 1'b1 : node2141;
											assign node2141 = (inp[14]) ? 1'b0 : 1'b1;
							assign node2146 = (inp[8]) ? node2184 : node2147;
								assign node2147 = (inp[0]) ? node2165 : node2148;
									assign node2148 = (inp[14]) ? node2154 : node2149;
										assign node2149 = (inp[13]) ? node2151 : 1'b1;
											assign node2151 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2154 = (inp[2]) ? node2160 : node2155;
											assign node2155 = (inp[11]) ? 1'b0 : node2156;
												assign node2156 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2160 = (inp[11]) ? 1'b1 : node2161;
												assign node2161 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2165 = (inp[4]) ? node2167 : 1'b0;
										assign node2167 = (inp[11]) ? node2179 : node2168;
											assign node2168 = (inp[13]) ? node2174 : node2169;
												assign node2169 = (inp[2]) ? 1'b1 : node2170;
													assign node2170 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2174 = (inp[2]) ? 1'b0 : node2175;
													assign node2175 = (inp[14]) ? 1'b1 : 1'b0;
											assign node2179 = (inp[2]) ? 1'b1 : node2180;
												assign node2180 = (inp[14]) ? 1'b0 : 1'b1;
								assign node2184 = (inp[0]) ? node2186 : 1'b0;
									assign node2186 = (inp[4]) ? 1'b0 : node2187;
										assign node2187 = (inp[2]) ? node2199 : node2188;
											assign node2188 = (inp[14]) ? node2194 : node2189;
												assign node2189 = (inp[13]) ? node2191 : 1'b1;
													assign node2191 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2194 = (inp[11]) ? 1'b0 : node2195;
													assign node2195 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2199 = (inp[13]) ? node2201 : 1'b1;
												assign node2201 = (inp[11]) ? 1'b1 : 1'b0;
						assign node2205 = (inp[10]) ? node2287 : node2206;
							assign node2206 = (inp[4]) ? node2266 : node2207;
								assign node2207 = (inp[0]) ? node2229 : node2208;
									assign node2208 = (inp[1]) ? node2210 : 1'b1;
										assign node2210 = (inp[8]) ? 1'b1 : node2211;
											assign node2211 = (inp[2]) ? node2223 : node2212;
												assign node2212 = (inp[14]) ? node2218 : node2213;
													assign node2213 = (inp[13]) ? node2215 : 1'b0;
														assign node2215 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2218 = (inp[13]) ? node2220 : 1'b1;
														assign node2220 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2223 = (inp[13]) ? node2225 : 1'b0;
													assign node2225 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2229 = (inp[8]) ? node2249 : node2230;
										assign node2230 = (inp[1]) ? 1'b1 : node2231;
											assign node2231 = (inp[14]) ? node2237 : node2232;
												assign node2232 = (inp[11]) ? 1'b0 : node2233;
													assign node2233 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2237 = (inp[2]) ? node2243 : node2238;
													assign node2238 = (inp[11]) ? 1'b1 : node2239;
														assign node2239 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2243 = (inp[11]) ? 1'b0 : node2244;
														assign node2244 = (inp[13]) ? 1'b1 : 1'b0;
										assign node2249 = (inp[2]) ? node2261 : node2250;
											assign node2250 = (inp[14]) ? node2256 : node2251;
												assign node2251 = (inp[13]) ? node2253 : 1'b0;
													assign node2253 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2256 = (inp[13]) ? node2258 : 1'b1;
													assign node2258 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2261 = (inp[11]) ? 1'b0 : node2262;
												assign node2262 = (inp[13]) ? 1'b1 : 1'b0;
								assign node2266 = (inp[8]) ? 1'b1 : node2267;
									assign node2267 = (inp[1]) ? node2269 : 1'b1;
										assign node2269 = (inp[11]) ? node2281 : node2270;
											assign node2270 = (inp[13]) ? node2276 : node2271;
												assign node2271 = (inp[2]) ? 1'b0 : node2272;
													assign node2272 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2276 = (inp[14]) ? node2278 : 1'b1;
													assign node2278 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2281 = (inp[2]) ? 1'b0 : node2282;
												assign node2282 = (inp[14]) ? 1'b1 : 1'b0;
							assign node2287 = (inp[4]) ? node2353 : node2288;
								assign node2288 = (inp[0]) ? node2310 : node2289;
									assign node2289 = (inp[8]) ? 1'b0 : node2290;
										assign node2290 = (inp[1]) ? node2292 : 1'b0;
											assign node2292 = (inp[13]) ? node2298 : node2293;
												assign node2293 = (inp[14]) ? node2295 : 1'b1;
													assign node2295 = (inp[2]) ? 1'b1 : 1'b0;
												assign node2298 = (inp[11]) ? node2304 : node2299;
													assign node2299 = (inp[14]) ? node2301 : 1'b0;
														assign node2301 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2304 = (inp[2]) ? 1'b1 : node2305;
														assign node2305 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2310 = (inp[8]) ? node2336 : node2311;
										assign node2311 = (inp[1]) ? 1'b0 : node2312;
											assign node2312 = (inp[14]) ? node2318 : node2313;
												assign node2313 = (inp[11]) ? 1'b1 : node2314;
													assign node2314 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2318 = (inp[11]) ? node2332 : node2319;
													assign node2319 = (inp[12]) ? node2327 : node2320;
														assign node2320 = (inp[2]) ? node2324 : node2321;
															assign node2321 = (inp[13]) ? 1'b1 : 1'b0;
															assign node2324 = (inp[13]) ? 1'b0 : 1'b1;
														assign node2327 = (inp[2]) ? node2329 : 1'b1;
															assign node2329 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2332 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2336 = (inp[2]) ? node2348 : node2337;
											assign node2337 = (inp[14]) ? node2343 : node2338;
												assign node2338 = (inp[11]) ? 1'b1 : node2339;
													assign node2339 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2343 = (inp[11]) ? 1'b0 : node2344;
													assign node2344 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2348 = (inp[11]) ? 1'b1 : node2349;
												assign node2349 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2353 = (inp[8]) ? 1'b0 : node2354;
									assign node2354 = (inp[1]) ? node2356 : 1'b0;
										assign node2356 = (inp[2]) ? node2368 : node2357;
											assign node2357 = (inp[14]) ? node2363 : node2358;
												assign node2358 = (inp[11]) ? 1'b1 : node2359;
													assign node2359 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2363 = (inp[13]) ? node2365 : 1'b0;
													assign node2365 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2368 = (inp[13]) ? node2370 : 1'b1;
												assign node2370 = (inp[11]) ? 1'b1 : 1'b0;
		assign node2374 = (inp[12]) ? node2456 : node2375;
			assign node2375 = (inp[1]) ? node2397 : node2376;
				assign node2376 = (inp[4]) ? 1'b1 : node2377;
					assign node2377 = (inp[0]) ? node2379 : 1'b1;
						assign node2379 = (inp[14]) ? node2385 : node2380;
							assign node2380 = (inp[11]) ? 1'b0 : node2381;
								assign node2381 = (inp[13]) ? 1'b1 : 1'b0;
							assign node2385 = (inp[2]) ? node2391 : node2386;
								assign node2386 = (inp[11]) ? 1'b1 : node2387;
									assign node2387 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2391 = (inp[13]) ? node2393 : 1'b0;
									assign node2393 = (inp[11]) ? 1'b0 : 1'b1;
				assign node2397 = (inp[8]) ? node2435 : node2398;
					assign node2398 = (inp[0]) ? node2416 : node2399;
						assign node2399 = (inp[2]) ? node2411 : node2400;
							assign node2400 = (inp[14]) ? node2406 : node2401;
								assign node2401 = (inp[11]) ? 1'b0 : node2402;
									assign node2402 = (inp[13]) ? 1'b1 : 1'b0;
								assign node2406 = (inp[13]) ? node2408 : 1'b1;
									assign node2408 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2411 = (inp[13]) ? node2413 : 1'b0;
								assign node2413 = (inp[11]) ? 1'b0 : 1'b1;
						assign node2416 = (inp[4]) ? node2418 : 1'b1;
							assign node2418 = (inp[14]) ? node2424 : node2419;
								assign node2419 = (inp[11]) ? 1'b0 : node2420;
									assign node2420 = (inp[13]) ? 1'b1 : 1'b0;
								assign node2424 = (inp[2]) ? node2430 : node2425;
									assign node2425 = (inp[13]) ? node2427 : 1'b1;
										assign node2427 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2430 = (inp[11]) ? 1'b0 : node2431;
										assign node2431 = (inp[13]) ? 1'b1 : 1'b0;
					assign node2435 = (inp[0]) ? node2437 : 1'b1;
						assign node2437 = (inp[4]) ? 1'b1 : node2438;
							assign node2438 = (inp[2]) ? node2450 : node2439;
								assign node2439 = (inp[14]) ? node2445 : node2440;
									assign node2440 = (inp[11]) ? 1'b0 : node2441;
										assign node2441 = (inp[13]) ? 1'b1 : 1'b0;
									assign node2445 = (inp[13]) ? node2447 : 1'b1;
										assign node2447 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2450 = (inp[13]) ? node2452 : 1'b0;
									assign node2452 = (inp[11]) ? 1'b0 : 1'b1;
			assign node2456 = (inp[15]) ? node3200 : node2457;
				assign node2457 = (inp[3]) ? node2705 : node2458;
					assign node2458 = (inp[10]) ? node2624 : node2459;
						assign node2459 = (inp[9]) ? node2543 : node2460;
							assign node2460 = (inp[1]) ? node2482 : node2461;
								assign node2461 = (inp[0]) ? node2463 : 1'b0;
									assign node2463 = (inp[4]) ? 1'b0 : node2464;
										assign node2464 = (inp[14]) ? node2470 : node2465;
											assign node2465 = (inp[13]) ? node2467 : 1'b1;
												assign node2467 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2470 = (inp[2]) ? node2476 : node2471;
												assign node2471 = (inp[13]) ? node2473 : 1'b0;
													assign node2473 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2476 = (inp[11]) ? 1'b1 : node2477;
													assign node2477 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2482 = (inp[8]) ? node2522 : node2483;
									assign node2483 = (inp[4]) ? node2505 : node2484;
										assign node2484 = (inp[0]) ? 1'b0 : node2485;
											assign node2485 = (inp[11]) ? node2499 : node2486;
												assign node2486 = (inp[13]) ? node2494 : node2487;
													assign node2487 = (inp[6]) ? 1'b1 : node2488;
														assign node2488 = (inp[14]) ? node2490 : 1'b1;
															assign node2490 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2494 = (inp[2]) ? 1'b0 : node2495;
														assign node2495 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2499 = (inp[14]) ? node2501 : 1'b1;
													assign node2501 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2505 = (inp[2]) ? node2517 : node2506;
											assign node2506 = (inp[14]) ? node2512 : node2507;
												assign node2507 = (inp[13]) ? node2509 : 1'b1;
													assign node2509 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2512 = (inp[13]) ? node2514 : 1'b0;
													assign node2514 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2517 = (inp[13]) ? node2519 : 1'b1;
												assign node2519 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2522 = (inp[4]) ? 1'b0 : node2523;
										assign node2523 = (inp[0]) ? node2525 : 1'b0;
											assign node2525 = (inp[13]) ? node2531 : node2526;
												assign node2526 = (inp[14]) ? node2528 : 1'b1;
													assign node2528 = (inp[2]) ? 1'b1 : 1'b0;
												assign node2531 = (inp[11]) ? node2537 : node2532;
													assign node2532 = (inp[2]) ? 1'b0 : node2533;
														assign node2533 = (inp[14]) ? 1'b1 : 1'b0;
													assign node2537 = (inp[14]) ? node2539 : 1'b1;
														assign node2539 = (inp[2]) ? 1'b1 : 1'b0;
							assign node2543 = (inp[0]) ? node2565 : node2544;
								assign node2544 = (inp[1]) ? node2546 : 1'b1;
									assign node2546 = (inp[8]) ? 1'b1 : node2547;
										assign node2547 = (inp[11]) ? node2559 : node2548;
											assign node2548 = (inp[13]) ? node2554 : node2549;
												assign node2549 = (inp[14]) ? node2551 : 1'b0;
													assign node2551 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2554 = (inp[2]) ? 1'b1 : node2555;
													assign node2555 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2559 = (inp[2]) ? 1'b0 : node2560;
												assign node2560 = (inp[14]) ? 1'b1 : 1'b0;
								assign node2565 = (inp[4]) ? node2603 : node2566;
									assign node2566 = (inp[8]) ? node2586 : node2567;
										assign node2567 = (inp[1]) ? 1'b1 : node2568;
											assign node2568 = (inp[13]) ? node2574 : node2569;
												assign node2569 = (inp[2]) ? 1'b0 : node2570;
													assign node2570 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2574 = (inp[11]) ? node2580 : node2575;
													assign node2575 = (inp[2]) ? 1'b1 : node2576;
														assign node2576 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2580 = (inp[2]) ? 1'b0 : node2581;
														assign node2581 = (inp[14]) ? 1'b1 : 1'b0;
										assign node2586 = (inp[13]) ? node2592 : node2587;
											assign node2587 = (inp[14]) ? node2589 : 1'b0;
												assign node2589 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2592 = (inp[11]) ? node2598 : node2593;
												assign node2593 = (inp[14]) ? node2595 : 1'b1;
													assign node2595 = (inp[2]) ? 1'b1 : 1'b0;
												assign node2598 = (inp[14]) ? node2600 : 1'b0;
													assign node2600 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2603 = (inp[8]) ? 1'b1 : node2604;
										assign node2604 = (inp[1]) ? node2606 : 1'b1;
											assign node2606 = (inp[2]) ? node2618 : node2607;
												assign node2607 = (inp[14]) ? node2613 : node2608;
													assign node2608 = (inp[13]) ? node2610 : 1'b0;
														assign node2610 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2613 = (inp[13]) ? node2615 : 1'b1;
														assign node2615 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2618 = (inp[13]) ? node2620 : 1'b0;
													assign node2620 = (inp[11]) ? 1'b0 : 1'b1;
						assign node2624 = (inp[4]) ? node2684 : node2625;
							assign node2625 = (inp[0]) ? node2647 : node2626;
								assign node2626 = (inp[8]) ? 1'b0 : node2627;
									assign node2627 = (inp[1]) ? node2629 : 1'b0;
										assign node2629 = (inp[2]) ? node2641 : node2630;
											assign node2630 = (inp[14]) ? node2636 : node2631;
												assign node2631 = (inp[11]) ? 1'b1 : node2632;
													assign node2632 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2636 = (inp[13]) ? node2638 : 1'b0;
													assign node2638 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2641 = (inp[11]) ? 1'b1 : node2642;
												assign node2642 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2647 = (inp[1]) ? node2665 : node2648;
									assign node2648 = (inp[13]) ? node2654 : node2649;
										assign node2649 = (inp[2]) ? 1'b1 : node2650;
											assign node2650 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2654 = (inp[11]) ? node2660 : node2655;
											assign node2655 = (inp[2]) ? 1'b0 : node2656;
												assign node2656 = (inp[14]) ? 1'b1 : 1'b0;
											assign node2660 = (inp[2]) ? 1'b1 : node2661;
												assign node2661 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2665 = (inp[8]) ? node2667 : 1'b0;
										assign node2667 = (inp[11]) ? node2679 : node2668;
											assign node2668 = (inp[13]) ? node2674 : node2669;
												assign node2669 = (inp[2]) ? 1'b1 : node2670;
													assign node2670 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2674 = (inp[14]) ? node2676 : 1'b0;
													assign node2676 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2679 = (inp[14]) ? node2681 : 1'b1;
												assign node2681 = (inp[2]) ? 1'b1 : 1'b0;
							assign node2684 = (inp[8]) ? 1'b0 : node2685;
								assign node2685 = (inp[1]) ? node2687 : 1'b0;
									assign node2687 = (inp[13]) ? node2693 : node2688;
										assign node2688 = (inp[2]) ? 1'b1 : node2689;
											assign node2689 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2693 = (inp[11]) ? node2699 : node2694;
											assign node2694 = (inp[2]) ? 1'b0 : node2695;
												assign node2695 = (inp[14]) ? 1'b1 : 1'b0;
											assign node2699 = (inp[2]) ? 1'b1 : node2700;
												assign node2700 = (inp[14]) ? 1'b0 : 1'b1;
					assign node2705 = (inp[7]) ? node2955 : node2706;
						assign node2706 = (inp[9]) ? node2796 : node2707;
							assign node2707 = (inp[8]) ? node2775 : node2708;
								assign node2708 = (inp[1]) ? node2738 : node2709;
									assign node2709 = (inp[0]) ? node2711 : 1'b1;
										assign node2711 = (inp[4]) ? 1'b1 : node2712;
											assign node2712 = (inp[11]) ? node2732 : node2713;
												assign node2713 = (inp[10]) ? node2723 : node2714;
													assign node2714 = (inp[2]) ? 1'b0 : node2715;
														assign node2715 = (inp[13]) ? node2719 : node2716;
															assign node2716 = (inp[14]) ? 1'b1 : 1'b0;
															assign node2719 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2723 = (inp[13]) ? node2727 : node2724;
														assign node2724 = (inp[2]) ? 1'b0 : 1'b1;
														assign node2727 = (inp[14]) ? node2729 : 1'b1;
															assign node2729 = (inp[2]) ? 1'b1 : 1'b0;
												assign node2732 = (inp[14]) ? node2734 : 1'b0;
													assign node2734 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2738 = (inp[4]) ? node2758 : node2739;
										assign node2739 = (inp[0]) ? 1'b1 : node2740;
											assign node2740 = (inp[2]) ? node2752 : node2741;
												assign node2741 = (inp[14]) ? node2747 : node2742;
													assign node2742 = (inp[11]) ? 1'b0 : node2743;
														assign node2743 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2747 = (inp[11]) ? 1'b1 : node2748;
														assign node2748 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2752 = (inp[13]) ? node2754 : 1'b0;
													assign node2754 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2758 = (inp[2]) ? node2770 : node2759;
											assign node2759 = (inp[14]) ? node2765 : node2760;
												assign node2760 = (inp[13]) ? node2762 : 1'b0;
													assign node2762 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2765 = (inp[11]) ? 1'b1 : node2766;
													assign node2766 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2770 = (inp[13]) ? node2772 : 1'b0;
												assign node2772 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2775 = (inp[0]) ? node2777 : 1'b1;
									assign node2777 = (inp[4]) ? 1'b1 : node2778;
										assign node2778 = (inp[2]) ? node2790 : node2779;
											assign node2779 = (inp[14]) ? node2785 : node2780;
												assign node2780 = (inp[11]) ? 1'b0 : node2781;
													assign node2781 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2785 = (inp[13]) ? node2787 : 1'b1;
													assign node2787 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2790 = (inp[11]) ? 1'b0 : node2791;
												assign node2791 = (inp[13]) ? 1'b1 : 1'b0;
							assign node2796 = (inp[10]) ? node2874 : node2797;
								assign node2797 = (inp[8]) ? node2853 : node2798;
									assign node2798 = (inp[1]) ? node2816 : node2799;
										assign node2799 = (inp[0]) ? node2801 : 1'b0;
											assign node2801 = (inp[4]) ? 1'b0 : node2802;
												assign node2802 = (inp[11]) ? node2810 : node2803;
													assign node2803 = (inp[13]) ? 1'b0 : node2804;
														assign node2804 = (inp[2]) ? 1'b1 : node2805;
															assign node2805 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2810 = (inp[2]) ? 1'b1 : node2811;
														assign node2811 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2816 = (inp[0]) ? node2834 : node2817;
											assign node2817 = (inp[2]) ? node2829 : node2818;
												assign node2818 = (inp[14]) ? node2824 : node2819;
													assign node2819 = (inp[13]) ? node2821 : 1'b1;
														assign node2821 = (inp[4]) ? 1'b0 : 1'b1;
													assign node2824 = (inp[11]) ? 1'b0 : node2825;
														assign node2825 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2829 = (inp[13]) ? node2831 : 1'b1;
													assign node2831 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2834 = (inp[4]) ? node2836 : 1'b0;
												assign node2836 = (inp[14]) ? node2842 : node2837;
													assign node2837 = (inp[11]) ? 1'b1 : node2838;
														assign node2838 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2842 = (inp[2]) ? node2848 : node2843;
														assign node2843 = (inp[13]) ? node2845 : 1'b0;
															assign node2845 = (inp[11]) ? 1'b0 : 1'b1;
														assign node2848 = (inp[13]) ? node2850 : 1'b1;
															assign node2850 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2853 = (inp[0]) ? node2855 : 1'b0;
										assign node2855 = (inp[4]) ? 1'b0 : node2856;
											assign node2856 = (inp[11]) ? node2868 : node2857;
												assign node2857 = (inp[13]) ? node2863 : node2858;
													assign node2858 = (inp[2]) ? 1'b1 : node2859;
														assign node2859 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2863 = (inp[14]) ? node2865 : 1'b0;
														assign node2865 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2868 = (inp[14]) ? node2870 : 1'b1;
													assign node2870 = (inp[2]) ? 1'b1 : 1'b0;
								assign node2874 = (inp[1]) ? node2896 : node2875;
									assign node2875 = (inp[0]) ? node2877 : 1'b1;
										assign node2877 = (inp[4]) ? 1'b1 : node2878;
											assign node2878 = (inp[2]) ? node2890 : node2879;
												assign node2879 = (inp[14]) ? node2885 : node2880;
													assign node2880 = (inp[11]) ? 1'b0 : node2881;
														assign node2881 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2885 = (inp[11]) ? 1'b1 : node2886;
														assign node2886 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2890 = (inp[13]) ? node2892 : 1'b0;
													assign node2892 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2896 = (inp[8]) ? node2934 : node2897;
										assign node2897 = (inp[4]) ? node2917 : node2898;
											assign node2898 = (inp[0]) ? 1'b1 : node2899;
												assign node2899 = (inp[14]) ? node2905 : node2900;
													assign node2900 = (inp[11]) ? 1'b0 : node2901;
														assign node2901 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2905 = (inp[2]) ? node2911 : node2906;
														assign node2906 = (inp[13]) ? node2908 : 1'b1;
															assign node2908 = (inp[11]) ? 1'b1 : 1'b0;
														assign node2911 = (inp[11]) ? 1'b0 : node2912;
															assign node2912 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2917 = (inp[2]) ? node2929 : node2918;
												assign node2918 = (inp[14]) ? node2924 : node2919;
													assign node2919 = (inp[13]) ? node2921 : 1'b0;
														assign node2921 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2924 = (inp[11]) ? 1'b1 : node2925;
														assign node2925 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2929 = (inp[11]) ? 1'b0 : node2930;
													assign node2930 = (inp[13]) ? 1'b1 : 1'b0;
										assign node2934 = (inp[4]) ? 1'b1 : node2935;
											assign node2935 = (inp[0]) ? node2937 : 1'b1;
												assign node2937 = (inp[11]) ? node2949 : node2938;
													assign node2938 = (inp[13]) ? node2944 : node2939;
														assign node2939 = (inp[14]) ? node2941 : 1'b0;
															assign node2941 = (inp[2]) ? 1'b0 : 1'b1;
														assign node2944 = (inp[2]) ? 1'b1 : node2945;
															assign node2945 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2949 = (inp[14]) ? node2951 : 1'b0;
														assign node2951 = (inp[2]) ? 1'b0 : 1'b1;
						assign node2955 = (inp[10]) ? node3121 : node2956;
							assign node2956 = (inp[9]) ? node3038 : node2957;
								assign node2957 = (inp[0]) ? node2979 : node2958;
									assign node2958 = (inp[1]) ? node2960 : 1'b0;
										assign node2960 = (inp[8]) ? 1'b0 : node2961;
											assign node2961 = (inp[13]) ? node2967 : node2962;
												assign node2962 = (inp[2]) ? 1'b1 : node2963;
													assign node2963 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2967 = (inp[11]) ? node2973 : node2968;
													assign node2968 = (inp[2]) ? 1'b0 : node2969;
														assign node2969 = (inp[14]) ? 1'b1 : 1'b0;
													assign node2973 = (inp[14]) ? node2975 : 1'b1;
														assign node2975 = (inp[2]) ? 1'b1 : 1'b0;
									assign node2979 = (inp[4]) ? node3017 : node2980;
										assign node2980 = (inp[8]) ? node3000 : node2981;
											assign node2981 = (inp[1]) ? 1'b0 : node2982;
												assign node2982 = (inp[11]) ? node2994 : node2983;
													assign node2983 = (inp[13]) ? node2989 : node2984;
														assign node2984 = (inp[14]) ? node2986 : 1'b1;
															assign node2986 = (inp[2]) ? 1'b1 : 1'b0;
														assign node2989 = (inp[14]) ? node2991 : 1'b0;
															assign node2991 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2994 = (inp[2]) ? 1'b1 : node2995;
														assign node2995 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3000 = (inp[2]) ? node3012 : node3001;
												assign node3001 = (inp[14]) ? node3007 : node3002;
													assign node3002 = (inp[13]) ? node3004 : 1'b1;
														assign node3004 = (inp[11]) ? 1'b1 : 1'b0;
													assign node3007 = (inp[13]) ? node3009 : 1'b0;
														assign node3009 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3012 = (inp[11]) ? 1'b1 : node3013;
													assign node3013 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3017 = (inp[8]) ? 1'b0 : node3018;
											assign node3018 = (inp[1]) ? node3020 : 1'b0;
												assign node3020 = (inp[14]) ? node3026 : node3021;
													assign node3021 = (inp[11]) ? 1'b1 : node3022;
														assign node3022 = (inp[13]) ? 1'b0 : 1'b1;
													assign node3026 = (inp[2]) ? node3032 : node3027;
														assign node3027 = (inp[11]) ? 1'b0 : node3028;
															assign node3028 = (inp[13]) ? 1'b1 : 1'b0;
														assign node3032 = (inp[11]) ? 1'b1 : node3033;
															assign node3033 = (inp[13]) ? 1'b0 : 1'b1;
								assign node3038 = (inp[8]) ? node3098 : node3039;
									assign node3039 = (inp[1]) ? node3061 : node3040;
										assign node3040 = (inp[0]) ? node3042 : 1'b1;
											assign node3042 = (inp[4]) ? 1'b1 : node3043;
												assign node3043 = (inp[13]) ? node3049 : node3044;
													assign node3044 = (inp[14]) ? node3046 : 1'b0;
														assign node3046 = (inp[2]) ? 1'b0 : 1'b1;
													assign node3049 = (inp[11]) ? node3055 : node3050;
														assign node3050 = (inp[14]) ? node3052 : 1'b1;
															assign node3052 = (inp[2]) ? 1'b1 : 1'b0;
														assign node3055 = (inp[14]) ? node3057 : 1'b0;
															assign node3057 = (inp[6]) ? 1'b1 : 1'b0;
										assign node3061 = (inp[4]) ? node3081 : node3062;
											assign node3062 = (inp[0]) ? 1'b1 : node3063;
												assign node3063 = (inp[11]) ? node3075 : node3064;
													assign node3064 = (inp[13]) ? node3070 : node3065;
														assign node3065 = (inp[2]) ? 1'b0 : node3066;
															assign node3066 = (inp[14]) ? 1'b1 : 1'b0;
														assign node3070 = (inp[2]) ? 1'b1 : node3071;
															assign node3071 = (inp[14]) ? 1'b0 : 1'b1;
													assign node3075 = (inp[14]) ? node3077 : 1'b0;
														assign node3077 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3081 = (inp[14]) ? node3087 : node3082;
												assign node3082 = (inp[11]) ? 1'b0 : node3083;
													assign node3083 = (inp[13]) ? 1'b1 : 1'b0;
												assign node3087 = (inp[2]) ? node3093 : node3088;
													assign node3088 = (inp[13]) ? node3090 : 1'b1;
														assign node3090 = (inp[11]) ? 1'b1 : 1'b0;
													assign node3093 = (inp[13]) ? node3095 : 1'b0;
														assign node3095 = (inp[0]) ? 1'b1 : 1'b0;
									assign node3098 = (inp[4]) ? 1'b1 : node3099;
										assign node3099 = (inp[0]) ? node3101 : 1'b1;
											assign node3101 = (inp[2]) ? node3115 : node3102;
												assign node3102 = (inp[14]) ? node3108 : node3103;
													assign node3103 = (inp[11]) ? 1'b0 : node3104;
														assign node3104 = (inp[13]) ? 1'b1 : 1'b0;
													assign node3108 = (inp[6]) ? 1'b1 : node3109;
														assign node3109 = (inp[13]) ? node3111 : 1'b1;
															assign node3111 = (inp[11]) ? 1'b1 : 1'b0;
												assign node3115 = (inp[13]) ? node3117 : 1'b0;
													assign node3117 = (inp[11]) ? 1'b0 : 1'b1;
							assign node3121 = (inp[8]) ? node3179 : node3122;
								assign node3122 = (inp[1]) ? node3144 : node3123;
									assign node3123 = (inp[4]) ? 1'b0 : node3124;
										assign node3124 = (inp[0]) ? node3126 : 1'b0;
											assign node3126 = (inp[2]) ? node3138 : node3127;
												assign node3127 = (inp[14]) ? node3133 : node3128;
													assign node3128 = (inp[11]) ? 1'b1 : node3129;
														assign node3129 = (inp[13]) ? 1'b0 : 1'b1;
													assign node3133 = (inp[11]) ? 1'b0 : node3134;
														assign node3134 = (inp[13]) ? 1'b1 : 1'b0;
												assign node3138 = (inp[11]) ? 1'b1 : node3139;
													assign node3139 = (inp[13]) ? 1'b0 : 1'b1;
									assign node3144 = (inp[4]) ? node3162 : node3145;
										assign node3145 = (inp[0]) ? 1'b0 : node3146;
											assign node3146 = (inp[14]) ? node3152 : node3147;
												assign node3147 = (inp[13]) ? node3149 : 1'b1;
													assign node3149 = (inp[11]) ? 1'b1 : 1'b0;
												assign node3152 = (inp[2]) ? node3158 : node3153;
													assign node3153 = (inp[13]) ? node3155 : 1'b0;
														assign node3155 = (inp[11]) ? 1'b0 : 1'b1;
													assign node3158 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3162 = (inp[11]) ? node3174 : node3163;
											assign node3163 = (inp[13]) ? node3169 : node3164;
												assign node3164 = (inp[2]) ? 1'b1 : node3165;
													assign node3165 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3169 = (inp[2]) ? 1'b0 : node3170;
													assign node3170 = (inp[14]) ? 1'b1 : 1'b0;
											assign node3174 = (inp[14]) ? node3176 : 1'b1;
												assign node3176 = (inp[2]) ? 1'b1 : 1'b0;
								assign node3179 = (inp[4]) ? 1'b0 : node3180;
									assign node3180 = (inp[0]) ? node3182 : 1'b0;
										assign node3182 = (inp[14]) ? node3188 : node3183;
											assign node3183 = (inp[11]) ? 1'b1 : node3184;
												assign node3184 = (inp[13]) ? 1'b0 : 1'b1;
											assign node3188 = (inp[2]) ? node3194 : node3189;
												assign node3189 = (inp[13]) ? node3191 : 1'b0;
													assign node3191 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3194 = (inp[11]) ? 1'b1 : node3195;
													assign node3195 = (inp[13]) ? 1'b0 : 1'b1;
				assign node3200 = (inp[8]) ? node3260 : node3201;
					assign node3201 = (inp[1]) ? node3223 : node3202;
						assign node3202 = (inp[0]) ? node3204 : 1'b1;
							assign node3204 = (inp[4]) ? 1'b1 : node3205;
								assign node3205 = (inp[14]) ? node3211 : node3206;
									assign node3206 = (inp[13]) ? node3208 : 1'b0;
										assign node3208 = (inp[11]) ? 1'b0 : 1'b1;
									assign node3211 = (inp[2]) ? node3217 : node3212;
										assign node3212 = (inp[13]) ? node3214 : 1'b1;
											assign node3214 = (inp[11]) ? 1'b1 : 1'b0;
										assign node3217 = (inp[13]) ? node3219 : 1'b0;
											assign node3219 = (inp[11]) ? 1'b0 : 1'b1;
						assign node3223 = (inp[4]) ? node3243 : node3224;
							assign node3224 = (inp[0]) ? 1'b1 : node3225;
								assign node3225 = (inp[13]) ? node3231 : node3226;
									assign node3226 = (inp[2]) ? 1'b0 : node3227;
										assign node3227 = (inp[14]) ? 1'b1 : 1'b0;
									assign node3231 = (inp[11]) ? node3237 : node3232;
										assign node3232 = (inp[2]) ? 1'b1 : node3233;
											assign node3233 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3237 = (inp[14]) ? node3239 : 1'b0;
											assign node3239 = (inp[2]) ? 1'b0 : 1'b1;
							assign node3243 = (inp[11]) ? node3255 : node3244;
								assign node3244 = (inp[13]) ? node3250 : node3245;
									assign node3245 = (inp[2]) ? 1'b0 : node3246;
										assign node3246 = (inp[14]) ? 1'b1 : 1'b0;
									assign node3250 = (inp[2]) ? 1'b1 : node3251;
										assign node3251 = (inp[14]) ? 1'b0 : 1'b1;
								assign node3255 = (inp[2]) ? 1'b0 : node3256;
									assign node3256 = (inp[14]) ? 1'b1 : 1'b0;
					assign node3260 = (inp[0]) ? node3262 : 1'b1;
						assign node3262 = (inp[4]) ? 1'b1 : node3263;
							assign node3263 = (inp[2]) ? node3275 : node3264;
								assign node3264 = (inp[14]) ? node3270 : node3265;
									assign node3265 = (inp[11]) ? 1'b0 : node3266;
										assign node3266 = (inp[13]) ? 1'b1 : 1'b0;
									assign node3270 = (inp[11]) ? 1'b1 : node3271;
										assign node3271 = (inp[13]) ? 1'b0 : 1'b1;
								assign node3275 = (inp[13]) ? node3277 : 1'b0;
									assign node3277 = (inp[11]) ? 1'b0 : 1'b1;

endmodule