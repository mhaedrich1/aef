module dtc_split875_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node465;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node639;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node700;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node754;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node839;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node856;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node997;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1021;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1038;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1136;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1175;
	wire [3-1:0] node1177;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1189;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1201;
	wire [3-1:0] node1204;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1261;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1384;
	wire [3-1:0] node1386;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1392;
	wire [3-1:0] node1393;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1403;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1426;
	wire [3-1:0] node1428;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1443;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1479;
	wire [3-1:0] node1481;
	wire [3-1:0] node1484;
	wire [3-1:0] node1486;
	wire [3-1:0] node1488;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1499;
	wire [3-1:0] node1502;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1535;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1542;
	wire [3-1:0] node1544;
	wire [3-1:0] node1547;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1553;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1561;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1571;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1579;
	wire [3-1:0] node1581;
	wire [3-1:0] node1584;
	wire [3-1:0] node1585;
	wire [3-1:0] node1586;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1593;
	wire [3-1:0] node1595;

	assign outp = (inp[6]) ? node546 : node1;
		assign node1 = (inp[9]) ? node375 : node2;
			assign node2 = (inp[3]) ? node242 : node3;
				assign node3 = (inp[0]) ? node41 : node4;
					assign node4 = (inp[7]) ? node26 : node5;
						assign node5 = (inp[10]) ? node15 : node6;
							assign node6 = (inp[5]) ? node8 : 3'b000;
								assign node8 = (inp[8]) ? 3'b000 : node9;
									assign node9 = (inp[11]) ? node11 : 3'b010;
										assign node11 = (inp[4]) ? 3'b010 : 3'b000;
							assign node15 = (inp[8]) ? node23 : node16;
								assign node16 = (inp[5]) ? node18 : 3'b010;
									assign node18 = (inp[11]) ? node20 : 3'b100;
										assign node20 = (inp[4]) ? 3'b100 : 3'b110;
								assign node23 = (inp[5]) ? 3'b010 : 3'b000;
						assign node26 = (inp[8]) ? 3'b000 : node27;
							assign node27 = (inp[5]) ? node29 : 3'b000;
								assign node29 = (inp[10]) ? node37 : node30;
									assign node30 = (inp[4]) ? node32 : 3'b000;
										assign node32 = (inp[2]) ? node34 : 3'b000;
											assign node34 = (inp[11]) ? 3'b000 : 3'b010;
									assign node37 = (inp[4]) ? 3'b000 : 3'b010;
					assign node41 = (inp[10]) ? node171 : node42;
						assign node42 = (inp[7]) ? node102 : node43;
							assign node43 = (inp[4]) ? node69 : node44;
								assign node44 = (inp[11]) ? node56 : node45;
									assign node45 = (inp[8]) ? node51 : node46;
										assign node46 = (inp[5]) ? node48 : 3'b110;
											assign node48 = (inp[1]) ? 3'b100 : 3'b000;
										assign node51 = (inp[5]) ? 3'b110 : node52;
											assign node52 = (inp[1]) ? 3'b110 : 3'b100;
									assign node56 = (inp[1]) ? node64 : node57;
										assign node57 = (inp[5]) ? node61 : node58;
											assign node58 = (inp[8]) ? 3'b100 : 3'b010;
											assign node61 = (inp[8]) ? 3'b010 : 3'b000;
										assign node64 = (inp[5]) ? 3'b010 : node65;
											assign node65 = (inp[8]) ? 3'b110 : 3'b010;
								assign node69 = (inp[1]) ? node87 : node70;
									assign node70 = (inp[11]) ? node80 : node71;
										assign node71 = (inp[2]) ? node73 : 3'b000;
											assign node73 = (inp[5]) ? node77 : node74;
												assign node74 = (inp[8]) ? 3'b000 : 3'b110;
												assign node77 = (inp[8]) ? 3'b110 : 3'b000;
										assign node80 = (inp[8]) ? node84 : node81;
											assign node81 = (inp[5]) ? 3'b000 : 3'b110;
											assign node84 = (inp[5]) ? 3'b110 : 3'b100;
									assign node87 = (inp[11]) ? node93 : node88;
										assign node88 = (inp[8]) ? node90 : 3'b100;
											assign node90 = (inp[5]) ? 3'b100 : 3'b010;
										assign node93 = (inp[5]) ? node99 : node94;
											assign node94 = (inp[8]) ? node96 : 3'b100;
												assign node96 = (inp[2]) ? 3'b100 : 3'b000;
											assign node99 = (inp[8]) ? 3'b100 : 3'b000;
							assign node102 = (inp[4]) ? node124 : node103;
								assign node103 = (inp[1]) ? node115 : node104;
									assign node104 = (inp[5]) ? node110 : node105;
										assign node105 = (inp[8]) ? 3'b010 : node106;
											assign node106 = (inp[11]) ? 3'b000 : 3'b001;
										assign node110 = (inp[8]) ? node112 : 3'b100;
											assign node112 = (inp[11]) ? 3'b000 : 3'b001;
									assign node115 = (inp[5]) ? node121 : node116;
										assign node116 = (inp[8]) ? node118 : 3'b001;
											assign node118 = (inp[11]) ? 3'b000 : 3'b100;
										assign node121 = (inp[8]) ? 3'b001 : 3'b110;
								assign node124 = (inp[1]) ? node148 : node125;
									assign node125 = (inp[11]) ? node141 : node126;
										assign node126 = (inp[2]) ? node134 : node127;
											assign node127 = (inp[8]) ? node131 : node128;
												assign node128 = (inp[5]) ? 3'b000 : 3'b001;
												assign node131 = (inp[5]) ? 3'b001 : 3'b100;
											assign node134 = (inp[5]) ? node138 : node135;
												assign node135 = (inp[8]) ? 3'b000 : 3'b111;
												assign node138 = (inp[8]) ? 3'b111 : 3'b000;
										assign node141 = (inp[5]) ? node145 : node142;
											assign node142 = (inp[8]) ? 3'b000 : 3'b010;
											assign node145 = (inp[8]) ? 3'b010 : 3'b100;
									assign node148 = (inp[2]) ? node158 : node149;
										assign node149 = (inp[8]) ? node155 : node150;
											assign node150 = (inp[5]) ? node152 : 3'b010;
												assign node152 = (inp[11]) ? 3'b000 : 3'b010;
											assign node155 = (inp[5]) ? 3'b010 : 3'b110;
										assign node158 = (inp[8]) ? node166 : node159;
											assign node159 = (inp[11]) ? node163 : node160;
												assign node160 = (inp[5]) ? 3'b010 : 3'b110;
												assign node163 = (inp[5]) ? 3'b100 : 3'b010;
											assign node166 = (inp[5]) ? node168 : 3'b110;
												assign node168 = (inp[11]) ? 3'b010 : 3'b110;
						assign node171 = (inp[7]) ? node203 : node172;
							assign node172 = (inp[4]) ? node194 : node173;
								assign node173 = (inp[1]) ? node183 : node174;
									assign node174 = (inp[11]) ? node176 : 3'b000;
										assign node176 = (inp[8]) ? node180 : node177;
											assign node177 = (inp[5]) ? 3'b000 : 3'b100;
											assign node180 = (inp[5]) ? 3'b100 : 3'b000;
									assign node183 = (inp[5]) ? node189 : node184;
										assign node184 = (inp[11]) ? node186 : 3'b010;
											assign node186 = (inp[8]) ? 3'b010 : 3'b100;
										assign node189 = (inp[8]) ? node191 : 3'b100;
											assign node191 = (inp[2]) ? 3'b010 : 3'b100;
								assign node194 = (inp[2]) ? node196 : 3'b000;
									assign node196 = (inp[11]) ? 3'b000 : node197;
										assign node197 = (inp[5]) ? 3'b000 : node198;
											assign node198 = (inp[8]) ? 3'b100 : 3'b000;
							assign node203 = (inp[4]) ? node223 : node204;
								assign node204 = (inp[1]) ? node210 : node205;
									assign node205 = (inp[5]) ? node207 : 3'b100;
										assign node207 = (inp[8]) ? 3'b100 : 3'b000;
									assign node210 = (inp[11]) ? node218 : node211;
										assign node211 = (inp[8]) ? node215 : node212;
											assign node212 = (inp[5]) ? 3'b010 : 3'b110;
											assign node215 = (inp[5]) ? 3'b110 : 3'b000;
										assign node218 = (inp[5]) ? node220 : 3'b110;
											assign node220 = (inp[8]) ? 3'b110 : 3'b010;
								assign node223 = (inp[8]) ? node231 : node224;
									assign node224 = (inp[5]) ? node228 : node225;
										assign node225 = (inp[1]) ? 3'b000 : 3'b010;
										assign node228 = (inp[11]) ? 3'b000 : 3'b100;
									assign node231 = (inp[5]) ? node237 : node232;
										assign node232 = (inp[11]) ? node234 : 3'b000;
											assign node234 = (inp[1]) ? 3'b010 : 3'b110;
										assign node237 = (inp[11]) ? node239 : 3'b010;
											assign node239 = (inp[1]) ? 3'b000 : 3'b010;
				assign node242 = (inp[7]) ? node274 : node243;
					assign node243 = (inp[4]) ? 3'b000 : node244;
						assign node244 = (inp[5]) ? 3'b000 : node245;
							assign node245 = (inp[11]) ? node263 : node246;
								assign node246 = (inp[1]) ? node254 : node247;
									assign node247 = (inp[0]) ? node249 : 3'b000;
										assign node249 = (inp[8]) ? node251 : 3'b000;
											assign node251 = (inp[10]) ? 3'b000 : 3'b100;
									assign node254 = (inp[0]) ? node258 : node255;
										assign node255 = (inp[8]) ? 3'b000 : 3'b100;
										assign node258 = (inp[10]) ? 3'b000 : node259;
											assign node259 = (inp[8]) ? 3'b100 : 3'b000;
								assign node263 = (inp[10]) ? 3'b000 : node264;
									assign node264 = (inp[1]) ? node266 : 3'b000;
										assign node266 = (inp[0]) ? 3'b000 : node267;
											assign node267 = (inp[8]) ? 3'b000 : 3'b100;
					assign node274 = (inp[8]) ? node314 : node275;
						assign node275 = (inp[0]) ? node299 : node276;
							assign node276 = (inp[4]) ? node288 : node277;
								assign node277 = (inp[1]) ? node283 : node278;
									assign node278 = (inp[10]) ? 3'b000 : node279;
										assign node279 = (inp[5]) ? 3'b010 : 3'b000;
									assign node283 = (inp[5]) ? node285 : 3'b010;
										assign node285 = (inp[10]) ? 3'b100 : 3'b110;
								assign node288 = (inp[11]) ? 3'b000 : node289;
									assign node289 = (inp[10]) ? 3'b000 : node290;
										assign node290 = (inp[1]) ? node294 : node291;
											assign node291 = (inp[5]) ? 3'b010 : 3'b000;
											assign node294 = (inp[5]) ? 3'b100 : 3'b010;
							assign node299 = (inp[5]) ? 3'b000 : node300;
								assign node300 = (inp[10]) ? 3'b000 : node301;
									assign node301 = (inp[11]) ? node307 : node302;
										assign node302 = (inp[4]) ? node304 : 3'b100;
											assign node304 = (inp[1]) ? 3'b000 : 3'b100;
										assign node307 = (inp[1]) ? node309 : 3'b000;
											assign node309 = (inp[4]) ? 3'b000 : 3'b100;
						assign node314 = (inp[0]) ? node348 : node315;
							assign node315 = (inp[5]) ? node317 : 3'b100;
								assign node317 = (inp[1]) ? node333 : node318;
									assign node318 = (inp[2]) ? node326 : node319;
										assign node319 = (inp[10]) ? node323 : node320;
											assign node320 = (inp[11]) ? 3'b100 : 3'b000;
											assign node323 = (inp[11]) ? 3'b000 : 3'b100;
										assign node326 = (inp[10]) ? node330 : node327;
											assign node327 = (inp[11]) ? 3'b100 : 3'b000;
											assign node330 = (inp[11]) ? 3'b000 : 3'b100;
									assign node333 = (inp[4]) ? node341 : node334;
										assign node334 = (inp[11]) ? node338 : node335;
											assign node335 = (inp[10]) ? 3'b110 : 3'b010;
											assign node338 = (inp[10]) ? 3'b010 : 3'b110;
										assign node341 = (inp[11]) ? node345 : node342;
											assign node342 = (inp[10]) ? 3'b100 : 3'b010;
											assign node345 = (inp[10]) ? 3'b000 : 3'b100;
							assign node348 = (inp[10]) ? node368 : node349;
								assign node349 = (inp[4]) ? node361 : node350;
									assign node350 = (inp[5]) ? node356 : node351;
										assign node351 = (inp[11]) ? 3'b100 : node352;
											assign node352 = (inp[1]) ? 3'b010 : 3'b110;
										assign node356 = (inp[11]) ? node358 : 3'b100;
											assign node358 = (inp[1]) ? 3'b100 : 3'b000;
									assign node361 = (inp[1]) ? 3'b000 : node362;
										assign node362 = (inp[5]) ? node364 : 3'b100;
											assign node364 = (inp[11]) ? 3'b000 : 3'b100;
								assign node368 = (inp[1]) ? node370 : 3'b000;
									assign node370 = (inp[5]) ? 3'b000 : node371;
										assign node371 = (inp[4]) ? 3'b000 : 3'b100;
			assign node375 = (inp[7]) ? node429 : node376;
				assign node376 = (inp[3]) ? 3'b000 : node377;
					assign node377 = (inp[0]) ? node391 : node378;
						assign node378 = (inp[10]) ? 3'b000 : node379;
							assign node379 = (inp[1]) ? node381 : 3'b000;
								assign node381 = (inp[4]) ? 3'b000 : node382;
									assign node382 = (inp[8]) ? 3'b000 : node383;
										assign node383 = (inp[11]) ? 3'b000 : node384;
											assign node384 = (inp[5]) ? 3'b010 : 3'b000;
						assign node391 = (inp[5]) ? node417 : node392;
							assign node392 = (inp[10]) ? node408 : node393;
								assign node393 = (inp[4]) ? node401 : node394;
									assign node394 = (inp[8]) ? 3'b100 : node395;
										assign node395 = (inp[11]) ? 3'b000 : node396;
											assign node396 = (inp[1]) ? 3'b100 : 3'b000;
									assign node401 = (inp[2]) ? node403 : 3'b000;
										assign node403 = (inp[8]) ? node405 : 3'b000;
											assign node405 = (inp[11]) ? 3'b100 : 3'b000;
								assign node408 = (inp[4]) ? node410 : 3'b000;
									assign node410 = (inp[11]) ? 3'b000 : node411;
										assign node411 = (inp[2]) ? node413 : 3'b000;
											assign node413 = (inp[8]) ? 3'b100 : 3'b000;
							assign node417 = (inp[11]) ? 3'b000 : node418;
								assign node418 = (inp[8]) ? node420 : 3'b000;
									assign node420 = (inp[4]) ? 3'b000 : node421;
										assign node421 = (inp[10]) ? 3'b000 : node422;
											assign node422 = (inp[1]) ? 3'b100 : 3'b000;
				assign node429 = (inp[3]) ? node519 : node430;
					assign node430 = (inp[0]) ? node446 : node431;
						assign node431 = (inp[5]) ? node433 : 3'b000;
							assign node433 = (inp[8]) ? 3'b000 : node434;
								assign node434 = (inp[4]) ? node438 : node435;
									assign node435 = (inp[10]) ? 3'b010 : 3'b000;
									assign node438 = (inp[11]) ? 3'b000 : node439;
										assign node439 = (inp[10]) ? 3'b000 : node440;
											assign node440 = (inp[2]) ? 3'b010 : 3'b000;
						assign node446 = (inp[4]) ? node472 : node447;
							assign node447 = (inp[8]) ? node457 : node448;
								assign node448 = (inp[5]) ? node454 : node449;
									assign node449 = (inp[10]) ? node451 : 3'b010;
										assign node451 = (inp[1]) ? 3'b100 : 3'b110;
									assign node454 = (inp[10]) ? 3'b000 : 3'b100;
								assign node457 = (inp[10]) ? node465 : node458;
									assign node458 = (inp[5]) ? 3'b010 : node459;
										assign node459 = (inp[1]) ? node461 : 3'b000;
											assign node461 = (inp[11]) ? 3'b010 : 3'b110;
									assign node465 = (inp[1]) ? node467 : 3'b110;
										assign node467 = (inp[5]) ? 3'b100 : node468;
											assign node468 = (inp[11]) ? 3'b100 : 3'b010;
							assign node472 = (inp[10]) ? node500 : node473;
								assign node473 = (inp[8]) ? node483 : node474;
									assign node474 = (inp[2]) ? node476 : 3'b000;
										assign node476 = (inp[5]) ? node480 : node477;
											assign node477 = (inp[11]) ? 3'b000 : 3'b100;
											assign node480 = (inp[11]) ? 3'b100 : 3'b000;
									assign node483 = (inp[1]) ? node493 : node484;
										assign node484 = (inp[5]) ? node488 : node485;
											assign node485 = (inp[11]) ? 3'b010 : 3'b110;
											assign node488 = (inp[11]) ? 3'b000 : node489;
												assign node489 = (inp[2]) ? 3'b100 : 3'b010;
										assign node493 = (inp[5]) ? node495 : 3'b100;
											assign node495 = (inp[2]) ? node497 : 3'b000;
												assign node497 = (inp[11]) ? 3'b000 : 3'b100;
								assign node500 = (inp[11]) ? node512 : node501;
									assign node501 = (inp[8]) ? node507 : node502;
										assign node502 = (inp[2]) ? node504 : 3'b000;
											assign node504 = (inp[5]) ? 3'b100 : 3'b000;
										assign node507 = (inp[5]) ? 3'b000 : node508;
											assign node508 = (inp[1]) ? 3'b000 : 3'b010;
									assign node512 = (inp[1]) ? 3'b000 : node513;
										assign node513 = (inp[8]) ? node515 : 3'b000;
											assign node515 = (inp[5]) ? 3'b000 : 3'b100;
					assign node519 = (inp[8]) ? node521 : 3'b000;
						assign node521 = (inp[0]) ? node537 : node522;
							assign node522 = (inp[5]) ? 3'b000 : node523;
								assign node523 = (inp[10]) ? node529 : node524;
									assign node524 = (inp[1]) ? node526 : 3'b100;
										assign node526 = (inp[4]) ? 3'b000 : 3'b100;
									assign node529 = (inp[1]) ? node531 : 3'b000;
										assign node531 = (inp[4]) ? 3'b100 : node532;
											assign node532 = (inp[11]) ? 3'b000 : 3'b100;
							assign node537 = (inp[4]) ? 3'b000 : node538;
								assign node538 = (inp[10]) ? 3'b000 : node539;
									assign node539 = (inp[5]) ? 3'b000 : node540;
										assign node540 = (inp[11]) ? 3'b000 : 3'b010;
		assign node546 = (inp[3]) ? node952 : node547;
			assign node547 = (inp[0]) ? node665 : node548;
				assign node548 = (inp[7]) ? node558 : node549;
					assign node549 = (inp[5]) ? node551 : 3'b001;
						assign node551 = (inp[8]) ? 3'b001 : node552;
							assign node552 = (inp[10]) ? node554 : 3'b000;
								assign node554 = (inp[9]) ? 3'b000 : 3'b001;
					assign node558 = (inp[5]) ? node620 : node559;
						assign node559 = (inp[9]) ? node569 : node560;
							assign node560 = (inp[11]) ? node562 : 3'b111;
								assign node562 = (inp[10]) ? node564 : 3'b111;
									assign node564 = (inp[8]) ? 3'b111 : node565;
										assign node565 = (inp[1]) ? 3'b011 : 3'b111;
							assign node569 = (inp[4]) ? node591 : node570;
								assign node570 = (inp[10]) ? node578 : node571;
									assign node571 = (inp[8]) ? 3'b111 : node572;
										assign node572 = (inp[11]) ? 3'b111 : node573;
											assign node573 = (inp[2]) ? 3'b011 : 3'b111;
									assign node578 = (inp[11]) ? node586 : node579;
										assign node579 = (inp[8]) ? node583 : node580;
											assign node580 = (inp[1]) ? 3'b011 : 3'b111;
											assign node583 = (inp[1]) ? 3'b111 : 3'b011;
										assign node586 = (inp[8]) ? 3'b011 : node587;
											assign node587 = (inp[1]) ? 3'b011 : 3'b111;
								assign node591 = (inp[1]) ? node607 : node592;
									assign node592 = (inp[10]) ? node600 : node593;
										assign node593 = (inp[8]) ? 3'b111 : node594;
											assign node594 = (inp[2]) ? 3'b011 : node595;
												assign node595 = (inp[11]) ? 3'b011 : 3'b111;
										assign node600 = (inp[8]) ? 3'b011 : node601;
											assign node601 = (inp[11]) ? 3'b101 : node602;
												assign node602 = (inp[2]) ? 3'b111 : 3'b011;
									assign node607 = (inp[10]) ? 3'b101 : node608;
										assign node608 = (inp[11]) ? node614 : node609;
											assign node609 = (inp[2]) ? node611 : 3'b011;
												assign node611 = (inp[8]) ? 3'b011 : 3'b111;
											assign node614 = (inp[8]) ? node616 : 3'b101;
												assign node616 = (inp[2]) ? 3'b001 : 3'b011;
						assign node620 = (inp[8]) ? node622 : 3'b000;
							assign node622 = (inp[9]) ? node630 : node623;
								assign node623 = (inp[10]) ? node625 : 3'b111;
									assign node625 = (inp[1]) ? node627 : 3'b111;
										assign node627 = (inp[11]) ? 3'b011 : 3'b111;
								assign node630 = (inp[4]) ? node644 : node631;
									assign node631 = (inp[11]) ? node639 : node632;
										assign node632 = (inp[2]) ? 3'b011 : node633;
											assign node633 = (inp[1]) ? 3'b111 : node634;
												assign node634 = (inp[10]) ? 3'b111 : 3'b011;
										assign node639 = (inp[10]) ? node641 : 3'b111;
											assign node641 = (inp[1]) ? 3'b011 : 3'b111;
									assign node644 = (inp[11]) ? node658 : node645;
										assign node645 = (inp[10]) ? node653 : node646;
											assign node646 = (inp[1]) ? node650 : node647;
												assign node647 = (inp[2]) ? 3'b011 : 3'b111;
												assign node650 = (inp[2]) ? 3'b111 : 3'b011;
											assign node653 = (inp[1]) ? 3'b101 : node654;
												assign node654 = (inp[2]) ? 3'b111 : 3'b011;
										assign node658 = (inp[10]) ? node662 : node659;
											assign node659 = (inp[1]) ? 3'b101 : 3'b011;
											assign node662 = (inp[1]) ? 3'b001 : 3'b101;
				assign node665 = (inp[10]) ? node831 : node666;
					assign node666 = (inp[4]) ? node730 : node667;
						assign node667 = (inp[5]) ? node695 : node668;
							assign node668 = (inp[11]) ? node682 : node669;
								assign node669 = (inp[8]) ? node677 : node670;
									assign node670 = (inp[7]) ? node672 : 3'b011;
										assign node672 = (inp[9]) ? node674 : 3'b111;
											assign node674 = (inp[1]) ? 3'b101 : 3'b011;
									assign node677 = (inp[1]) ? node679 : 3'b111;
										assign node679 = (inp[7]) ? 3'b011 : 3'b111;
								assign node682 = (inp[7]) ? node684 : 3'b111;
									assign node684 = (inp[9]) ? node688 : node685;
										assign node685 = (inp[1]) ? 3'b011 : 3'b111;
										assign node688 = (inp[1]) ? node692 : node689;
											assign node689 = (inp[8]) ? 3'b111 : 3'b011;
											assign node692 = (inp[8]) ? 3'b111 : 3'b110;
							assign node695 = (inp[8]) ? node711 : node696;
								assign node696 = (inp[7]) ? node704 : node697;
									assign node697 = (inp[9]) ? 3'b101 : node698;
										assign node698 = (inp[1]) ? node700 : 3'b001;
											assign node700 = (inp[11]) ? 3'b001 : 3'b101;
									assign node704 = (inp[9]) ? 3'b111 : node705;
										assign node705 = (inp[1]) ? 3'b011 : node706;
											assign node706 = (inp[11]) ? 3'b111 : 3'b011;
								assign node711 = (inp[11]) ? node721 : node712;
									assign node712 = (inp[7]) ? node714 : 3'b011;
										assign node714 = (inp[1]) ? node718 : node715;
											assign node715 = (inp[9]) ? 3'b011 : 3'b111;
											assign node718 = (inp[9]) ? 3'b101 : 3'b111;
									assign node721 = (inp[7]) ? node723 : 3'b111;
										assign node723 = (inp[1]) ? node727 : node724;
											assign node724 = (inp[9]) ? 3'b011 : 3'b111;
											assign node727 = (inp[9]) ? 3'b110 : 3'b011;
						assign node730 = (inp[11]) ? node786 : node731;
							assign node731 = (inp[7]) ? node749 : node732;
								assign node732 = (inp[8]) ? node746 : node733;
									assign node733 = (inp[5]) ? node735 : 3'b001;
										assign node735 = (inp[2]) ? node741 : node736;
											assign node736 = (inp[1]) ? 3'b100 : node737;
												assign node737 = (inp[9]) ? 3'b100 : 3'b000;
											assign node741 = (inp[9]) ? 3'b110 : node742;
												assign node742 = (inp[1]) ? 3'b110 : 3'b010;
									assign node746 = (inp[5]) ? 3'b001 : 3'b101;
								assign node749 = (inp[9]) ? node767 : node750;
									assign node750 = (inp[1]) ? node758 : node751;
										assign node751 = (inp[8]) ? 3'b111 : node752;
											assign node752 = (inp[5]) ? node754 : 3'b111;
												assign node754 = (inp[2]) ? 3'b001 : 3'b011;
										assign node758 = (inp[5]) ? node762 : node759;
											assign node759 = (inp[8]) ? 3'b011 : 3'b101;
											assign node762 = (inp[8]) ? 3'b101 : node763;
												assign node763 = (inp[2]) ? 3'b101 : 3'b111;
									assign node767 = (inp[8]) ? node777 : node768;
										assign node768 = (inp[5]) ? node774 : node769;
											assign node769 = (inp[2]) ? 3'b001 : node770;
												assign node770 = (inp[1]) ? 3'b001 : 3'b101;
											assign node774 = (inp[2]) ? 3'b101 : 3'b111;
										assign node777 = (inp[1]) ? 3'b001 : node778;
											assign node778 = (inp[5]) ? node782 : node779;
												assign node779 = (inp[2]) ? 3'b101 : 3'b011;
												assign node782 = (inp[2]) ? 3'b001 : 3'b101;
							assign node786 = (inp[7]) ? node798 : node787;
								assign node787 = (inp[5]) ? node791 : node788;
									assign node788 = (inp[8]) ? 3'b111 : 3'b011;
									assign node791 = (inp[8]) ? 3'b011 : node792;
										assign node792 = (inp[9]) ? 3'b110 : node793;
											assign node793 = (inp[1]) ? 3'b110 : 3'b010;
								assign node798 = (inp[9]) ? node816 : node799;
									assign node799 = (inp[5]) ? node807 : node800;
										assign node800 = (inp[1]) ? node804 : node801;
											assign node801 = (inp[8]) ? 3'b111 : 3'b011;
											assign node804 = (inp[8]) ? 3'b011 : 3'b101;
										assign node807 = (inp[8]) ? node813 : node808;
											assign node808 = (inp[2]) ? node810 : 3'b101;
												assign node810 = (inp[1]) ? 3'b001 : 3'b101;
											assign node813 = (inp[1]) ? 3'b101 : 3'b011;
									assign node816 = (inp[1]) ? node822 : node817;
										assign node817 = (inp[8]) ? node819 : 3'b101;
											assign node819 = (inp[5]) ? 3'b001 : 3'b101;
										assign node822 = (inp[5]) ? node828 : node823;
											assign node823 = (inp[8]) ? node825 : 3'b110;
												assign node825 = (inp[2]) ? 3'b000 : 3'b001;
											assign node828 = (inp[8]) ? 3'b110 : 3'b101;
					assign node831 = (inp[7]) ? node861 : node832;
						assign node832 = (inp[11]) ? node844 : node833;
							assign node833 = (inp[5]) ? node835 : 3'b110;
								assign node835 = (inp[8]) ? 3'b110 : node836;
									assign node836 = (inp[4]) ? 3'b110 : node837;
										assign node837 = (inp[1]) ? node839 : 3'b100;
											assign node839 = (inp[9]) ? 3'b100 : 3'b000;
							assign node844 = (inp[4]) ? node856 : node845;
								assign node845 = (inp[5]) ? node849 : node846;
									assign node846 = (inp[8]) ? 3'b110 : 3'b010;
									assign node849 = (inp[8]) ? 3'b010 : node850;
										assign node850 = (inp[1]) ? node852 : 3'b100;
											assign node852 = (inp[9]) ? 3'b100 : 3'b000;
								assign node856 = (inp[5]) ? node858 : 3'b100;
									assign node858 = (inp[8]) ? 3'b100 : 3'b110;
						assign node861 = (inp[8]) ? node907 : node862;
							assign node862 = (inp[5]) ? node892 : node863;
								assign node863 = (inp[9]) ? node879 : node864;
									assign node864 = (inp[11]) ? node872 : node865;
										assign node865 = (inp[1]) ? node869 : node866;
											assign node866 = (inp[4]) ? 3'b011 : 3'b111;
											assign node869 = (inp[4]) ? 3'b001 : 3'b011;
										assign node872 = (inp[1]) ? node876 : node873;
											assign node873 = (inp[4]) ? 3'b101 : 3'b111;
											assign node876 = (inp[4]) ? 3'b001 : 3'b101;
									assign node879 = (inp[1]) ? node887 : node880;
										assign node880 = (inp[11]) ? node884 : node881;
											assign node881 = (inp[4]) ? 3'b001 : 3'b101;
											assign node884 = (inp[4]) ? 3'b110 : 3'b101;
										assign node887 = (inp[11]) ? node889 : 3'b110;
											assign node889 = (inp[2]) ? 3'b010 : 3'b110;
								assign node892 = (inp[4]) ? node898 : node893;
									assign node893 = (inp[9]) ? 3'b110 : node894;
										assign node894 = (inp[1]) ? 3'b010 : 3'b110;
									assign node898 = (inp[9]) ? 3'b100 : node899;
										assign node899 = (inp[1]) ? node901 : 3'b100;
											assign node901 = (inp[11]) ? node903 : 3'b000;
												assign node903 = (inp[2]) ? 3'b100 : 3'b000;
							assign node907 = (inp[9]) ? node927 : node908;
								assign node908 = (inp[1]) ? node918 : node909;
									assign node909 = (inp[4]) ? node911 : 3'b111;
										assign node911 = (inp[11]) ? node915 : node912;
											assign node912 = (inp[5]) ? 3'b011 : 3'b111;
											assign node915 = (inp[5]) ? 3'b101 : 3'b011;
									assign node918 = (inp[5]) ? node920 : 3'b101;
										assign node920 = (inp[11]) ? node924 : node921;
											assign node921 = (inp[4]) ? 3'b001 : 3'b011;
											assign node924 = (inp[4]) ? 3'b001 : 3'b101;
								assign node927 = (inp[1]) ? node939 : node928;
									assign node928 = (inp[5]) ? node934 : node929;
										assign node929 = (inp[4]) ? node931 : 3'b011;
											assign node931 = (inp[11]) ? 3'b001 : 3'b101;
										assign node934 = (inp[4]) ? node936 : 3'b101;
											assign node936 = (inp[11]) ? 3'b110 : 3'b001;
									assign node939 = (inp[5]) ? node947 : node940;
										assign node940 = (inp[4]) ? node944 : node941;
											assign node941 = (inp[11]) ? 3'b001 : 3'b101;
											assign node944 = (inp[11]) ? 3'b110 : 3'b100;
										assign node947 = (inp[11]) ? node949 : 3'b110;
											assign node949 = (inp[4]) ? 3'b010 : 3'b110;
			assign node952 = (inp[7]) ? node1220 : node953;
				assign node953 = (inp[0]) ? node1095 : node954;
					assign node954 = (inp[10]) ? node1068 : node955;
						assign node955 = (inp[11]) ? node1001 : node956;
							assign node956 = (inp[2]) ? node990 : node957;
								assign node957 = (inp[1]) ? node973 : node958;
									assign node958 = (inp[9]) ? node966 : node959;
										assign node959 = (inp[5]) ? node963 : node960;
											assign node960 = (inp[8]) ? 3'b000 : 3'b110;
											assign node963 = (inp[8]) ? 3'b110 : 3'b000;
										assign node966 = (inp[5]) ? node970 : node967;
											assign node967 = (inp[8]) ? 3'b000 : 3'b110;
											assign node970 = (inp[8]) ? 3'b110 : 3'b000;
									assign node973 = (inp[9]) ? node983 : node974;
										assign node974 = (inp[8]) ? node980 : node975;
											assign node975 = (inp[5]) ? node977 : 3'b110;
												assign node977 = (inp[4]) ? 3'b000 : 3'b010;
											assign node980 = (inp[5]) ? 3'b110 : 3'b000;
										assign node983 = (inp[8]) ? node987 : node984;
											assign node984 = (inp[5]) ? 3'b000 : 3'b110;
											assign node987 = (inp[5]) ? 3'b110 : 3'b000;
								assign node990 = (inp[5]) ? node994 : node991;
									assign node991 = (inp[8]) ? 3'b000 : 3'b110;
									assign node994 = (inp[8]) ? 3'b110 : node995;
										assign node995 = (inp[1]) ? node997 : 3'b000;
											assign node997 = (inp[9]) ? 3'b000 : 3'b010;
							assign node1001 = (inp[4]) ? node1031 : node1002;
								assign node1002 = (inp[2]) ? node1016 : node1003;
									assign node1003 = (inp[1]) ? node1009 : node1004;
										assign node1004 = (inp[8]) ? 3'b000 : node1005;
											assign node1005 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1009 = (inp[8]) ? node1013 : node1010;
											assign node1010 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1013 = (inp[5]) ? 3'b010 : 3'b000;
									assign node1016 = (inp[9]) ? node1024 : node1017;
										assign node1017 = (inp[5]) ? node1021 : node1018;
											assign node1018 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1021 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1024 = (inp[8]) ? node1028 : node1025;
											assign node1025 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1028 = (inp[5]) ? 3'b010 : 3'b000;
								assign node1031 = (inp[1]) ? node1055 : node1032;
									assign node1032 = (inp[9]) ? node1048 : node1033;
										assign node1033 = (inp[2]) ? node1041 : node1034;
											assign node1034 = (inp[8]) ? node1038 : node1035;
												assign node1035 = (inp[5]) ? 3'b000 : 3'b010;
												assign node1038 = (inp[5]) ? 3'b010 : 3'b000;
											assign node1041 = (inp[8]) ? node1045 : node1042;
												assign node1042 = (inp[5]) ? 3'b000 : 3'b010;
												assign node1045 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1048 = (inp[5]) ? node1052 : node1049;
											assign node1049 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1052 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1055 = (inp[9]) ? node1061 : node1056;
										assign node1056 = (inp[8]) ? node1058 : 3'b010;
											assign node1058 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1061 = (inp[8]) ? node1065 : node1062;
											assign node1062 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1065 = (inp[5]) ? 3'b010 : 3'b000;
						assign node1068 = (inp[11]) ? node1084 : node1069;
							assign node1069 = (inp[8]) ? node1081 : node1070;
								assign node1070 = (inp[5]) ? node1072 : 3'b010;
									assign node1072 = (inp[9]) ? 3'b100 : node1073;
										assign node1073 = (inp[1]) ? node1075 : 3'b110;
											assign node1075 = (inp[2]) ? 3'b100 : node1076;
												assign node1076 = (inp[4]) ? 3'b110 : 3'b100;
								assign node1081 = (inp[5]) ? 3'b010 : 3'b000;
							assign node1084 = (inp[5]) ? node1088 : node1085;
								assign node1085 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1088 = (inp[9]) ? 3'b100 : node1089;
									assign node1089 = (inp[8]) ? 3'b100 : node1090;
										assign node1090 = (inp[1]) ? 3'b100 : 3'b110;
					assign node1095 = (inp[9]) ? node1193 : node1096;
						assign node1096 = (inp[10]) ? node1160 : node1097;
							assign node1097 = (inp[4]) ? node1121 : node1098;
								assign node1098 = (inp[11]) ? node1112 : node1099;
									assign node1099 = (inp[5]) ? node1105 : node1100;
										assign node1100 = (inp[8]) ? 3'b100 : node1101;
											assign node1101 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1105 = (inp[1]) ? node1109 : node1106;
											assign node1106 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1109 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1112 = (inp[8]) ? node1116 : node1113;
										assign node1113 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1116 = (inp[5]) ? 3'b010 : node1117;
											assign node1117 = (inp[1]) ? 3'b110 : 3'b100;
								assign node1121 = (inp[2]) ? node1141 : node1122;
									assign node1122 = (inp[5]) ? node1132 : node1123;
										assign node1123 = (inp[8]) ? node1127 : node1124;
											assign node1124 = (inp[1]) ? 3'b000 : 3'b010;
											assign node1127 = (inp[11]) ? 3'b000 : node1128;
												assign node1128 = (inp[1]) ? 3'b010 : 3'b000;
										assign node1132 = (inp[1]) ? node1136 : node1133;
											assign node1133 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1136 = (inp[11]) ? node1138 : 3'b000;
												assign node1138 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1141 = (inp[1]) ? node1151 : node1142;
										assign node1142 = (inp[5]) ? node1148 : node1143;
											assign node1143 = (inp[8]) ? node1145 : 3'b010;
												assign node1145 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1148 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1151 = (inp[5]) ? node1157 : node1152;
											assign node1152 = (inp[11]) ? 3'b100 : node1153;
												assign node1153 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1157 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1160 = (inp[1]) ? node1168 : node1161;
								assign node1161 = (inp[8]) ? node1165 : node1162;
									assign node1162 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1165 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1168 = (inp[4]) ? node1180 : node1169;
									assign node1169 = (inp[8]) ? node1175 : node1170;
										assign node1170 = (inp[5]) ? 3'b100 : node1171;
											assign node1171 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1175 = (inp[11]) ? node1177 : 3'b010;
											assign node1177 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1180 = (inp[11]) ? 3'b000 : node1181;
										assign node1181 = (inp[5]) ? node1187 : node1182;
											assign node1182 = (inp[2]) ? node1184 : 3'b100;
												assign node1184 = (inp[8]) ? 3'b100 : 3'b000;
											assign node1187 = (inp[8]) ? node1189 : 3'b000;
												assign node1189 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1193 = (inp[5]) ? node1211 : node1194;
							assign node1194 = (inp[8]) ? node1196 : 3'b000;
								assign node1196 = (inp[10]) ? node1204 : node1197;
									assign node1197 = (inp[4]) ? node1199 : 3'b100;
										assign node1199 = (inp[11]) ? node1201 : 3'b000;
											assign node1201 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1204 = (inp[4]) ? node1206 : 3'b000;
										assign node1206 = (inp[2]) ? node1208 : 3'b000;
											assign node1208 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1211 = (inp[4]) ? 3'b000 : node1212;
								assign node1212 = (inp[10]) ? 3'b000 : node1213;
									assign node1213 = (inp[8]) ? 3'b000 : node1214;
										assign node1214 = (inp[11]) ? 3'b000 : 3'b010;
				assign node1220 = (inp[0]) ? node1418 : node1221;
					assign node1221 = (inp[9]) ? node1321 : node1222;
						assign node1222 = (inp[4]) ? node1264 : node1223;
							assign node1223 = (inp[1]) ? node1241 : node1224;
								assign node1224 = (inp[8]) ? node1234 : node1225;
									assign node1225 = (inp[5]) ? node1229 : node1226;
										assign node1226 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1229 = (inp[10]) ? 3'b110 : node1230;
											assign node1230 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1234 = (inp[10]) ? node1236 : 3'b111;
										assign node1236 = (inp[5]) ? 3'b011 : node1237;
											assign node1237 = (inp[11]) ? 3'b011 : 3'b111;
								assign node1241 = (inp[10]) ? node1255 : node1242;
									assign node1242 = (inp[8]) ? node1250 : node1243;
										assign node1243 = (inp[11]) ? node1247 : node1244;
											assign node1244 = (inp[5]) ? 3'b001 : 3'b011;
											assign node1247 = (inp[5]) ? 3'b111 : 3'b011;
										assign node1250 = (inp[5]) ? 3'b011 : node1251;
											assign node1251 = (inp[11]) ? 3'b011 : 3'b111;
									assign node1255 = (inp[5]) ? node1261 : node1256;
										assign node1256 = (inp[8]) ? node1258 : 3'b101;
											assign node1258 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1261 = (inp[8]) ? 3'b101 : 3'b111;
							assign node1264 = (inp[10]) ? node1294 : node1265;
								assign node1265 = (inp[8]) ? node1281 : node1266;
									assign node1266 = (inp[5]) ? node1276 : node1267;
										assign node1267 = (inp[1]) ? node1271 : node1268;
											assign node1268 = (inp[2]) ? 3'b101 : 3'b011;
											assign node1271 = (inp[11]) ? 3'b001 : node1272;
												assign node1272 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1276 = (inp[11]) ? 3'b110 : node1277;
											assign node1277 = (inp[1]) ? 3'b001 : 3'b000;
									assign node1281 = (inp[5]) ? node1287 : node1282;
										assign node1282 = (inp[11]) ? node1284 : 3'b011;
											assign node1284 = (inp[1]) ? 3'b111 : 3'b001;
										assign node1287 = (inp[1]) ? 3'b001 : node1288;
											assign node1288 = (inp[11]) ? 3'b101 : node1289;
												assign node1289 = (inp[2]) ? 3'b101 : 3'b011;
								assign node1294 = (inp[8]) ? node1306 : node1295;
									assign node1295 = (inp[5]) ? 3'b110 : node1296;
										assign node1296 = (inp[1]) ? node1300 : node1297;
											assign node1297 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1300 = (inp[11]) ? 3'b110 : node1301;
												assign node1301 = (inp[2]) ? 3'b110 : 3'b001;
									assign node1306 = (inp[1]) ? node1312 : node1307;
										assign node1307 = (inp[11]) ? node1309 : 3'b101;
											assign node1309 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1312 = (inp[5]) ? node1316 : node1313;
											assign node1313 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1316 = (inp[11]) ? 3'b110 : node1317;
												assign node1317 = (inp[2]) ? 3'b110 : 3'b001;
						assign node1321 = (inp[4]) ? node1357 : node1322;
							assign node1322 = (inp[8]) ? node1336 : node1323;
								assign node1323 = (inp[5]) ? node1331 : node1324;
									assign node1324 = (inp[1]) ? node1328 : node1325;
										assign node1325 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1328 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1331 = (inp[10]) ? 3'b110 : node1332;
										assign node1332 = (inp[11]) ? 3'b110 : 3'b000;
								assign node1336 = (inp[10]) ? node1348 : node1337;
									assign node1337 = (inp[1]) ? node1343 : node1338;
										assign node1338 = (inp[11]) ? 3'b101 : node1339;
											assign node1339 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1343 = (inp[5]) ? 3'b001 : node1344;
											assign node1344 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1348 = (inp[1]) ? node1354 : node1349;
										assign node1349 = (inp[5]) ? 3'b001 : node1350;
											assign node1350 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1354 = (inp[5]) ? 3'b110 : 3'b001;
							assign node1357 = (inp[10]) ? node1389 : node1358;
								assign node1358 = (inp[11]) ? node1374 : node1359;
									assign node1359 = (inp[8]) ? node1363 : node1360;
										assign node1360 = (inp[5]) ? 3'b000 : 3'b110;
										assign node1363 = (inp[5]) ? node1367 : node1364;
											assign node1364 = (inp[2]) ? 3'b101 : 3'b001;
											assign node1367 = (inp[1]) ? node1371 : node1368;
												assign node1368 = (inp[2]) ? 3'b110 : 3'b001;
												assign node1371 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1374 = (inp[5]) ? node1384 : node1375;
										assign node1375 = (inp[1]) ? node1381 : node1376;
											assign node1376 = (inp[8]) ? node1378 : 3'b110;
												assign node1378 = (inp[2]) ? 3'b000 : 3'b001;
											assign node1381 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1384 = (inp[8]) ? node1386 : 3'b110;
											assign node1386 = (inp[1]) ? 3'b010 : 3'b110;
								assign node1389 = (inp[11]) ? node1403 : node1390;
									assign node1390 = (inp[1]) ? node1392 : 3'b110;
										assign node1392 = (inp[5]) ? node1398 : node1393;
											assign node1393 = (inp[2]) ? node1395 : 3'b010;
												assign node1395 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1398 = (inp[2]) ? 3'b110 : node1399;
												assign node1399 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1403 = (inp[1]) ? node1411 : node1404;
										assign node1404 = (inp[8]) ? node1408 : node1405;
											assign node1405 = (inp[5]) ? 3'b110 : 3'b010;
											assign node1408 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1411 = (inp[5]) ? node1415 : node1412;
											assign node1412 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1415 = (inp[8]) ? 3'b100 : 3'b110;
					assign node1418 = (inp[9]) ? node1526 : node1419;
						assign node1419 = (inp[4]) ? node1455 : node1420;
							assign node1420 = (inp[5]) ? node1440 : node1421;
								assign node1421 = (inp[10]) ? node1431 : node1422;
									assign node1422 = (inp[1]) ? node1426 : node1423;
										assign node1423 = (inp[8]) ? 3'b011 : 3'b101;
										assign node1426 = (inp[8]) ? node1428 : 3'b001;
											assign node1428 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1431 = (inp[1]) ? node1435 : node1432;
										assign node1432 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1435 = (inp[11]) ? 3'b110 : node1436;
											assign node1436 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1440 = (inp[8]) ? node1448 : node1441;
									assign node1441 = (inp[1]) ? 3'b110 : node1442;
										assign node1442 = (inp[11]) ? 3'b010 : node1443;
											assign node1443 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1448 = (inp[10]) ? node1452 : node1449;
										assign node1449 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1452 = (inp[1]) ? 3'b110 : 3'b001;
							assign node1455 = (inp[10]) ? node1491 : node1456;
								assign node1456 = (inp[1]) ? node1474 : node1457;
									assign node1457 = (inp[8]) ? node1463 : node1458;
										assign node1458 = (inp[11]) ? node1460 : 3'b110;
											assign node1460 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1463 = (inp[5]) ? node1469 : node1464;
											assign node1464 = (inp[11]) ? 3'b001 : node1465;
												assign node1465 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1469 = (inp[2]) ? 3'b110 : node1470;
												assign node1470 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1474 = (inp[8]) ? node1484 : node1475;
										assign node1475 = (inp[11]) ? node1479 : node1476;
											assign node1476 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1479 = (inp[5]) ? node1481 : 3'b010;
												assign node1481 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1484 = (inp[5]) ? node1486 : 3'b110;
											assign node1486 = (inp[2]) ? node1488 : 3'b110;
												assign node1488 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1491 = (inp[1]) ? node1509 : node1492;
									assign node1492 = (inp[5]) ? node1502 : node1493;
										assign node1493 = (inp[11]) ? node1499 : node1494;
											assign node1494 = (inp[8]) ? 3'b001 : node1495;
												assign node1495 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1499 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1502 = (inp[8]) ? node1504 : 3'b010;
											assign node1504 = (inp[2]) ? 3'b010 : node1505;
												assign node1505 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1509 = (inp[5]) ? node1517 : node1510;
										assign node1510 = (inp[8]) ? 3'b010 : node1511;
											assign node1511 = (inp[2]) ? 3'b010 : node1512;
												assign node1512 = (inp[11]) ? 3'b100 : 3'b110;
										assign node1517 = (inp[8]) ? node1523 : node1518;
											assign node1518 = (inp[11]) ? node1520 : 3'b100;
												assign node1520 = (inp[2]) ? 3'b000 : 3'b100;
											assign node1523 = (inp[11]) ? 3'b100 : 3'b010;
						assign node1526 = (inp[4]) ? node1556 : node1527;
							assign node1527 = (inp[5]) ? node1547 : node1528;
								assign node1528 = (inp[10]) ? node1538 : node1529;
									assign node1529 = (inp[8]) ? node1533 : node1530;
										assign node1530 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1533 = (inp[1]) ? node1535 : 3'b001;
											assign node1535 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1538 = (inp[1]) ? node1542 : node1539;
										assign node1539 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1542 = (inp[8]) ? node1544 : 3'b100;
											assign node1544 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1547 = (inp[8]) ? node1549 : 3'b000;
									assign node1549 = (inp[10]) ? node1553 : node1550;
										assign node1550 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1553 = (inp[1]) ? 3'b100 : 3'b010;
							assign node1556 = (inp[1]) ? node1584 : node1557;
								assign node1557 = (inp[8]) ? node1565 : node1558;
									assign node1558 = (inp[5]) ? 3'b000 : node1559;
										assign node1559 = (inp[11]) ? node1561 : 3'b100;
											assign node1561 = (inp[10]) ? 3'b000 : 3'b100;
									assign node1565 = (inp[5]) ? node1579 : node1566;
										assign node1566 = (inp[10]) ? node1574 : node1567;
											assign node1567 = (inp[11]) ? node1571 : node1568;
												assign node1568 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1571 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1574 = (inp[11]) ? 3'b100 : node1575;
												assign node1575 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1579 = (inp[10]) ? node1581 : 3'b100;
											assign node1581 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1584 = (inp[10]) ? 3'b000 : node1585;
									assign node1585 = (inp[8]) ? node1593 : node1586;
										assign node1586 = (inp[2]) ? node1588 : 3'b000;
											assign node1588 = (inp[11]) ? 3'b000 : node1589;
												assign node1589 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1593 = (inp[5]) ? node1595 : 3'b100;
											assign node1595 = (inp[11]) ? 3'b000 : 3'b100;

endmodule