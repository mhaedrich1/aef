module dtc_split05_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;

	assign outp = (inp[2]) ? node52 : node1;
		assign node1 = (inp[3]) ? node29 : node2;
			assign node2 = (inp[10]) ? node14 : node3;
				assign node3 = (inp[5]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node6 : 3'b111;
						assign node6 = (inp[6]) ? node8 : 3'b110;
							assign node8 = (inp[11]) ? node10 : 3'b110;
								assign node10 = (inp[8]) ? 3'b111 : 3'b110;
				assign node14 = (inp[9]) ? node22 : node15;
					assign node15 = (inp[11]) ? 3'b110 : node16;
						assign node16 = (inp[1]) ? node18 : 3'b110;
							assign node18 = (inp[7]) ? 3'b110 : 3'b111;
					assign node22 = (inp[5]) ? node24 : 3'b110;
						assign node24 = (inp[4]) ? 3'b011 : node25;
							assign node25 = (inp[0]) ? 3'b111 : 3'b110;
			assign node29 = (inp[4]) ? node45 : node30;
				assign node30 = (inp[10]) ? node40 : node31;
					assign node31 = (inp[0]) ? 3'b111 : node32;
						assign node32 = (inp[6]) ? 3'b111 : node33;
							assign node33 = (inp[11]) ? 3'b111 : node34;
								assign node34 = (inp[1]) ? 3'b111 : 3'b110;
					assign node40 = (inp[5]) ? node42 : 3'b110;
						assign node42 = (inp[11]) ? 3'b011 : 3'b110;
				assign node45 = (inp[5]) ? 3'b010 : node46;
					assign node46 = (inp[0]) ? 3'b011 : node47;
						assign node47 = (inp[1]) ? 3'b011 : 3'b010;
		assign node52 = (inp[4]) ? node82 : node53;
			assign node53 = (inp[3]) ? node71 : node54;
				assign node54 = (inp[10]) ? node62 : node55;
					assign node55 = (inp[5]) ? node57 : 3'b011;
						assign node57 = (inp[9]) ? 3'b010 : node58;
							assign node58 = (inp[6]) ? 3'b010 : 3'b011;
					assign node62 = (inp[5]) ? 3'b011 : node63;
						assign node63 = (inp[9]) ? node65 : 3'b010;
							assign node65 = (inp[7]) ? node67 : 3'b010;
								assign node67 = (inp[0]) ? 3'b011 : 3'b010;
				assign node71 = (inp[10]) ? node77 : node72;
					assign node72 = (inp[5]) ? 3'b010 : node73;
						assign node73 = (inp[9]) ? 3'b010 : 3'b011;
					assign node77 = (inp[8]) ? node79 : 3'b111;
						assign node79 = (inp[9]) ? 3'b110 : 3'b111;
			assign node82 = (inp[3]) ? node100 : node83;
				assign node83 = (inp[5]) ? node93 : node84;
					assign node84 = (inp[11]) ? node86 : 3'b101;
						assign node86 = (inp[9]) ? node88 : 3'b101;
							assign node88 = (inp[7]) ? 3'b100 : node89;
								assign node89 = (inp[1]) ? 3'b101 : 3'b100;
					assign node93 = (inp[9]) ? node95 : 3'b100;
						assign node95 = (inp[10]) ? 3'b001 : node96;
							assign node96 = (inp[8]) ? 3'b101 : 3'b100;
				assign node100 = (inp[5]) ? node106 : node101;
					assign node101 = (inp[10]) ? node103 : 3'b000;
						assign node103 = (inp[9]) ? 3'b100 : 3'b101;
					assign node106 = (inp[9]) ? node108 : 3'b001;
						assign node108 = (inp[11]) ? 3'b000 : node109;
							assign node109 = (inp[7]) ? node111 : 3'b001;
								assign node111 = (inp[6]) ? 3'b001 : 3'b000;

endmodule