module dtc_split75_bm28 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node7;
	wire [10-1:0] node10;
	wire [10-1:0] node11;
	wire [10-1:0] node15;
	wire [10-1:0] node16;
	wire [10-1:0] node18;
	wire [10-1:0] node21;
	wire [10-1:0] node22;
	wire [10-1:0] node25;
	wire [10-1:0] node28;
	wire [10-1:0] node29;
	wire [10-1:0] node30;
	wire [10-1:0] node33;
	wire [10-1:0] node34;
	wire [10-1:0] node37;
	wire [10-1:0] node40;
	wire [10-1:0] node41;
	wire [10-1:0] node44;
	wire [10-1:0] node46;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node52;
	wire [10-1:0] node55;
	wire [10-1:0] node58;
	wire [10-1:0] node59;
	wire [10-1:0] node61;
	wire [10-1:0] node64;
	wire [10-1:0] node67;
	wire [10-1:0] node68;
	wire [10-1:0] node69;
	wire [10-1:0] node72;
	wire [10-1:0] node73;
	wire [10-1:0] node76;
	wire [10-1:0] node79;
	wire [10-1:0] node80;
	wire [10-1:0] node81;
	wire [10-1:0] node84;
	wire [10-1:0] node87;
	wire [10-1:0] node88;
	wire [10-1:0] node91;
	wire [10-1:0] node94;
	wire [10-1:0] node95;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node99;
	wire [10-1:0] node103;
	wire [10-1:0] node104;
	wire [10-1:0] node107;
	wire [10-1:0] node110;
	wire [10-1:0] node111;
	wire [10-1:0] node113;
	wire [10-1:0] node116;
	wire [10-1:0] node119;
	wire [10-1:0] node120;
	wire [10-1:0] node121;
	wire [10-1:0] node123;
	wire [10-1:0] node126;
	wire [10-1:0] node127;
	wire [10-1:0] node130;
	wire [10-1:0] node133;
	wire [10-1:0] node134;
	wire [10-1:0] node135;
	wire [10-1:0] node138;
	wire [10-1:0] node141;
	wire [10-1:0] node143;
	wire [10-1:0] node146;
	wire [10-1:0] node147;
	wire [10-1:0] node148;
	wire [10-1:0] node149;
	wire [10-1:0] node150;
	wire [10-1:0] node154;
	wire [10-1:0] node157;
	wire [10-1:0] node158;
	wire [10-1:0] node159;
	wire [10-1:0] node163;
	wire [10-1:0] node166;
	wire [10-1:0] node167;
	wire [10-1:0] node168;
	wire [10-1:0] node169;
	wire [10-1:0] node173;
	wire [10-1:0] node174;
	wire [10-1:0] node177;
	wire [10-1:0] node180;
	wire [10-1:0] node181;
	wire [10-1:0] node183;
	wire [10-1:0] node186;
	wire [10-1:0] node188;

	assign outp = (inp[4]) ? node94 : node1;
		assign node1 = (inp[2]) ? node49 : node2;
			assign node2 = (inp[5]) ? node28 : node3;
				assign node3 = (inp[3]) ? node15 : node4;
					assign node4 = (inp[6]) ? node10 : node5;
						assign node5 = (inp[1]) ? node7 : 10'b0101011001;
							assign node7 = (inp[0]) ? 10'b0011110001 : 10'b0001010101;
						assign node10 = (inp[1]) ? 10'b0111010000 : node11;
							assign node11 = (inp[0]) ? 10'b0011011000 : 10'b0111111000;
					assign node15 = (inp[1]) ? node21 : node16;
						assign node16 = (inp[6]) ? node18 : 10'b0001100101;
							assign node18 = (inp[0]) ? 10'b0011000000 : 10'b0111100000;
						assign node21 = (inp[6]) ? node25 : node22;
							assign node22 = (inp[0]) ? 10'b0011101000 : 10'b0001001100;
							assign node25 = (inp[0]) ? 10'b0001001001 : 10'b0101101001;
				assign node28 = (inp[3]) ? node40 : node29;
					assign node29 = (inp[6]) ? node33 : node30;
						assign node30 = (inp[0]) ? 10'b0010110000 : 10'b0000010100;
						assign node33 = (inp[1]) ? node37 : node34;
							assign node34 = (inp[0]) ? 10'b0000111001 : 10'b0110011001;
							assign node37 = (inp[0]) ? 10'b0000010001 : 10'b0100110001;
					assign node40 = (inp[1]) ? node44 : node41;
						assign node41 = (inp[6]) ? 10'b0110000001 : 10'b0100000000;
						assign node44 = (inp[6]) ? node46 : 10'b0010001001;
							assign node46 = (inp[0]) ? 10'b0000001000 : 10'b0100101000;
			assign node49 = (inp[3]) ? node67 : node50;
				assign node50 = (inp[5]) ? node58 : node51;
					assign node51 = (inp[6]) ? node55 : node52;
						assign node52 = (inp[1]) ? 10'b1000000101 : 10'b1000101101;
						assign node55 = (inp[0]) ? 10'b1010001000 : 10'b1110101000;
					assign node58 = (inp[1]) ? node64 : node59;
						assign node59 = (inp[0]) ? node61 : 10'b1111000001;
							assign node61 = (inp[6]) ? 10'b1001100001 : 10'b1101000000;
						assign node64 = (inp[0]) ? 10'b1001001000 : 10'b1101101000;
				assign node67 = (inp[5]) ? node79 : node68;
					assign node68 = (inp[1]) ? node72 : node69;
						assign node69 = (inp[6]) ? 10'b1111011001 : 10'b1101011000;
						assign node72 = (inp[6]) ? node76 : node73;
							assign node73 = (inp[0]) ? 10'b1011110000 : 10'b1001010100;
							assign node76 = (inp[0]) ? 10'b1001010001 : 10'b1101110001;
					assign node79 = (inp[6]) ? node87 : node80;
						assign node80 = (inp[1]) ? node84 : node81;
							assign node81 = (inp[0]) ? 10'b1010111001 : 10'b1000011101;
							assign node84 = (inp[0]) ? 10'b1010010001 : 10'b1110110001;
						assign node87 = (inp[1]) ? node91 : node88;
							assign node88 = (inp[0]) ? 10'b1000111000 : 10'b1110011000;
							assign node91 = (inp[0]) ? 10'b1000010000 : 10'b1100110000;
		assign node94 = (inp[3]) ? node146 : node95;
			assign node95 = (inp[2]) ? node119 : node96;
				assign node96 = (inp[5]) ? node110 : node97;
					assign node97 = (inp[6]) ? node103 : node98;
						assign node98 = (inp[1]) ? 10'b1010110011 : node99;
							assign node99 = (inp[0]) ? 10'b1100011011 : 10'b1000111111;
						assign node103 = (inp[1]) ? node107 : node104;
							assign node104 = (inp[0]) ? 10'b1010011010 : 10'b1110111010;
							assign node107 = (inp[0]) ? 10'b1000110010 : 10'b1110010010;
					assign node110 = (inp[0]) ? node116 : node111;
						assign node111 = (inp[1]) ? node113 : 10'b1111010011;
							assign node113 = (inp[6]) ? 10'b1101111010 : 10'b1111111011;
						assign node116 = (inp[6]) ? 10'b1001011010 : 10'b1011011011;
				assign node119 = (inp[5]) ? node133 : node120;
					assign node120 = (inp[1]) ? node126 : node121;
						assign node121 = (inp[6]) ? node123 : 10'b0001110111;
							assign node123 = (inp[0]) ? 10'b0011010010 : 10'b0111110010;
						assign node126 = (inp[6]) ? node130 : node127;
							assign node127 = (inp[0]) ? 10'b0011111010 : 10'b0001011110;
							assign node130 = (inp[0]) ? 10'b0001011011 : 10'b0101111011;
					assign node133 = (inp[1]) ? node141 : node134;
						assign node134 = (inp[6]) ? node138 : node135;
							assign node135 = (inp[0]) ? 10'b0100010010 : 10'b0000110110;
							assign node138 = (inp[0]) ? 10'b0000110011 : 10'b0110010011;
						assign node141 = (inp[0]) ? node143 : 10'b0100111010;
							assign node143 = (inp[6]) ? 10'b0000011010 : 10'b0010011011;
			assign node146 = (inp[2]) ? node166 : node147;
				assign node147 = (inp[5]) ? node157 : node148;
					assign node148 = (inp[6]) ? node154 : node149;
						assign node149 = (inp[1]) ? 10'b1000001110 : node150;
							assign node150 = (inp[0]) ? 10'b1100000011 : 10'b1000100111;
						assign node154 = (inp[1]) ? 10'b1100101011 : 10'b1110100010;
					assign node157 = (inp[6]) ? node163 : node158;
						assign node158 = (inp[1]) ? 10'b1111100011 : node159;
							assign node159 = (inp[0]) ? 10'b1011101011 : 10'b1001001111;
						assign node163 = (inp[1]) ? 10'b1001000010 : 10'b1001101010;
				assign node166 = (inp[5]) ? node180 : node167;
					assign node167 = (inp[6]) ? node173 : node168;
						assign node168 = (inp[1]) ? 10'b0011100010 : node169;
							assign node169 = (inp[0]) ? 10'b0101001010 : 10'b0001101110;
						assign node173 = (inp[1]) ? node177 : node174;
							assign node174 = (inp[0]) ? 10'b0001101011 : 10'b0111001011;
							assign node177 = (inp[0]) ? 10'b0001000011 : 10'b0101100011;
					assign node180 = (inp[6]) ? node186 : node181;
						assign node181 = (inp[0]) ? node183 : 10'b0000001111;
							assign node183 = (inp[1]) ? 10'b0010000011 : 10'b0010101011;
						assign node186 = (inp[1]) ? node188 : 10'b0110001010;
							assign node188 = (inp[0]) ? 10'b0000000010 : 10'b0100100010;

endmodule