module dtc_split33_bm28 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node9;
	wire [10-1:0] node10;
	wire [10-1:0] node14;
	wire [10-1:0] node15;
	wire [10-1:0] node16;
	wire [10-1:0] node17;
	wire [10-1:0] node22;
	wire [10-1:0] node23;
	wire [10-1:0] node27;
	wire [10-1:0] node28;
	wire [10-1:0] node29;
	wire [10-1:0] node31;
	wire [10-1:0] node34;
	wire [10-1:0] node37;
	wire [10-1:0] node38;
	wire [10-1:0] node41;
	wire [10-1:0] node44;
	wire [10-1:0] node45;
	wire [10-1:0] node46;
	wire [10-1:0] node48;
	wire [10-1:0] node49;
	wire [10-1:0] node52;
	wire [10-1:0] node54;
	wire [10-1:0] node57;
	wire [10-1:0] node58;
	wire [10-1:0] node59;
	wire [10-1:0] node63;
	wire [10-1:0] node65;
	wire [10-1:0] node68;
	wire [10-1:0] node69;
	wire [10-1:0] node71;
	wire [10-1:0] node73;
	wire [10-1:0] node76;
	wire [10-1:0] node77;
	wire [10-1:0] node80;
	wire [10-1:0] node82;

	assign outp = (inp[4]) ? node44 : node1;
		assign node1 = (inp[2]) ? node27 : node2;
			assign node2 = (inp[5]) ? node14 : node3;
				assign node3 = (inp[3]) ? node9 : node4;
					assign node4 = (inp[6]) ? 10'b0111010000 : node5;
						assign node5 = (inp[0]) ? 10'b0101011001 : 10'b0001111101;
					assign node9 = (inp[6]) ? 10'b0101101001 : node10;
						assign node10 = (inp[1]) ? 10'b0001001100 : 10'b0001100101;
				assign node14 = (inp[3]) ? node22 : node15;
					assign node15 = (inp[6]) ? 10'b0110011001 : node16;
						assign node16 = (inp[0]) ? 10'b0010110000 : node17;
							assign node17 = (inp[1]) ? 10'b0000010100 : 10'b0000111100;
					assign node22 = (inp[0]) ? 10'b0000100001 : node23;
						assign node23 = (inp[6]) ? 10'b0110000001 : 10'b0110101001;
			assign node27 = (inp[3]) ? node37 : node28;
				assign node28 = (inp[5]) ? node34 : node29;
					assign node29 = (inp[1]) ? node31 : 10'b1010001000;
						assign node31 = (inp[0]) ? 10'b1000100000 : 10'b1110000000;
					assign node34 = (inp[6]) ? 10'b1001100001 : 10'b1001100100;
				assign node37 = (inp[0]) ? node41 : node38;
					assign node38 = (inp[1]) ? 10'b1101110001 : 10'b1111011001;
					assign node41 = (inp[6]) ? 10'b1000010000 : 10'b1010010001;
		assign node44 = (inp[3]) ? node68 : node45;
			assign node45 = (inp[2]) ? node57 : node46;
				assign node46 = (inp[5]) ? node48 : 10'b1010110011;
					assign node48 = (inp[0]) ? node52 : node49;
						assign node49 = (inp[6]) ? 10'b1101111010 : 10'b1111111011;
						assign node52 = (inp[6]) ? node54 : 10'b1101010010;
							assign node54 = (inp[1]) ? 10'b1001011010 : 10'b1001110011;
				assign node57 = (inp[1]) ? node63 : node58;
					assign node58 = (inp[5]) ? 10'b0110010011 : node59;
						assign node59 = (inp[6]) ? 10'b0011010010 : 10'b0101010011;
					assign node63 = (inp[5]) ? node65 : 10'b0101111011;
						assign node65 = (inp[0]) ? 10'b0010011011 : 10'b0110111011;
			assign node68 = (inp[2]) ? node76 : node69;
				assign node69 = (inp[0]) ? node71 : 10'b1000001110;
					assign node71 = (inp[1]) ? node73 : 10'b1010000010;
						assign node73 = (inp[6]) ? 10'b1001000010 : 10'b1011000011;
				assign node76 = (inp[5]) ? node80 : node77;
					assign node77 = (inp[6]) ? 10'b0101100011 : 10'b0001000110;
					assign node80 = (inp[6]) ? node82 : 10'b0110100011;
						assign node82 = (inp[0]) ? 10'b0000101010 : 10'b0110001010;

endmodule