module dtc_split875_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node6;
	wire [2-1:0] node9;
	wire [2-1:0] node11;
	wire [2-1:0] node14;
	wire [2-1:0] node15;
	wire [2-1:0] node16;
	wire [2-1:0] node19;
	wire [2-1:0] node22;
	wire [2-1:0] node24;
	wire [2-1:0] node27;
	wire [2-1:0] node28;
	wire [2-1:0] node29;
	wire [2-1:0] node32;
	wire [2-1:0] node35;
	wire [2-1:0] node36;
	wire [2-1:0] node37;
	wire [2-1:0] node40;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node47;
	wire [2-1:0] node50;
	wire [2-1:0] node51;
	wire [2-1:0] node52;
	wire [2-1:0] node55;
	wire [2-1:0] node58;
	wire [2-1:0] node59;
	wire [2-1:0] node60;
	wire [2-1:0] node61;
	wire [2-1:0] node64;
	wire [2-1:0] node67;
	wire [2-1:0] node68;
	wire [2-1:0] node72;
	wire [2-1:0] node73;
	wire [2-1:0] node74;
	wire [2-1:0] node77;
	wire [2-1:0] node80;
	wire [2-1:0] node81;
	wire [2-1:0] node84;
	wire [2-1:0] node87;
	wire [2-1:0] node88;
	wire [2-1:0] node89;
	wire [2-1:0] node90;
	wire [2-1:0] node91;
	wire [2-1:0] node94;
	wire [2-1:0] node97;
	wire [2-1:0] node98;
	wire [2-1:0] node99;
	wire [2-1:0] node102;
	wire [2-1:0] node105;
	wire [2-1:0] node106;
	wire [2-1:0] node109;
	wire [2-1:0] node112;
	wire [2-1:0] node113;
	wire [2-1:0] node115;
	wire [2-1:0] node118;
	wire [2-1:0] node119;
	wire [2-1:0] node120;
	wire [2-1:0] node124;
	wire [2-1:0] node125;
	wire [2-1:0] node129;
	wire [2-1:0] node130;
	wire [2-1:0] node131;
	wire [2-1:0] node132;
	wire [2-1:0] node133;
	wire [2-1:0] node137;
	wire [2-1:0] node138;
	wire [2-1:0] node142;
	wire [2-1:0] node143;
	wire [2-1:0] node144;
	wire [2-1:0] node148;
	wire [2-1:0] node151;
	wire [2-1:0] node152;
	wire [2-1:0] node153;
	wire [2-1:0] node154;
	wire [2-1:0] node158;
	wire [2-1:0] node161;
	wire [2-1:0] node162;
	wire [2-1:0] node163;
	wire [2-1:0] node167;
	wire [2-1:0] node168;
	wire [2-1:0] node172;
	wire [2-1:0] node173;
	wire [2-1:0] node174;
	wire [2-1:0] node175;
	wire [2-1:0] node176;
	wire [2-1:0] node177;
	wire [2-1:0] node178;
	wire [2-1:0] node182;
	wire [2-1:0] node183;
	wire [2-1:0] node186;
	wire [2-1:0] node189;
	wire [2-1:0] node190;
	wire [2-1:0] node191;
	wire [2-1:0] node194;
	wire [2-1:0] node197;
	wire [2-1:0] node198;
	wire [2-1:0] node201;
	wire [2-1:0] node204;
	wire [2-1:0] node205;
	wire [2-1:0] node206;
	wire [2-1:0] node207;
	wire [2-1:0] node211;
	wire [2-1:0] node212;
	wire [2-1:0] node215;
	wire [2-1:0] node218;
	wire [2-1:0] node219;
	wire [2-1:0] node222;
	wire [2-1:0] node225;
	wire [2-1:0] node226;
	wire [2-1:0] node227;
	wire [2-1:0] node228;
	wire [2-1:0] node232;
	wire [2-1:0] node233;
	wire [2-1:0] node237;
	wire [2-1:0] node239;
	wire [2-1:0] node240;
	wire [2-1:0] node244;
	wire [2-1:0] node245;
	wire [2-1:0] node246;
	wire [2-1:0] node247;
	wire [2-1:0] node248;
	wire [2-1:0] node249;
	wire [2-1:0] node252;
	wire [2-1:0] node256;
	wire [2-1:0] node257;
	wire [2-1:0] node260;
	wire [2-1:0] node263;
	wire [2-1:0] node264;
	wire [2-1:0] node266;
	wire [2-1:0] node267;
	wire [2-1:0] node270;
	wire [2-1:0] node273;
	wire [2-1:0] node274;
	wire [2-1:0] node276;
	wire [2-1:0] node279;
	wire [2-1:0] node281;
	wire [2-1:0] node284;
	wire [2-1:0] node285;
	wire [2-1:0] node286;
	wire [2-1:0] node287;
	wire [2-1:0] node288;
	wire [2-1:0] node291;
	wire [2-1:0] node294;
	wire [2-1:0] node295;
	wire [2-1:0] node298;
	wire [2-1:0] node301;
	wire [2-1:0] node302;
	wire [2-1:0] node303;
	wire [2-1:0] node306;
	wire [2-1:0] node309;
	wire [2-1:0] node310;
	wire [2-1:0] node313;
	wire [2-1:0] node316;
	wire [2-1:0] node317;
	wire [2-1:0] node319;
	wire [2-1:0] node322;
	wire [2-1:0] node323;
	wire [2-1:0] node326;

	assign outp = (inp[7]) ? node172 : node1;
		assign node1 = (inp[0]) ? node87 : node2;
			assign node2 = (inp[6]) ? node50 : node3;
				assign node3 = (inp[2]) ? node27 : node4;
					assign node4 = (inp[4]) ? node14 : node5;
						assign node5 = (inp[3]) ? node9 : node6;
							assign node6 = (inp[5]) ? 2'b01 : 2'b11;
							assign node9 = (inp[1]) ? node11 : 2'b01;
								assign node11 = (inp[5]) ? 2'b11 : 2'b01;
						assign node14 = (inp[5]) ? node22 : node15;
							assign node15 = (inp[1]) ? node19 : node16;
								assign node16 = (inp[3]) ? 2'b01 : 2'b11;
								assign node19 = (inp[3]) ? 2'b11 : 2'b01;
							assign node22 = (inp[3]) ? node24 : 2'b11;
								assign node24 = (inp[1]) ? 2'b01 : 2'b11;
					assign node27 = (inp[3]) ? node35 : node28;
						assign node28 = (inp[5]) ? node32 : node29;
							assign node29 = (inp[1]) ? 2'b00 : 2'b10;
							assign node32 = (inp[1]) ? 2'b10 : 2'b00;
						assign node35 = (inp[4]) ? node43 : node36;
							assign node36 = (inp[5]) ? node40 : node37;
								assign node37 = (inp[1]) ? 2'b00 : 2'b10;
								assign node40 = (inp[1]) ? 2'b10 : 2'b00;
							assign node43 = (inp[1]) ? node47 : node44;
								assign node44 = (inp[5]) ? 2'b10 : 2'b00;
								assign node47 = (inp[5]) ? 2'b00 : 2'b10;
				assign node50 = (inp[4]) ? node58 : node51;
					assign node51 = (inp[5]) ? node55 : node52;
						assign node52 = (inp[1]) ? 2'b00 : 2'b10;
						assign node55 = (inp[1]) ? 2'b10 : 2'b00;
					assign node58 = (inp[1]) ? node72 : node59;
						assign node59 = (inp[2]) ? node67 : node60;
							assign node60 = (inp[5]) ? node64 : node61;
								assign node61 = (inp[3]) ? 2'b00 : 2'b10;
								assign node64 = (inp[3]) ? 2'b10 : 2'b00;
							assign node67 = (inp[5]) ? 2'b10 : node68;
								assign node68 = (inp[3]) ? 2'b00 : 2'b10;
						assign node72 = (inp[2]) ? node80 : node73;
							assign node73 = (inp[3]) ? node77 : node74;
								assign node74 = (inp[5]) ? 2'b10 : 2'b00;
								assign node77 = (inp[5]) ? 2'b00 : 2'b10;
							assign node80 = (inp[3]) ? node84 : node81;
								assign node81 = (inp[5]) ? 2'b10 : 2'b00;
								assign node84 = (inp[5]) ? 2'b00 : 2'b10;
			assign node87 = (inp[6]) ? node129 : node88;
				assign node88 = (inp[2]) ? node112 : node89;
					assign node89 = (inp[4]) ? node97 : node90;
						assign node90 = (inp[1]) ? node94 : node91;
							assign node91 = (inp[5]) ? 2'b00 : 2'b10;
							assign node94 = (inp[5]) ? 2'b10 : 2'b00;
						assign node97 = (inp[1]) ? node105 : node98;
							assign node98 = (inp[5]) ? node102 : node99;
								assign node99 = (inp[3]) ? 2'b00 : 2'b10;
								assign node102 = (inp[3]) ? 2'b10 : 2'b00;
							assign node105 = (inp[3]) ? node109 : node106;
								assign node106 = (inp[5]) ? 2'b10 : 2'b00;
								assign node109 = (inp[5]) ? 2'b00 : 2'b10;
					assign node112 = (inp[1]) ? node118 : node113;
						assign node113 = (inp[5]) ? node115 : 2'b01;
							assign node115 = (inp[3]) ? 2'b11 : 2'b01;
						assign node118 = (inp[5]) ? node124 : node119;
							assign node119 = (inp[3]) ? 2'b11 : node120;
								assign node120 = (inp[4]) ? 2'b11 : 2'b01;
							assign node124 = (inp[4]) ? 2'b01 : node125;
								assign node125 = (inp[3]) ? 2'b01 : 2'b11;
				assign node129 = (inp[2]) ? node151 : node130;
					assign node130 = (inp[5]) ? node142 : node131;
						assign node131 = (inp[1]) ? node137 : node132;
							assign node132 = (inp[4]) ? 2'b01 : node133;
								assign node133 = (inp[3]) ? 2'b01 : 2'b11;
							assign node137 = (inp[3]) ? 2'b11 : node138;
								assign node138 = (inp[4]) ? 2'b11 : 2'b01;
						assign node142 = (inp[1]) ? node148 : node143;
							assign node143 = (inp[4]) ? 2'b11 : node144;
								assign node144 = (inp[3]) ? 2'b11 : 2'b01;
							assign node148 = (inp[3]) ? 2'b01 : 2'b11;
					assign node151 = (inp[5]) ? node161 : node152;
						assign node152 = (inp[1]) ? node158 : node153;
							assign node153 = (inp[3]) ? 2'b01 : node154;
								assign node154 = (inp[4]) ? 2'b01 : 2'b11;
							assign node158 = (inp[3]) ? 2'b11 : 2'b01;
						assign node161 = (inp[1]) ? node167 : node162;
							assign node162 = (inp[3]) ? 2'b11 : node163;
								assign node163 = (inp[4]) ? 2'b11 : 2'b01;
							assign node167 = (inp[4]) ? 2'b01 : node168;
								assign node168 = (inp[3]) ? 2'b01 : 2'b11;
		assign node172 = (inp[0]) ? node244 : node173;
			assign node173 = (inp[6]) ? node225 : node174;
				assign node174 = (inp[2]) ? node204 : node175;
					assign node175 = (inp[4]) ? node189 : node176;
						assign node176 = (inp[3]) ? node182 : node177;
							assign node177 = (inp[5]) ? 2'b00 : node178;
								assign node178 = (inp[1]) ? 2'b00 : 2'b10;
							assign node182 = (inp[1]) ? node186 : node183;
								assign node183 = (inp[5]) ? 2'b00 : 2'b10;
								assign node186 = (inp[5]) ? 2'b10 : 2'b00;
						assign node189 = (inp[5]) ? node197 : node190;
							assign node190 = (inp[1]) ? node194 : node191;
								assign node191 = (inp[3]) ? 2'b00 : 2'b10;
								assign node194 = (inp[3]) ? 2'b10 : 2'b00;
							assign node197 = (inp[3]) ? node201 : node198;
								assign node198 = (inp[1]) ? 2'b10 : 2'b00;
								assign node201 = (inp[1]) ? 2'b00 : 2'b10;
					assign node204 = (inp[3]) ? node218 : node205;
						assign node205 = (inp[4]) ? node211 : node206;
							assign node206 = (inp[1]) ? 2'b01 : node207;
								assign node207 = (inp[5]) ? 2'b01 : 2'b11;
							assign node211 = (inp[5]) ? node215 : node212;
								assign node212 = (inp[1]) ? 2'b11 : 2'b01;
								assign node215 = (inp[1]) ? 2'b01 : 2'b11;
						assign node218 = (inp[1]) ? node222 : node219;
							assign node219 = (inp[5]) ? 2'b11 : 2'b01;
							assign node222 = (inp[5]) ? 2'b01 : 2'b11;
				assign node225 = (inp[1]) ? node237 : node226;
					assign node226 = (inp[5]) ? node232 : node227;
						assign node227 = (inp[3]) ? 2'b01 : node228;
							assign node228 = (inp[4]) ? 2'b01 : 2'b11;
						assign node232 = (inp[3]) ? 2'b11 : node233;
							assign node233 = (inp[4]) ? 2'b11 : 2'b01;
					assign node237 = (inp[5]) ? node239 : 2'b11;
						assign node239 = (inp[4]) ? 2'b01 : node240;
							assign node240 = (inp[3]) ? 2'b01 : 2'b11;
			assign node244 = (inp[6]) ? node284 : node245;
				assign node245 = (inp[2]) ? node263 : node246;
					assign node246 = (inp[3]) ? node256 : node247;
						assign node247 = (inp[1]) ? 2'b11 : node248;
							assign node248 = (inp[4]) ? node252 : node249;
								assign node249 = (inp[5]) ? 2'b01 : 2'b11;
								assign node252 = (inp[5]) ? 2'b11 : 2'b01;
						assign node256 = (inp[1]) ? node260 : node257;
							assign node257 = (inp[5]) ? 2'b11 : 2'b01;
							assign node260 = (inp[5]) ? 2'b01 : 2'b11;
					assign node263 = (inp[3]) ? node273 : node264;
						assign node264 = (inp[4]) ? node266 : 2'b10;
							assign node266 = (inp[5]) ? node270 : node267;
								assign node267 = (inp[1]) ? 2'b10 : 2'b00;
								assign node270 = (inp[1]) ? 2'b00 : 2'b10;
						assign node273 = (inp[4]) ? node279 : node274;
							assign node274 = (inp[5]) ? node276 : 2'b00;
								assign node276 = (inp[1]) ? 2'b00 : 2'b10;
							assign node279 = (inp[1]) ? node281 : 2'b10;
								assign node281 = (inp[5]) ? 2'b00 : 2'b10;
				assign node284 = (inp[3]) ? node316 : node285;
					assign node285 = (inp[2]) ? node301 : node286;
						assign node286 = (inp[1]) ? node294 : node287;
							assign node287 = (inp[5]) ? node291 : node288;
								assign node288 = (inp[4]) ? 2'b00 : 2'b10;
								assign node291 = (inp[4]) ? 2'b10 : 2'b00;
							assign node294 = (inp[5]) ? node298 : node295;
								assign node295 = (inp[4]) ? 2'b10 : 2'b00;
								assign node298 = (inp[4]) ? 2'b00 : 2'b10;
						assign node301 = (inp[5]) ? node309 : node302;
							assign node302 = (inp[4]) ? node306 : node303;
								assign node303 = (inp[1]) ? 2'b00 : 2'b10;
								assign node306 = (inp[1]) ? 2'b10 : 2'b00;
							assign node309 = (inp[1]) ? node313 : node310;
								assign node310 = (inp[4]) ? 2'b10 : 2'b00;
								assign node313 = (inp[4]) ? 2'b00 : 2'b10;
					assign node316 = (inp[2]) ? node322 : node317;
						assign node317 = (inp[5]) ? node319 : 2'b10;
							assign node319 = (inp[1]) ? 2'b00 : 2'b10;
						assign node322 = (inp[1]) ? node326 : node323;
							assign node323 = (inp[5]) ? 2'b10 : 2'b00;
							assign node326 = (inp[5]) ? 2'b00 : 2'b10;

endmodule