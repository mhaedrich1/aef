module dtc_split33_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;

	assign outp = (inp[9]) ? node326 : node1;
		assign node1 = (inp[6]) ? node145 : node2;
			assign node2 = (inp[10]) ? node60 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? node13 : 3'b111;
										assign node13 = (inp[5]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node37 : node18;
						assign node18 = (inp[8]) ? node28 : node19;
							assign node19 = (inp[4]) ? node21 : 3'b111;
								assign node21 = (inp[0]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? node25 : 3'b111;
										assign node25 = (inp[3]) ? 3'b011 : 3'b111;
							assign node28 = (inp[3]) ? 3'b011 : node29;
								assign node29 = (inp[4]) ? node31 : 3'b111;
									assign node31 = (inp[2]) ? 3'b011 : node32;
										assign node32 = (inp[0]) ? 3'b011 : 3'b111;
						assign node37 = (inp[8]) ? node45 : node38;
							assign node38 = (inp[1]) ? node40 : 3'b011;
								assign node40 = (inp[4]) ? 3'b101 : node41;
									assign node41 = (inp[3]) ? 3'b011 : 3'b111;
							assign node45 = (inp[3]) ? node51 : node46;
								assign node46 = (inp[4]) ? node48 : 3'b011;
									assign node48 = (inp[0]) ? 3'b101 : 3'b011;
								assign node51 = (inp[1]) ? node53 : 3'b101;
									assign node53 = (inp[0]) ? node55 : 3'b101;
										assign node55 = (inp[5]) ? node57 : 3'b101;
											assign node57 = (inp[4]) ? 3'b001 : 3'b101;
				assign node60 = (inp[7]) ? node88 : node61;
					assign node61 = (inp[11]) ? node73 : node62;
						assign node62 = (inp[3]) ? node66 : node63;
							assign node63 = (inp[8]) ? 3'b011 : 3'b111;
							assign node66 = (inp[8]) ? node68 : 3'b011;
								assign node68 = (inp[4]) ? 3'b101 : node69;
									assign node69 = (inp[0]) ? 3'b101 : 3'b011;
						assign node73 = (inp[3]) ? node77 : node74;
							assign node74 = (inp[8]) ? 3'b101 : 3'b011;
							assign node77 = (inp[8]) ? node79 : 3'b101;
								assign node79 = (inp[4]) ? 3'b001 : node80;
									assign node80 = (inp[1]) ? 3'b001 : node81;
										assign node81 = (inp[5]) ? node83 : 3'b101;
											assign node83 = (inp[2]) ? 3'b001 : 3'b101;
					assign node88 = (inp[11]) ? node116 : node89;
						assign node89 = (inp[8]) ? node101 : node90;
							assign node90 = (inp[1]) ? 3'b101 : node91;
								assign node91 = (inp[4]) ? node95 : node92;
									assign node92 = (inp[3]) ? 3'b101 : 3'b011;
									assign node95 = (inp[3]) ? node97 : 3'b101;
										assign node97 = (inp[5]) ? 3'b001 : 3'b101;
							assign node101 = (inp[4]) ? node109 : node102;
								assign node102 = (inp[3]) ? 3'b001 : node103;
									assign node103 = (inp[2]) ? node105 : 3'b101;
										assign node105 = (inp[1]) ? 3'b001 : 3'b101;
								assign node109 = (inp[1]) ? node111 : 3'b001;
									assign node111 = (inp[3]) ? node113 : 3'b001;
										assign node113 = (inp[5]) ? 3'b110 : 3'b001;
						assign node116 = (inp[8]) ? node130 : node117;
							assign node117 = (inp[4]) ? node125 : node118;
								assign node118 = (inp[3]) ? 3'b001 : node119;
									assign node119 = (inp[0]) ? 3'b001 : node120;
										assign node120 = (inp[5]) ? 3'b001 : 3'b101;
								assign node125 = (inp[3]) ? node127 : 3'b001;
									assign node127 = (inp[1]) ? 3'b001 : 3'b110;
							assign node130 = (inp[3]) ? node138 : node131;
								assign node131 = (inp[4]) ? 3'b110 : node132;
									assign node132 = (inp[1]) ? node134 : 3'b001;
										assign node134 = (inp[0]) ? 3'b110 : 3'b001;
								assign node138 = (inp[1]) ? node140 : 3'b110;
									assign node140 = (inp[5]) ? node142 : 3'b110;
										assign node142 = (inp[0]) ? 3'b010 : 3'b110;
			assign node145 = (inp[10]) ? node229 : node146;
				assign node146 = (inp[7]) ? node186 : node147;
					assign node147 = (inp[11]) ? node161 : node148;
						assign node148 = (inp[8]) ? node152 : node149;
							assign node149 = (inp[3]) ? 3'b101 : 3'b011;
							assign node152 = (inp[3]) ? node154 : 3'b101;
								assign node154 = (inp[4]) ? 3'b001 : node155;
									assign node155 = (inp[5]) ? node157 : 3'b101;
										assign node157 = (inp[0]) ? 3'b001 : 3'b101;
						assign node161 = (inp[5]) ? node171 : node162;
							assign node162 = (inp[8]) ? node166 : node163;
								assign node163 = (inp[3]) ? 3'b001 : 3'b101;
								assign node166 = (inp[4]) ? node168 : 3'b001;
									assign node168 = (inp[3]) ? 3'b110 : 3'b001;
							assign node171 = (inp[8]) ? node179 : node172;
								assign node172 = (inp[3]) ? 3'b001 : node173;
									assign node173 = (inp[2]) ? node175 : 3'b101;
										assign node175 = (inp[4]) ? 3'b001 : 3'b101;
								assign node179 = (inp[3]) ? node181 : 3'b001;
									assign node181 = (inp[0]) ? 3'b110 : node182;
										assign node182 = (inp[1]) ? 3'b110 : 3'b001;
					assign node186 = (inp[11]) ? node206 : node187;
						assign node187 = (inp[8]) ? node195 : node188;
							assign node188 = (inp[3]) ? node192 : node189;
								assign node189 = (inp[4]) ? 3'b001 : 3'b101;
								assign node192 = (inp[4]) ? 3'b110 : 3'b001;
							assign node195 = (inp[3]) ? node201 : node196;
								assign node196 = (inp[4]) ? node198 : 3'b001;
									assign node198 = (inp[0]) ? 3'b110 : 3'b001;
								assign node201 = (inp[1]) ? node203 : 3'b110;
									assign node203 = (inp[4]) ? 3'b010 : 3'b110;
						assign node206 = (inp[8]) ? node222 : node207;
							assign node207 = (inp[3]) ? node215 : node208;
								assign node208 = (inp[0]) ? 3'b110 : node209;
									assign node209 = (inp[4]) ? 3'b110 : node210;
										assign node210 = (inp[5]) ? 3'b110 : 3'b001;
								assign node215 = (inp[4]) ? node217 : 3'b110;
									assign node217 = (inp[5]) ? 3'b010 : node218;
										assign node218 = (inp[0]) ? 3'b010 : 3'b110;
							assign node222 = (inp[3]) ? 3'b010 : node223;
								assign node223 = (inp[4]) ? 3'b010 : node224;
									assign node224 = (inp[1]) ? 3'b010 : 3'b110;
				assign node229 = (inp[7]) ? node265 : node230;
					assign node230 = (inp[3]) ? node252 : node231;
						assign node231 = (inp[8]) ? node249 : node232;
							assign node232 = (inp[11]) ? node240 : node233;
								assign node233 = (inp[5]) ? node235 : 3'b001;
									assign node235 = (inp[4]) ? node237 : 3'b001;
										assign node237 = (inp[0]) ? 3'b110 : 3'b001;
								assign node240 = (inp[2]) ? node242 : 3'b110;
									assign node242 = (inp[1]) ? node244 : 3'b110;
										assign node244 = (inp[0]) ? 3'b010 : node245;
											assign node245 = (inp[5]) ? 3'b010 : 3'b110;
							assign node249 = (inp[11]) ? 3'b010 : 3'b110;
						assign node252 = (inp[11]) ? node262 : node253;
							assign node253 = (inp[8]) ? node255 : 3'b110;
								assign node255 = (inp[0]) ? 3'b010 : node256;
									assign node256 = (inp[5]) ? node258 : 3'b010;
										assign node258 = (inp[1]) ? 3'b010 : 3'b110;
							assign node262 = (inp[8]) ? 3'b100 : 3'b010;
					assign node265 = (inp[11]) ? node297 : node266;
						assign node266 = (inp[8]) ? node284 : node267;
							assign node267 = (inp[3]) ? node273 : node268;
								assign node268 = (inp[4]) ? 3'b010 : node269;
									assign node269 = (inp[5]) ? 3'b010 : 3'b110;
								assign node273 = (inp[4]) ? node279 : node274;
									assign node274 = (inp[2]) ? node276 : 3'b010;
										assign node276 = (inp[1]) ? 3'b100 : 3'b010;
									assign node279 = (inp[0]) ? 3'b100 : node280;
										assign node280 = (inp[1]) ? 3'b100 : 3'b010;
							assign node284 = (inp[3]) ? node292 : node285;
								assign node285 = (inp[1]) ? 3'b100 : node286;
									assign node286 = (inp[4]) ? node288 : 3'b010;
										assign node288 = (inp[0]) ? 3'b100 : 3'b010;
								assign node292 = (inp[5]) ? node294 : 3'b100;
									assign node294 = (inp[4]) ? 3'b000 : 3'b100;
						assign node297 = (inp[8]) ? node315 : node298;
							assign node298 = (inp[3]) ? node306 : node299;
								assign node299 = (inp[4]) ? 3'b100 : node300;
									assign node300 = (inp[0]) ? 3'b100 : node301;
										assign node301 = (inp[5]) ? 3'b100 : 3'b010;
								assign node306 = (inp[4]) ? 3'b000 : node307;
									assign node307 = (inp[0]) ? node309 : 3'b100;
										assign node309 = (inp[5]) ? node311 : 3'b100;
											assign node311 = (inp[1]) ? 3'b000 : 3'b100;
							assign node315 = (inp[3]) ? 3'b000 : node316;
								assign node316 = (inp[5]) ? node320 : node317;
									assign node317 = (inp[4]) ? 3'b000 : 3'b100;
									assign node320 = (inp[0]) ? 3'b000 : node321;
										assign node321 = (inp[4]) ? 3'b000 : 3'b100;
		assign node326 = (inp[6]) ? node476 : node327;
			assign node327 = (inp[10]) ? node413 : node328;
				assign node328 = (inp[7]) ? node358 : node329;
					assign node329 = (inp[11]) ? node341 : node330;
						assign node330 = (inp[3]) ? node334 : node331;
							assign node331 = (inp[8]) ? 3'b001 : 3'b101;
							assign node334 = (inp[8]) ? node336 : 3'b001;
								assign node336 = (inp[4]) ? 3'b110 : node337;
									assign node337 = (inp[5]) ? 3'b110 : 3'b001;
						assign node341 = (inp[8]) ? node349 : node342;
							assign node342 = (inp[3]) ? 3'b110 : node343;
								assign node343 = (inp[2]) ? node345 : 3'b001;
									assign node345 = (inp[0]) ? 3'b110 : 3'b001;
							assign node349 = (inp[3]) ? node351 : 3'b110;
								assign node351 = (inp[2]) ? 3'b010 : node352;
									assign node352 = (inp[5]) ? 3'b010 : node353;
										assign node353 = (inp[4]) ? 3'b010 : 3'b110;
					assign node358 = (inp[11]) ? node382 : node359;
						assign node359 = (inp[8]) ? node369 : node360;
							assign node360 = (inp[4]) ? node362 : 3'b110;
								assign node362 = (inp[3]) ? node364 : 3'b110;
									assign node364 = (inp[1]) ? 3'b010 : node365;
										assign node365 = (inp[5]) ? 3'b010 : 3'b110;
							assign node369 = (inp[4]) ? node377 : node370;
								assign node370 = (inp[3]) ? 3'b010 : node371;
									assign node371 = (inp[1]) ? node373 : 3'b110;
										assign node373 = (inp[0]) ? 3'b010 : 3'b110;
								assign node377 = (inp[0]) ? node379 : 3'b010;
									assign node379 = (inp[3]) ? 3'b100 : 3'b010;
						assign node382 = (inp[8]) ? node392 : node383;
							assign node383 = (inp[3]) ? node385 : 3'b010;
								assign node385 = (inp[4]) ? 3'b100 : node386;
									assign node386 = (inp[5]) ? node388 : 3'b010;
										assign node388 = (inp[0]) ? 3'b100 : 3'b010;
							assign node392 = (inp[3]) ? node404 : node393;
								assign node393 = (inp[4]) ? 3'b100 : node394;
									assign node394 = (inp[0]) ? 3'b100 : node395;
										assign node395 = (inp[2]) ? node397 : 3'b010;
											assign node397 = (inp[1]) ? node399 : 3'b010;
												assign node399 = (inp[5]) ? 3'b100 : 3'b010;
								assign node404 = (inp[4]) ? node406 : 3'b100;
									assign node406 = (inp[5]) ? node408 : 3'b100;
										assign node408 = (inp[0]) ? 3'b000 : node409;
											assign node409 = (inp[1]) ? 3'b000 : 3'b100;
				assign node413 = (inp[7]) ? node455 : node414;
					assign node414 = (inp[11]) ? node424 : node415;
						assign node415 = (inp[8]) ? node421 : node416;
							assign node416 = (inp[3]) ? 3'b010 : node417;
								assign node417 = (inp[4]) ? 3'b010 : 3'b110;
							assign node421 = (inp[3]) ? 3'b100 : 3'b010;
						assign node424 = (inp[1]) ? node438 : node425;
							assign node425 = (inp[4]) ? 3'b100 : node426;
								assign node426 = (inp[5]) ? 3'b010 : node427;
									assign node427 = (inp[0]) ? node429 : 3'b100;
										assign node429 = (inp[3]) ? node433 : node430;
											assign node430 = (inp[8]) ? 3'b100 : 3'b010;
											assign node433 = (inp[8]) ? 3'b000 : 3'b100;
							assign node438 = (inp[8]) ? node450 : node439;
								assign node439 = (inp[3]) ? node443 : node440;
									assign node440 = (inp[4]) ? 3'b100 : 3'b010;
									assign node443 = (inp[2]) ? node445 : 3'b100;
										assign node445 = (inp[4]) ? node447 : 3'b100;
											assign node447 = (inp[0]) ? 3'b000 : 3'b100;
								assign node450 = (inp[3]) ? 3'b000 : node451;
									assign node451 = (inp[4]) ? 3'b000 : 3'b100;
					assign node455 = (inp[11]) ? 3'b000 : node456;
						assign node456 = (inp[8]) ? node468 : node457;
							assign node457 = (inp[3]) ? node459 : 3'b100;
								assign node459 = (inp[4]) ? 3'b000 : node460;
									assign node460 = (inp[5]) ? node462 : 3'b100;
										assign node462 = (inp[2]) ? 3'b000 : node463;
											assign node463 = (inp[0]) ? 3'b000 : 3'b100;
							assign node468 = (inp[3]) ? 3'b000 : node469;
								assign node469 = (inp[0]) ? 3'b000 : node470;
									assign node470 = (inp[4]) ? 3'b000 : 3'b100;
			assign node476 = (inp[10]) ? 3'b000 : node477;
				assign node477 = (inp[7]) ? node505 : node478;
					assign node478 = (inp[11]) ? node496 : node479;
						assign node479 = (inp[8]) ? node487 : node480;
							assign node480 = (inp[3]) ? 3'b100 : node481;
								assign node481 = (inp[4]) ? node483 : 3'b010;
									assign node483 = (inp[1]) ? 3'b100 : 3'b010;
							assign node487 = (inp[3]) ? node489 : 3'b100;
								assign node489 = (inp[0]) ? 3'b000 : node490;
									assign node490 = (inp[5]) ? 3'b000 : node491;
										assign node491 = (inp[2]) ? 3'b000 : 3'b100;
						assign node496 = (inp[3]) ? 3'b000 : node497;
							assign node497 = (inp[8]) ? 3'b000 : node498;
								assign node498 = (inp[4]) ? node500 : 3'b100;
									assign node500 = (inp[0]) ? 3'b000 : 3'b100;
					assign node505 = (inp[5]) ? 3'b000 : node506;
						assign node506 = (inp[4]) ? 3'b000 : node507;
							assign node507 = (inp[1]) ? 3'b000 : node508;
								assign node508 = (inp[8]) ? 3'b000 : 3'b100;

endmodule