module dtc_split05_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node20;
	wire [4-1:0] node22;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node28;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node60;
	wire [4-1:0] node61;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node72;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node77;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node96;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node106;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node114;
	wire [4-1:0] node116;
	wire [4-1:0] node118;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node129;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node136;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node145;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node151;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node165;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node188;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node195;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node213;
	wire [4-1:0] node216;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node233;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node240;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node277;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node287;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node342;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node349;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node365;
	wire [4-1:0] node367;
	wire [4-1:0] node371;
	wire [4-1:0] node373;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node401;
	wire [4-1:0] node404;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node430;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node461;
	wire [4-1:0] node466;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node479;
	wire [4-1:0] node481;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node499;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node508;
	wire [4-1:0] node511;
	wire [4-1:0] node512;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node530;
	wire [4-1:0] node532;
	wire [4-1:0] node534;
	wire [4-1:0] node535;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node332 : node3;
			assign node3 = (inp[3]) ? node121 : node4;
				assign node4 = (inp[0]) ? node38 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node20 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[5]) ? node14 : node9;
									assign node9 = (inp[1]) ? 4'b0010 : node10;
										assign node10 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node14 = (inp[13]) ? node16 : 4'b0000;
										assign node16 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node20 = (inp[7]) ? node22 : 4'b0000;
								assign node22 = (inp[5]) ? node28 : node23;
									assign node23 = (inp[9]) ? 4'b0010 : node24;
										assign node24 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node28 = (inp[9]) ? node30 : 4'b0000;
										assign node30 = (inp[13]) ? 4'b0010 : node31;
											assign node31 = (inp[2]) ? 4'b0000 : node32;
												assign node32 = (inp[15]) ? 4'b0000 : 4'b0010;
					assign node38 = (inp[4]) ? node96 : node39;
						assign node39 = (inp[10]) ? node65 : node40;
							assign node40 = (inp[11]) ? node52 : node41;
								assign node41 = (inp[7]) ? node47 : node42;
									assign node42 = (inp[9]) ? 4'b0000 : node43;
										assign node43 = (inp[8]) ? 4'b0010 : 4'b0000;
									assign node47 = (inp[9]) ? 4'b0010 : node48;
										assign node48 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node52 = (inp[7]) ? node60 : node53;
									assign node53 = (inp[2]) ? 4'b0010 : node54;
										assign node54 = (inp[9]) ? node56 : 4'b0010;
											assign node56 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node60 = (inp[2]) ? 4'b0000 : node61;
										assign node61 = (inp[9]) ? 4'b0010 : 4'b0000;
							assign node65 = (inp[7]) ? node81 : node66;
								assign node66 = (inp[11]) ? node72 : node67;
									assign node67 = (inp[9]) ? 4'b0000 : node68;
										assign node68 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node72 = (inp[2]) ? node74 : 4'b0010;
										assign node74 = (inp[8]) ? 4'b0000 : node75;
											assign node75 = (inp[9]) ? node77 : 4'b0010;
												assign node77 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node81 = (inp[9]) ? node83 : 4'b0000;
									assign node83 = (inp[5]) ? node89 : node84;
										assign node84 = (inp[8]) ? 4'b0010 : node85;
											assign node85 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node89 = (inp[11]) ? 4'b0000 : node90;
											assign node90 = (inp[6]) ? 4'b0010 : node91;
												assign node91 = (inp[13]) ? 4'b0010 : 4'b0000;
						assign node96 = (inp[7]) ? node98 : 4'b0010;
							assign node98 = (inp[11]) ? node106 : node99;
								assign node99 = (inp[5]) ? node101 : 4'b0000;
									assign node101 = (inp[9]) ? 4'b0000 : node102;
										assign node102 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node106 = (inp[9]) ? node108 : 4'b0010;
									assign node108 = (inp[13]) ? node114 : node109;
										assign node109 = (inp[5]) ? 4'b0010 : node110;
											assign node110 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node114 = (inp[10]) ? node116 : 4'b0000;
											assign node116 = (inp[15]) ? node118 : 4'b0000;
												assign node118 = (inp[1]) ? 4'b0000 : 4'b0010;
				assign node121 = (inp[0]) ? node155 : node122;
					assign node122 = (inp[4]) ? node124 : 4'b0010;
						assign node124 = (inp[7]) ? node140 : node125;
							assign node125 = (inp[11]) ? 4'b0000 : node126;
								assign node126 = (inp[9]) ? node132 : node127;
									assign node127 = (inp[13]) ? node129 : 4'b0000;
										assign node129 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node132 = (inp[5]) ? node134 : 4'b0010;
										assign node134 = (inp[13]) ? node136 : 4'b0000;
											assign node136 = (inp[1]) ? 4'b0010 : 4'b0000;
							assign node140 = (inp[11]) ? node142 : 4'b0010;
								assign node142 = (inp[9]) ? node148 : node143;
									assign node143 = (inp[13]) ? node145 : 4'b0000;
										assign node145 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node148 = (inp[1]) ? 4'b0010 : node149;
										assign node149 = (inp[6]) ? node151 : 4'b0010;
											assign node151 = (inp[10]) ? 4'b0010 : 4'b0000;
					assign node155 = (inp[9]) ? node223 : node156;
						assign node156 = (inp[7]) ? node178 : node157;
							assign node157 = (inp[4]) ? node165 : node158;
								assign node158 = (inp[11]) ? 4'b0010 : node159;
									assign node159 = (inp[2]) ? 4'b1000 : node160;
										assign node160 = (inp[10]) ? 4'b1000 : 4'b0010;
								assign node165 = (inp[11]) ? 4'b0000 : node166;
									assign node166 = (inp[13]) ? 4'b0010 : node167;
										assign node167 = (inp[1]) ? node173 : node168;
											assign node168 = (inp[8]) ? node170 : 4'b0000;
												assign node170 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node173 = (inp[2]) ? 4'b0010 : 4'b0000;
							assign node178 = (inp[4]) ? node206 : node179;
								assign node179 = (inp[1]) ? node191 : node180;
									assign node180 = (inp[6]) ? node182 : 4'b0000;
										assign node182 = (inp[11]) ? node188 : node183;
											assign node183 = (inp[8]) ? 4'b0010 : node184;
												assign node184 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node188 = (inp[13]) ? 4'b0000 : 4'b1010;
									assign node191 = (inp[11]) ? node199 : node192;
										assign node192 = (inp[6]) ? 4'b1000 : node193;
											assign node193 = (inp[10]) ? node195 : 4'b1010;
												assign node195 = (inp[2]) ? 4'b1010 : 4'b1000;
										assign node199 = (inp[6]) ? node201 : 4'b0010;
											assign node201 = (inp[15]) ? 4'b0000 : node202;
												assign node202 = (inp[10]) ? 4'b1010 : 4'b1000;
								assign node206 = (inp[11]) ? node210 : node207;
									assign node207 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node210 = (inp[8]) ? node216 : node211;
										assign node211 = (inp[1]) ? node213 : 4'b1010;
											assign node213 = (inp[13]) ? 4'b0010 : 4'b1010;
										assign node216 = (inp[5]) ? node218 : 4'b1000;
											assign node218 = (inp[13]) ? 4'b1010 : node219;
												assign node219 = (inp[15]) ? 4'b1000 : 4'b1010;
						assign node223 = (inp[7]) ? node273 : node224;
							assign node224 = (inp[4]) ? node252 : node225;
								assign node225 = (inp[8]) ? node237 : node226;
									assign node226 = (inp[13]) ? 4'b1000 : node227;
										assign node227 = (inp[5]) ? node233 : node228;
											assign node228 = (inp[2]) ? 4'b1000 : node229;
												assign node229 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node233 = (inp[11]) ? 4'b1000 : 4'b1010;
									assign node237 = (inp[10]) ? node243 : node238;
										assign node238 = (inp[1]) ? node240 : 4'b1010;
											assign node240 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node243 = (inp[5]) ? node247 : node244;
											assign node244 = (inp[13]) ? 4'b1000 : 4'b1010;
											assign node247 = (inp[13]) ? 4'b1010 : node248;
												assign node248 = (inp[11]) ? 4'b1000 : 4'b1010;
								assign node252 = (inp[6]) ? node262 : node253;
									assign node253 = (inp[15]) ? 4'b0010 : node254;
										assign node254 = (inp[2]) ? node258 : node255;
											assign node255 = (inp[5]) ? 4'b0000 : 4'b1000;
											assign node258 = (inp[8]) ? 4'b0010 : 4'b1010;
									assign node262 = (inp[10]) ? node268 : node263;
										assign node263 = (inp[13]) ? 4'b1000 : node264;
											assign node264 = (inp[1]) ? 4'b1000 : 4'b0010;
										assign node268 = (inp[11]) ? 4'b0010 : node269;
											assign node269 = (inp[8]) ? 4'b1000 : 4'b1010;
							assign node273 = (inp[4]) ? node295 : node274;
								assign node274 = (inp[1]) ? node282 : node275;
									assign node275 = (inp[5]) ? node277 : 4'b0011;
										assign node277 = (inp[13]) ? node279 : 4'b0001;
											assign node279 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node282 = (inp[6]) ? node290 : node283;
										assign node283 = (inp[15]) ? node287 : node284;
											assign node284 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node287 = (inp[11]) ? 4'b0011 : 4'b0111;
										assign node290 = (inp[8]) ? 4'b0000 : node291;
											assign node291 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node295 = (inp[13]) ? node317 : node296;
									assign node296 = (inp[1]) ? node306 : node297;
										assign node297 = (inp[15]) ? node301 : node298;
											assign node298 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node301 = (inp[6]) ? 4'b1000 : node302;
												assign node302 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node306 = (inp[11]) ? node314 : node307;
											assign node307 = (inp[6]) ? node311 : node308;
												assign node308 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node311 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node314 = (inp[6]) ? 4'b0011 : 4'b1010;
									assign node317 = (inp[6]) ? node325 : node318;
										assign node318 = (inp[10]) ? 4'b1011 : node319;
											assign node319 = (inp[5]) ? 4'b1110 : node320;
												assign node320 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node325 = (inp[1]) ? 4'b0000 : node326;
											assign node326 = (inp[5]) ? 4'b0010 : node327;
												assign node327 = (inp[8]) ? 4'b1000 : 4'b1010;
			assign node332 = (inp[0]) ? node334 : 4'b0000;
				assign node334 = (inp[4]) ? node466 : node335;
					assign node335 = (inp[7]) ? node395 : node336;
						assign node336 = (inp[9]) ? node360 : node337;
							assign node337 = (inp[11]) ? node357 : node338;
								assign node338 = (inp[8]) ? node346 : node339;
									assign node339 = (inp[3]) ? 4'b0000 : node340;
										assign node340 = (inp[6]) ? node342 : 4'b0000;
											assign node342 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node346 = (inp[6]) ? node352 : node347;
										assign node347 = (inp[3]) ? node349 : 4'b0000;
											assign node349 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node352 = (inp[10]) ? node354 : 4'b0010;
											assign node354 = (inp[3]) ? 4'b0010 : 4'b0000;
								assign node357 = (inp[3]) ? 4'b0010 : 4'b0000;
							assign node360 = (inp[11]) ? node380 : node361;
								assign node361 = (inp[13]) ? node371 : node362;
									assign node362 = (inp[3]) ? 4'b0000 : node363;
										assign node363 = (inp[5]) ? node365 : 4'b0010;
											assign node365 = (inp[6]) ? node367 : 4'b0000;
												assign node367 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node371 = (inp[5]) ? node373 : 4'b0010;
										assign node373 = (inp[15]) ? node375 : 4'b0010;
											assign node375 = (inp[6]) ? 4'b0000 : node376;
												assign node376 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node380 = (inp[3]) ? node382 : 4'b0000;
									assign node382 = (inp[15]) ? node388 : node383;
										assign node383 = (inp[1]) ? 4'b0000 : node384;
											assign node384 = (inp[13]) ? 4'b0000 : 4'b0010;
										assign node388 = (inp[5]) ? 4'b0010 : node389;
											assign node389 = (inp[13]) ? 4'b0000 : node390;
												assign node390 = (inp[6]) ? 4'b0000 : 4'b0010;
						assign node395 = (inp[3]) ? node411 : node396;
							assign node396 = (inp[11]) ? node398 : 4'b0010;
								assign node398 = (inp[9]) ? node404 : node399;
									assign node399 = (inp[1]) ? node401 : 4'b0000;
										assign node401 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node404 = (inp[6]) ? node406 : 4'b0010;
										assign node406 = (inp[1]) ? 4'b0010 : node407;
											assign node407 = (inp[5]) ? 4'b0000 : 4'b0010;
							assign node411 = (inp[13]) ? node439 : node412;
								assign node412 = (inp[11]) ? node424 : node413;
									assign node413 = (inp[5]) ? node415 : 4'b1000;
										assign node415 = (inp[2]) ? node421 : node416;
											assign node416 = (inp[9]) ? node418 : 4'b0010;
												assign node418 = (inp[6]) ? 4'b0000 : 4'b1010;
											assign node421 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node424 = (inp[8]) ? node434 : node425;
										assign node425 = (inp[1]) ? 4'b0010 : node426;
											assign node426 = (inp[15]) ? node430 : node427;
												assign node427 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node430 = (inp[6]) ? 4'b1010 : 4'b1000;
										assign node434 = (inp[9]) ? 4'b0000 : node435;
											assign node435 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node439 = (inp[9]) ? node453 : node440;
									assign node440 = (inp[8]) ? node448 : node441;
										assign node441 = (inp[1]) ? node445 : node442;
											assign node442 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node445 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node448 = (inp[6]) ? 4'b1000 : node449;
											assign node449 = (inp[11]) ? 4'b1000 : 4'b1010;
									assign node453 = (inp[11]) ? node459 : node454;
										assign node454 = (inp[1]) ? 4'b0000 : node455;
											assign node455 = (inp[6]) ? 4'b1001 : 4'b0001;
										assign node459 = (inp[6]) ? 4'b0001 : node460;
											assign node460 = (inp[15]) ? 4'b0010 : node461;
												assign node461 = (inp[10]) ? 4'b1000 : 4'b1010;
					assign node466 = (inp[3]) ? node468 : 4'b0000;
						assign node468 = (inp[7]) ? node486 : node469;
							assign node469 = (inp[11]) ? 4'b0000 : node470;
								assign node470 = (inp[5]) ? node476 : node471;
									assign node471 = (inp[13]) ? 4'b0010 : node472;
										assign node472 = (inp[9]) ? 4'b0010 : 4'b0000;
									assign node476 = (inp[10]) ? 4'b0000 : node477;
										assign node477 = (inp[15]) ? node479 : 4'b0010;
											assign node479 = (inp[1]) ? node481 : 4'b0000;
												assign node481 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node486 = (inp[2]) ? node516 : node487;
								assign node487 = (inp[9]) ? node503 : node488;
									assign node488 = (inp[15]) ? node498 : node489;
										assign node489 = (inp[8]) ? node491 : 4'b0010;
											assign node491 = (inp[6]) ? node495 : node492;
												assign node492 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node495 = (inp[10]) ? 4'b0010 : 4'b0000;
										assign node498 = (inp[1]) ? 4'b0000 : node499;
											assign node499 = (inp[11]) ? 4'b0000 : 4'b0010;
									assign node503 = (inp[10]) ? node511 : node504;
										assign node504 = (inp[11]) ? node506 : 4'b0011;
											assign node506 = (inp[1]) ? node508 : 4'b0010;
												assign node508 = (inp[15]) ? 4'b0010 : 4'b1010;
										assign node511 = (inp[8]) ? 4'b1000 : node512;
											assign node512 = (inp[6]) ? 4'b1010 : 4'b0010;
								assign node516 = (inp[1]) ? node530 : node517;
									assign node517 = (inp[15]) ? 4'b0000 : node518;
										assign node518 = (inp[6]) ? node526 : node519;
											assign node519 = (inp[13]) ? node523 : node520;
												assign node520 = (inp[11]) ? 4'b0010 : 4'b1000;
												assign node523 = (inp[11]) ? 4'b1000 : 4'b0010;
											assign node526 = (inp[9]) ? 4'b1000 : 4'b0000;
									assign node530 = (inp[10]) ? node532 : 4'b0010;
										assign node532 = (inp[15]) ? node534 : 4'b0010;
											assign node534 = (inp[8]) ? 4'b0000 : node535;
												assign node535 = (inp[9]) ? 4'b1000 : 4'b0000;

endmodule