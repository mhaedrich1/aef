module dtc_split875_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node511;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node813;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node896;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1006;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1038;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1047;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1073;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1083;
	wire [3-1:0] node1086;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1112;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1132;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1143;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1168;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;

	assign outp = (inp[6]) ? node248 : node1;
		assign node1 = (inp[7]) ? node39 : node2;
			assign node2 = (inp[1]) ? 3'b000 : node3;
				assign node3 = (inp[10]) ? 3'b000 : node4;
					assign node4 = (inp[9]) ? 3'b000 : node5;
						assign node5 = (inp[0]) ? node7 : 3'b000;
							assign node7 = (inp[8]) ? node9 : 3'b000;
								assign node9 = (inp[3]) ? node29 : node10;
									assign node10 = (inp[5]) ? node18 : node11;
										assign node11 = (inp[11]) ? node15 : node12;
											assign node12 = (inp[2]) ? 3'b000 : 3'b100;
											assign node15 = (inp[2]) ? 3'b100 : 3'b000;
										assign node18 = (inp[4]) ? node24 : node19;
											assign node19 = (inp[2]) ? 3'b000 : node20;
												assign node20 = (inp[11]) ? 3'b000 : 3'b100;
											assign node24 = (inp[2]) ? node26 : 3'b000;
												assign node26 = (inp[11]) ? 3'b100 : 3'b000;
									assign node29 = (inp[11]) ? node33 : node30;
										assign node30 = (inp[2]) ? 3'b000 : 3'b100;
										assign node33 = (inp[2]) ? 3'b100 : 3'b000;
			assign node39 = (inp[9]) ? node207 : node40;
				assign node40 = (inp[0]) ? node130 : node41;
					assign node41 = (inp[10]) ? node89 : node42;
						assign node42 = (inp[1]) ? node46 : node43;
							assign node43 = (inp[11]) ? 3'b001 : 3'b101;
							assign node46 = (inp[8]) ? node62 : node47;
								assign node47 = (inp[11]) ? node55 : node48;
									assign node48 = (inp[2]) ? node50 : 3'b110;
										assign node50 = (inp[3]) ? 3'b010 : node51;
											assign node51 = (inp[4]) ? 3'b010 : 3'b110;
									assign node55 = (inp[2]) ? node57 : 3'b010;
										assign node57 = (inp[3]) ? 3'b110 : node58;
											assign node58 = (inp[4]) ? 3'b110 : 3'b010;
								assign node62 = (inp[11]) ? node76 : node63;
									assign node63 = (inp[4]) ? 3'b001 : node64;
										assign node64 = (inp[2]) ? node70 : node65;
											assign node65 = (inp[5]) ? 3'b001 : node66;
												assign node66 = (inp[3]) ? 3'b001 : 3'b101;
											assign node70 = (inp[5]) ? 3'b110 : node71;
												assign node71 = (inp[3]) ? 3'b110 : 3'b001;
									assign node76 = (inp[4]) ? 3'b110 : node77;
										assign node77 = (inp[3]) ? node83 : node78;
											assign node78 = (inp[2]) ? node80 : 3'b001;
												assign node80 = (inp[5]) ? 3'b010 : 3'b110;
											assign node83 = (inp[2]) ? node85 : 3'b110;
												assign node85 = (inp[5]) ? 3'b010 : 3'b110;
						assign node89 = (inp[1]) ? node91 : 3'b110;
							assign node91 = (inp[8]) ? node95 : node92;
								assign node92 = (inp[11]) ? 3'b000 : 3'b100;
								assign node95 = (inp[11]) ? node115 : node96;
									assign node96 = (inp[2]) ? node104 : node97;
										assign node97 = (inp[3]) ? 3'b010 : node98;
											assign node98 = (inp[5]) ? 3'b010 : node99;
												assign node99 = (inp[4]) ? 3'b010 : 3'b110;
										assign node104 = (inp[3]) ? node110 : node105;
											assign node105 = (inp[5]) ? node107 : 3'b010;
												assign node107 = (inp[4]) ? 3'b010 : 3'b110;
											assign node110 = (inp[5]) ? 3'b100 : node111;
												assign node111 = (inp[4]) ? 3'b100 : 3'b010;
									assign node115 = (inp[4]) ? 3'b100 : node116;
										assign node116 = (inp[5]) ? node122 : node117;
											assign node117 = (inp[2]) ? 3'b110 : node118;
												assign node118 = (inp[3]) ? 3'b110 : 3'b010;
											assign node122 = (inp[3]) ? node126 : node123;
												assign node123 = (inp[2]) ? 3'b010 : 3'b110;
												assign node126 = (inp[2]) ? 3'b000 : 3'b100;
					assign node130 = (inp[10]) ? node194 : node131;
						assign node131 = (inp[1]) ? node165 : node132;
							assign node132 = (inp[11]) ? node150 : node133;
								assign node133 = (inp[8]) ? node143 : node134;
									assign node134 = (inp[2]) ? node136 : 3'b010;
										assign node136 = (inp[5]) ? node138 : 3'b100;
											assign node138 = (inp[4]) ? 3'b100 : node139;
												assign node139 = (inp[3]) ? 3'b100 : 3'b010;
									assign node143 = (inp[2]) ? node145 : 3'b110;
										assign node145 = (inp[4]) ? 3'b010 : node146;
											assign node146 = (inp[3]) ? 3'b010 : 3'b110;
								assign node150 = (inp[8]) ? node158 : node151;
									assign node151 = (inp[2]) ? node153 : 3'b100;
										assign node153 = (inp[4]) ? 3'b010 : node154;
											assign node154 = (inp[3]) ? 3'b010 : 3'b100;
									assign node158 = (inp[2]) ? node160 : 3'b010;
										assign node160 = (inp[3]) ? 3'b100 : node161;
											assign node161 = (inp[4]) ? 3'b100 : 3'b010;
							assign node165 = (inp[8]) ? node173 : node166;
								assign node166 = (inp[2]) ? 3'b000 : node167;
									assign node167 = (inp[11]) ? 3'b000 : node168;
										assign node168 = (inp[3]) ? 3'b000 : 3'b100;
								assign node173 = (inp[11]) ? node183 : node174;
									assign node174 = (inp[2]) ? 3'b100 : node175;
										assign node175 = (inp[3]) ? 3'b100 : node176;
											assign node176 = (inp[5]) ? node178 : 3'b010;
												assign node178 = (inp[4]) ? 3'b010 : 3'b100;
									assign node183 = (inp[2]) ? node189 : node184;
										assign node184 = (inp[3]) ? node186 : 3'b100;
											assign node186 = (inp[4]) ? 3'b000 : 3'b100;
										assign node189 = (inp[4]) ? 3'b000 : node190;
											assign node190 = (inp[5]) ? 3'b100 : 3'b000;
						assign node194 = (inp[1]) ? 3'b000 : node195;
							assign node195 = (inp[11]) ? 3'b000 : node196;
								assign node196 = (inp[8]) ? node198 : 3'b000;
									assign node198 = (inp[2]) ? node200 : 3'b100;
										assign node200 = (inp[3]) ? 3'b000 : node201;
											assign node201 = (inp[4]) ? 3'b000 : 3'b100;
				assign node207 = (inp[10]) ? 3'b000 : node208;
					assign node208 = (inp[0]) ? 3'b000 : node209;
						assign node209 = (inp[1]) ? node217 : node210;
							assign node210 = (inp[2]) ? node214 : node211;
								assign node211 = (inp[11]) ? 3'b110 : 3'b010;
								assign node214 = (inp[11]) ? 3'b000 : 3'b100;
							assign node217 = (inp[8]) ? node219 : 3'b000;
								assign node219 = (inp[3]) ? node235 : node220;
									assign node220 = (inp[4]) ? 3'b000 : node221;
										assign node221 = (inp[5]) ? node227 : node222;
											assign node222 = (inp[11]) ? node224 : 3'b000;
												assign node224 = (inp[2]) ? 3'b100 : 3'b000;
											assign node227 = (inp[11]) ? node231 : node228;
												assign node228 = (inp[2]) ? 3'b000 : 3'b100;
												assign node231 = (inp[2]) ? 3'b100 : 3'b000;
									assign node235 = (inp[11]) ? node241 : node236;
										assign node236 = (inp[2]) ? node238 : 3'b000;
											assign node238 = (inp[4]) ? 3'b100 : 3'b000;
										assign node241 = (inp[4]) ? node243 : 3'b100;
											assign node243 = (inp[2]) ? 3'b000 : 3'b100;
		assign node248 = (inp[9]) ? node804 : node249;
			assign node249 = (inp[0]) ? node545 : node250;
				assign node250 = (inp[7]) ? node442 : node251;
					assign node251 = (inp[10]) ? node337 : node252;
						assign node252 = (inp[1]) ? node282 : node253;
							assign node253 = (inp[8]) ? node265 : node254;
								assign node254 = (inp[11]) ? node260 : node255;
									assign node255 = (inp[2]) ? 3'b011 : node256;
										assign node256 = (inp[3]) ? 3'b011 : 3'b111;
									assign node260 = (inp[2]) ? 3'b101 : node261;
										assign node261 = (inp[3]) ? 3'b101 : 3'b001;
								assign node265 = (inp[11]) ? node273 : node266;
									assign node266 = (inp[2]) ? 3'b111 : node267;
										assign node267 = (inp[3]) ? node269 : 3'b011;
											assign node269 = (inp[4]) ? 3'b111 : 3'b011;
									assign node273 = (inp[2]) ? 3'b011 : node274;
										assign node274 = (inp[3]) ? node276 : 3'b111;
											assign node276 = (inp[4]) ? 3'b011 : node277;
												assign node277 = (inp[5]) ? 3'b011 : 3'b111;
							assign node282 = (inp[8]) ? node314 : node283;
								assign node283 = (inp[11]) ? node301 : node284;
									assign node284 = (inp[2]) ? node292 : node285;
										assign node285 = (inp[4]) ? 3'b101 : node286;
											assign node286 = (inp[3]) ? 3'b101 : node287;
												assign node287 = (inp[5]) ? 3'b110 : 3'b010;
										assign node292 = (inp[3]) ? node298 : node293;
											assign node293 = (inp[5]) ? node295 : 3'b101;
												assign node295 = (inp[4]) ? 3'b101 : 3'b001;
											assign node298 = (inp[4]) ? 3'b001 : 3'b101;
									assign node301 = (inp[3]) ? node307 : node302;
										assign node302 = (inp[4]) ? 3'b001 : node303;
											assign node303 = (inp[2]) ? 3'b001 : 3'b101;
										assign node307 = (inp[5]) ? node309 : 3'b001;
											assign node309 = (inp[2]) ? node311 : 3'b001;
												assign node311 = (inp[4]) ? 3'b110 : 3'b001;
								assign node314 = (inp[11]) ? node326 : node315;
									assign node315 = (inp[4]) ? node321 : node316;
										assign node316 = (inp[3]) ? 3'b011 : node317;
											assign node317 = (inp[2]) ? 3'b011 : 3'b101;
										assign node321 = (inp[2]) ? node323 : 3'b011;
											assign node323 = (inp[3]) ? 3'b101 : 3'b011;
									assign node326 = (inp[3]) ? node332 : node327;
										assign node327 = (inp[2]) ? 3'b101 : node328;
											assign node328 = (inp[4]) ? 3'b101 : 3'b011;
										assign node332 = (inp[2]) ? node334 : 3'b101;
											assign node334 = (inp[4]) ? 3'b001 : 3'b101;
						assign node337 = (inp[1]) ? node389 : node338;
							assign node338 = (inp[8]) ? node370 : node339;
								assign node339 = (inp[11]) ? node351 : node340;
									assign node340 = (inp[2]) ? 3'b001 : node341;
										assign node341 = (inp[5]) ? node347 : node342;
											assign node342 = (inp[4]) ? node344 : 3'b101;
												assign node344 = (inp[3]) ? 3'b001 : 3'b101;
											assign node347 = (inp[4]) ? 3'b101 : 3'b001;
									assign node351 = (inp[5]) ? node361 : node352;
										assign node352 = (inp[2]) ? node358 : node353;
											assign node353 = (inp[3]) ? node355 : 3'b001;
												assign node355 = (inp[4]) ? 3'b101 : 3'b001;
											assign node358 = (inp[4]) ? 3'b101 : 3'b111;
										assign node361 = (inp[2]) ? node367 : node362;
											assign node362 = (inp[3]) ? node364 : 3'b001;
												assign node364 = (inp[4]) ? 3'b110 : 3'b000;
											assign node367 = (inp[4]) ? 3'b110 : 3'b010;
								assign node370 = (inp[11]) ? node378 : node371;
									assign node371 = (inp[2]) ? 3'b101 : node372;
										assign node372 = (inp[3]) ? node374 : 3'b011;
											assign node374 = (inp[4]) ? 3'b101 : 3'b011;
									assign node378 = (inp[2]) ? node384 : node379;
										assign node379 = (inp[4]) ? node381 : 3'b101;
											assign node381 = (inp[3]) ? 3'b001 : 3'b101;
										assign node384 = (inp[5]) ? 3'b001 : node385;
											assign node385 = (inp[4]) ? 3'b011 : 3'b001;
							assign node389 = (inp[8]) ? node413 : node390;
								assign node390 = (inp[11]) ? node402 : node391;
									assign node391 = (inp[3]) ? node397 : node392;
										assign node392 = (inp[4]) ? 3'b110 : node393;
											assign node393 = (inp[2]) ? 3'b110 : 3'b001;
										assign node397 = (inp[2]) ? node399 : 3'b110;
											assign node399 = (inp[4]) ? 3'b010 : 3'b110;
									assign node402 = (inp[3]) ? node408 : node403;
										assign node403 = (inp[2]) ? 3'b010 : node404;
											assign node404 = (inp[4]) ? 3'b010 : 3'b110;
										assign node408 = (inp[2]) ? node410 : 3'b010;
											assign node410 = (inp[4]) ? 3'b100 : 3'b010;
								assign node413 = (inp[11]) ? node427 : node414;
									assign node414 = (inp[3]) ? node420 : node415;
										assign node415 = (inp[2]) ? 3'b001 : node416;
											assign node416 = (inp[4]) ? 3'b001 : 3'b101;
										assign node420 = (inp[4]) ? node422 : 3'b001;
											assign node422 = (inp[2]) ? node424 : 3'b001;
												assign node424 = (inp[5]) ? 3'b110 : 3'b101;
									assign node427 = (inp[4]) ? node433 : node428;
										assign node428 = (inp[3]) ? 3'b110 : node429;
											assign node429 = (inp[2]) ? 3'b110 : 3'b010;
										assign node433 = (inp[3]) ? node435 : 3'b001;
											assign node435 = (inp[5]) ? node439 : node436;
												assign node436 = (inp[2]) ? 3'b001 : 3'b101;
												assign node439 = (inp[2]) ? 3'b010 : 3'b110;
					assign node442 = (inp[10]) ? node480 : node443;
						assign node443 = (inp[8]) ? 3'b111 : node444;
							assign node444 = (inp[1]) ? node446 : 3'b111;
								assign node446 = (inp[11]) ? node462 : node447;
									assign node447 = (inp[2]) ? node455 : node448;
										assign node448 = (inp[3]) ? 3'b111 : node449;
											assign node449 = (inp[4]) ? node451 : 3'b011;
												assign node451 = (inp[5]) ? 3'b011 : 3'b111;
										assign node455 = (inp[5]) ? node457 : 3'b111;
											assign node457 = (inp[3]) ? node459 : 3'b111;
												assign node459 = (inp[4]) ? 3'b011 : 3'b111;
									assign node462 = (inp[5]) ? node470 : node463;
										assign node463 = (inp[3]) ? 3'b011 : node464;
											assign node464 = (inp[2]) ? 3'b011 : node465;
												assign node465 = (inp[4]) ? 3'b011 : 3'b111;
										assign node470 = (inp[2]) ? node474 : node471;
											assign node471 = (inp[3]) ? 3'b011 : 3'b111;
											assign node474 = (inp[4]) ? node476 : 3'b011;
												assign node476 = (inp[3]) ? 3'b101 : 3'b011;
						assign node480 = (inp[1]) ? node516 : node481;
							assign node481 = (inp[8]) ? node511 : node482;
								assign node482 = (inp[5]) ? node492 : node483;
									assign node483 = (inp[11]) ? node487 : node484;
										assign node484 = (inp[2]) ? 3'b011 : 3'b111;
										assign node487 = (inp[2]) ? node489 : 3'b011;
											assign node489 = (inp[4]) ? 3'b111 : 3'b011;
									assign node492 = (inp[11]) ? node500 : node493;
										assign node493 = (inp[2]) ? 3'b011 : node494;
											assign node494 = (inp[3]) ? node496 : 3'b111;
												assign node496 = (inp[4]) ? 3'b011 : 3'b111;
										assign node500 = (inp[4]) ? node506 : node501;
											assign node501 = (inp[3]) ? 3'b001 : node502;
												assign node502 = (inp[2]) ? 3'b001 : 3'b011;
											assign node506 = (inp[3]) ? 3'b101 : node507;
												assign node507 = (inp[2]) ? 3'b101 : 3'b011;
								assign node511 = (inp[2]) ? node513 : 3'b111;
									assign node513 = (inp[11]) ? 3'b011 : 3'b111;
							assign node516 = (inp[11]) ? node532 : node517;
								assign node517 = (inp[8]) ? node523 : node518;
									assign node518 = (inp[2]) ? 3'b101 : node519;
										assign node519 = (inp[3]) ? 3'b101 : 3'b011;
									assign node523 = (inp[2]) ? 3'b011 : node524;
										assign node524 = (inp[3]) ? node526 : 3'b111;
											assign node526 = (inp[5]) ? 3'b011 : node527;
												assign node527 = (inp[4]) ? 3'b011 : 3'b111;
								assign node532 = (inp[8]) ? node538 : node533;
									assign node533 = (inp[3]) ? 3'b001 : node534;
										assign node534 = (inp[2]) ? 3'b001 : 3'b101;
									assign node538 = (inp[2]) ? 3'b101 : node539;
										assign node539 = (inp[3]) ? node541 : 3'b001;
											assign node541 = (inp[5]) ? 3'b101 : 3'b001;
				assign node545 = (inp[7]) ? node675 : node546;
					assign node546 = (inp[10]) ? node616 : node547;
						assign node547 = (inp[1]) ? node579 : node548;
							assign node548 = (inp[8]) ? node564 : node549;
								assign node549 = (inp[11]) ? node557 : node550;
									assign node550 = (inp[2]) ? node552 : 3'b001;
										assign node552 = (inp[3]) ? 3'b110 : node553;
											assign node553 = (inp[4]) ? 3'b110 : 3'b001;
									assign node557 = (inp[2]) ? node559 : 3'b110;
										assign node559 = (inp[3]) ? 3'b010 : node560;
											assign node560 = (inp[5]) ? 3'b010 : 3'b110;
								assign node564 = (inp[11]) ? node572 : node565;
									assign node565 = (inp[2]) ? node567 : 3'b101;
										assign node567 = (inp[3]) ? 3'b001 : node568;
											assign node568 = (inp[4]) ? 3'b001 : 3'b101;
									assign node572 = (inp[2]) ? node574 : 3'b001;
										assign node574 = (inp[3]) ? 3'b110 : node575;
											assign node575 = (inp[4]) ? 3'b101 : 3'b001;
							assign node579 = (inp[8]) ? node597 : node580;
								assign node580 = (inp[11]) ? node586 : node581;
									assign node581 = (inp[2]) ? 3'b010 : node582;
										assign node582 = (inp[4]) ? 3'b010 : 3'b110;
									assign node586 = (inp[2]) ? node592 : node587;
										assign node587 = (inp[3]) ? node589 : 3'b010;
											assign node589 = (inp[5]) ? 3'b100 : 3'b010;
										assign node592 = (inp[4]) ? node594 : 3'b100;
											assign node594 = (inp[5]) ? 3'b100 : 3'b010;
								assign node597 = (inp[2]) ? node609 : node598;
									assign node598 = (inp[11]) ? node604 : node599;
										assign node599 = (inp[4]) ? node601 : 3'b001;
											assign node601 = (inp[3]) ? 3'b110 : 3'b001;
										assign node604 = (inp[4]) ? node606 : 3'b110;
											assign node606 = (inp[3]) ? 3'b010 : 3'b110;
									assign node609 = (inp[11]) ? node611 : 3'b110;
										assign node611 = (inp[4]) ? node613 : 3'b110;
											assign node613 = (inp[5]) ? 3'b010 : 3'b001;
						assign node616 = (inp[11]) ? node648 : node617;
							assign node617 = (inp[1]) ? node633 : node618;
								assign node618 = (inp[8]) ? node626 : node619;
									assign node619 = (inp[2]) ? node621 : 3'b010;
										assign node621 = (inp[4]) ? 3'b100 : node622;
											assign node622 = (inp[3]) ? 3'b100 : 3'b010;
									assign node626 = (inp[2]) ? node628 : 3'b110;
										assign node628 = (inp[4]) ? 3'b010 : node629;
											assign node629 = (inp[3]) ? 3'b010 : 3'b110;
								assign node633 = (inp[8]) ? node641 : node634;
									assign node634 = (inp[4]) ? node636 : 3'b100;
										assign node636 = (inp[2]) ? 3'b000 : node637;
											assign node637 = (inp[3]) ? 3'b000 : 3'b100;
									assign node641 = (inp[2]) ? node643 : 3'b010;
										assign node643 = (inp[4]) ? 3'b100 : node644;
											assign node644 = (inp[3]) ? 3'b100 : 3'b110;
							assign node648 = (inp[2]) ? node666 : node649;
								assign node649 = (inp[1]) ? node661 : node650;
									assign node650 = (inp[8]) ? node656 : node651;
										assign node651 = (inp[3]) ? 3'b100 : node652;
											assign node652 = (inp[4]) ? 3'b100 : 3'b000;
										assign node656 = (inp[3]) ? 3'b010 : node657;
											assign node657 = (inp[4]) ? 3'b010 : 3'b110;
									assign node661 = (inp[8]) ? 3'b100 : node662;
										assign node662 = (inp[4]) ? 3'b000 : 3'b100;
								assign node666 = (inp[1]) ? node670 : node667;
									assign node667 = (inp[8]) ? 3'b100 : 3'b000;
									assign node670 = (inp[8]) ? 3'b000 : node671;
										assign node671 = (inp[4]) ? 3'b000 : 3'b100;
					assign node675 = (inp[10]) ? node735 : node676;
						assign node676 = (inp[1]) ? node714 : node677;
							assign node677 = (inp[8]) ? node701 : node678;
								assign node678 = (inp[11]) ? node690 : node679;
									assign node679 = (inp[2]) ? node685 : node680;
										assign node680 = (inp[4]) ? 3'b011 : node681;
											assign node681 = (inp[3]) ? 3'b011 : 3'b101;
										assign node685 = (inp[3]) ? 3'b101 : node686;
											assign node686 = (inp[4]) ? 3'b101 : 3'b111;
									assign node690 = (inp[2]) ? node696 : node691;
										assign node691 = (inp[3]) ? 3'b101 : node692;
											assign node692 = (inp[4]) ? 3'b101 : 3'b011;
										assign node696 = (inp[5]) ? 3'b001 : node697;
											assign node697 = (inp[3]) ? 3'b001 : 3'b101;
								assign node701 = (inp[4]) ? node707 : node702;
									assign node702 = (inp[2]) ? 3'b011 : node703;
										assign node703 = (inp[11]) ? 3'b011 : 3'b111;
									assign node707 = (inp[11]) ? node711 : node708;
										assign node708 = (inp[2]) ? 3'b011 : 3'b111;
										assign node711 = (inp[2]) ? 3'b101 : 3'b011;
							assign node714 = (inp[8]) ? node728 : node715;
								assign node715 = (inp[11]) ? node719 : node716;
									assign node716 = (inp[2]) ? 3'b001 : 3'b101;
									assign node719 = (inp[2]) ? node721 : 3'b001;
										assign node721 = (inp[5]) ? node723 : 3'b111;
											assign node723 = (inp[4]) ? node725 : 3'b111;
												assign node725 = (inp[3]) ? 3'b110 : 3'b111;
								assign node728 = (inp[2]) ? node732 : node729;
									assign node729 = (inp[11]) ? 3'b101 : 3'b011;
									assign node732 = (inp[11]) ? 3'b001 : 3'b101;
						assign node735 = (inp[1]) ? node777 : node736;
							assign node736 = (inp[2]) ? node760 : node737;
								assign node737 = (inp[4]) ? node749 : node738;
									assign node738 = (inp[11]) ? node744 : node739;
										assign node739 = (inp[8]) ? 3'b101 : node740;
											assign node740 = (inp[3]) ? 3'b001 : 3'b101;
										assign node744 = (inp[3]) ? node746 : 3'b001;
											assign node746 = (inp[8]) ? 3'b001 : 3'b101;
									assign node749 = (inp[8]) ? node755 : node750;
										assign node750 = (inp[11]) ? node752 : 3'b001;
											assign node752 = (inp[5]) ? 3'b110 : 3'b101;
										assign node755 = (inp[3]) ? node757 : 3'b101;
											assign node757 = (inp[11]) ? 3'b001 : 3'b101;
								assign node760 = (inp[4]) ? node768 : node761;
									assign node761 = (inp[8]) ? node765 : node762;
										assign node762 = (inp[11]) ? 3'b101 : 3'b001;
										assign node765 = (inp[11]) ? 3'b010 : 3'b101;
									assign node768 = (inp[11]) ? node774 : node769;
										assign node769 = (inp[8]) ? node771 : 3'b110;
											assign node771 = (inp[3]) ? 3'b001 : 3'b101;
										assign node774 = (inp[8]) ? 3'b110 : 3'b010;
							assign node777 = (inp[8]) ? node785 : node778;
								assign node778 = (inp[11]) ? node782 : node779;
									assign node779 = (inp[2]) ? 3'b010 : 3'b110;
									assign node782 = (inp[2]) ? 3'b100 : 3'b010;
								assign node785 = (inp[11]) ? node797 : node786;
									assign node786 = (inp[2]) ? node792 : node787;
										assign node787 = (inp[3]) ? 3'b001 : node788;
											assign node788 = (inp[4]) ? 3'b001 : 3'b000;
										assign node792 = (inp[4]) ? node794 : 3'b111;
											assign node794 = (inp[3]) ? 3'b110 : 3'b111;
									assign node797 = (inp[2]) ? 3'b010 : node798;
										assign node798 = (inp[4]) ? 3'b110 : node799;
											assign node799 = (inp[3]) ? 3'b110 : 3'b111;
			assign node804 = (inp[0]) ? node1100 : node805;
				assign node805 = (inp[7]) ? node945 : node806;
					assign node806 = (inp[10]) ? node886 : node807;
						assign node807 = (inp[11]) ? node851 : node808;
							assign node808 = (inp[8]) ? node832 : node809;
								assign node809 = (inp[1]) ? node817 : node810;
									assign node810 = (inp[2]) ? 3'b010 : node811;
										assign node811 = (inp[3]) ? node813 : 3'b110;
											assign node813 = (inp[4]) ? 3'b010 : 3'b110;
									assign node817 = (inp[2]) ? node825 : node818;
										assign node818 = (inp[4]) ? node822 : node819;
											assign node819 = (inp[3]) ? 3'b100 : 3'b010;
											assign node822 = (inp[5]) ? 3'b100 : 3'b000;
										assign node825 = (inp[5]) ? node827 : 3'b100;
											assign node827 = (inp[4]) ? node829 : 3'b100;
												assign node829 = (inp[3]) ? 3'b000 : 3'b100;
								assign node832 = (inp[1]) ? node846 : node833;
									assign node833 = (inp[2]) ? node841 : node834;
										assign node834 = (inp[4]) ? node836 : 3'b001;
											assign node836 = (inp[3]) ? 3'b110 : node837;
												assign node837 = (inp[5]) ? 3'b010 : 3'b110;
										assign node841 = (inp[4]) ? node843 : 3'b110;
											assign node843 = (inp[5]) ? 3'b110 : 3'b010;
									assign node846 = (inp[2]) ? 3'b010 : node847;
										assign node847 = (inp[3]) ? 3'b010 : 3'b110;
							assign node851 = (inp[8]) ? node871 : node852;
								assign node852 = (inp[1]) ? node860 : node853;
									assign node853 = (inp[2]) ? 3'b100 : node854;
										assign node854 = (inp[3]) ? node856 : 3'b000;
											assign node856 = (inp[4]) ? 3'b100 : 3'b000;
									assign node860 = (inp[2]) ? 3'b000 : node861;
										assign node861 = (inp[5]) ? node865 : node862;
											assign node862 = (inp[4]) ? 3'b100 : 3'b000;
											assign node865 = (inp[3]) ? 3'b000 : node866;
												assign node866 = (inp[4]) ? 3'b000 : 3'b100;
								assign node871 = (inp[1]) ? node881 : node872;
									assign node872 = (inp[2]) ? 3'b010 : node873;
										assign node873 = (inp[4]) ? node875 : 3'b101;
											assign node875 = (inp[3]) ? node877 : 3'b110;
												assign node877 = (inp[5]) ? 3'b010 : 3'b110;
									assign node881 = (inp[2]) ? 3'b100 : node882;
										assign node882 = (inp[3]) ? 3'b100 : 3'b010;
						assign node886 = (inp[1]) ? node934 : node887;
							assign node887 = (inp[8]) ? node923 : node888;
								assign node888 = (inp[4]) ? node916 : node889;
									assign node889 = (inp[3]) ? node901 : node890;
										assign node890 = (inp[5]) ? node896 : node891;
											assign node891 = (inp[11]) ? 3'b000 : node892;
												assign node892 = (inp[2]) ? 3'b000 : 3'b100;
											assign node896 = (inp[2]) ? node898 : 3'b000;
												assign node898 = (inp[11]) ? 3'b100 : 3'b000;
										assign node901 = (inp[5]) ? node909 : node902;
											assign node902 = (inp[11]) ? node906 : node903;
												assign node903 = (inp[2]) ? 3'b000 : 3'b100;
												assign node906 = (inp[2]) ? 3'b100 : 3'b000;
											assign node909 = (inp[2]) ? node913 : node910;
												assign node910 = (inp[11]) ? 3'b000 : 3'b100;
												assign node913 = (inp[11]) ? 3'b100 : 3'b000;
									assign node916 = (inp[11]) ? node920 : node917;
										assign node917 = (inp[2]) ? 3'b000 : 3'b100;
										assign node920 = (inp[2]) ? 3'b100 : 3'b000;
								assign node923 = (inp[11]) ? node931 : node924;
									assign node924 = (inp[2]) ? node926 : 3'b010;
										assign node926 = (inp[3]) ? 3'b100 : node927;
											assign node927 = (inp[4]) ? 3'b100 : 3'b110;
									assign node931 = (inp[2]) ? 3'b000 : 3'b100;
							assign node934 = (inp[4]) ? node936 : 3'b000;
								assign node936 = (inp[8]) ? node938 : 3'b000;
									assign node938 = (inp[11]) ? 3'b000 : node939;
										assign node939 = (inp[3]) ? 3'b000 : node940;
											assign node940 = (inp[2]) ? 3'b000 : 3'b100;
					assign node945 = (inp[10]) ? node1041 : node946;
						assign node946 = (inp[1]) ? node992 : node947;
							assign node947 = (inp[8]) ? node977 : node948;
								assign node948 = (inp[2]) ? node968 : node949;
									assign node949 = (inp[3]) ? node957 : node950;
										assign node950 = (inp[5]) ? node952 : 3'b101;
											assign node952 = (inp[11]) ? node954 : 3'b101;
												assign node954 = (inp[4]) ? 3'b001 : 3'b101;
										assign node957 = (inp[5]) ? node963 : node958;
											assign node958 = (inp[4]) ? 3'b101 : node959;
												assign node959 = (inp[11]) ? 3'b001 : 3'b101;
											assign node963 = (inp[11]) ? 3'b001 : node964;
												assign node964 = (inp[4]) ? 3'b001 : 3'b101;
									assign node968 = (inp[11]) ? 3'b110 : node969;
										assign node969 = (inp[3]) ? 3'b001 : node970;
											assign node970 = (inp[5]) ? node972 : 3'b101;
												assign node972 = (inp[4]) ? 3'b001 : 3'b101;
								assign node977 = (inp[11]) ? node985 : node978;
									assign node978 = (inp[2]) ? node980 : 3'b011;
										assign node980 = (inp[3]) ? 3'b101 : node981;
											assign node981 = (inp[5]) ? 3'b011 : 3'b101;
									assign node985 = (inp[2]) ? 3'b001 : node986;
										assign node986 = (inp[4]) ? 3'b101 : node987;
											assign node987 = (inp[3]) ? 3'b101 : 3'b001;
							assign node992 = (inp[11]) ? node1010 : node993;
								assign node993 = (inp[8]) ? node1003 : node994;
									assign node994 = (inp[2]) ? 3'b110 : node995;
										assign node995 = (inp[5]) ? node997 : 3'b001;
											assign node997 = (inp[4]) ? node999 : 3'b110;
												assign node999 = (inp[3]) ? 3'b110 : 3'b001;
									assign node1003 = (inp[2]) ? 3'b001 : node1004;
										assign node1004 = (inp[3]) ? node1006 : 3'b101;
											assign node1006 = (inp[4]) ? 3'b001 : 3'b101;
								assign node1010 = (inp[5]) ? node1024 : node1011;
									assign node1011 = (inp[2]) ? node1019 : node1012;
										assign node1012 = (inp[8]) ? node1014 : 3'b110;
											assign node1014 = (inp[3]) ? node1016 : 3'b010;
												assign node1016 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1019 = (inp[8]) ? 3'b110 : node1020;
											assign node1020 = (inp[4]) ? 3'b010 : 3'b001;
									assign node1024 = (inp[2]) ? node1036 : node1025;
										assign node1025 = (inp[8]) ? node1031 : node1026;
											assign node1026 = (inp[4]) ? node1028 : 3'b110;
												assign node1028 = (inp[3]) ? 3'b010 : 3'b110;
											assign node1031 = (inp[3]) ? node1033 : 3'b010;
												assign node1033 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1036 = (inp[4]) ? node1038 : 3'b110;
											assign node1038 = (inp[8]) ? 3'b110 : 3'b010;
						assign node1041 = (inp[1]) ? node1061 : node1042;
							assign node1042 = (inp[11]) ? node1054 : node1043;
								assign node1043 = (inp[2]) ? node1047 : node1044;
									assign node1044 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1047 = (inp[8]) ? node1049 : 3'b010;
										assign node1049 = (inp[3]) ? 3'b110 : node1050;
											assign node1050 = (inp[4]) ? 3'b110 : 3'b111;
								assign node1054 = (inp[2]) ? node1058 : node1055;
									assign node1055 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1058 = (inp[8]) ? 3'b010 : 3'b100;
							assign node1061 = (inp[8]) ? node1077 : node1062;
								assign node1062 = (inp[11]) ? node1070 : node1063;
									assign node1063 = (inp[2]) ? 3'b100 : node1064;
										assign node1064 = (inp[3]) ? node1066 : 3'b010;
											assign node1066 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1070 = (inp[2]) ? 3'b000 : node1071;
										assign node1071 = (inp[4]) ? node1073 : 3'b100;
											assign node1073 = (inp[3]) ? 3'b000 : 3'b100;
								assign node1077 = (inp[2]) ? node1093 : node1078;
									assign node1078 = (inp[11]) ? node1086 : node1079;
										assign node1079 = (inp[4]) ? node1081 : 3'b100;
											assign node1081 = (inp[5]) ? node1083 : 3'b010;
												assign node1083 = (inp[3]) ? 3'b010 : 3'b110;
										assign node1086 = (inp[3]) ? node1088 : 3'b010;
											assign node1088 = (inp[4]) ? node1090 : 3'b010;
												assign node1090 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1093 = (inp[11]) ? 3'b100 : node1094;
										assign node1094 = (inp[5]) ? 3'b010 : node1095;
											assign node1095 = (inp[4]) ? 3'b100 : 3'b010;
				assign node1100 = (inp[10]) ? node1180 : node1101;
					assign node1101 = (inp[7]) ? node1125 : node1102;
						assign node1102 = (inp[1]) ? 3'b000 : node1103;
							assign node1103 = (inp[8]) ? node1105 : 3'b000;
								assign node1105 = (inp[11]) ? node1117 : node1106;
									assign node1106 = (inp[2]) ? node1112 : node1107;
										assign node1107 = (inp[3]) ? 3'b100 : node1108;
											assign node1108 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1112 = (inp[4]) ? node1114 : 3'b100;
											assign node1114 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1117 = (inp[4]) ? 3'b000 : node1118;
										assign node1118 = (inp[2]) ? 3'b010 : node1119;
											assign node1119 = (inp[3]) ? 3'b010 : 3'b100;
						assign node1125 = (inp[1]) ? node1153 : node1126;
							assign node1126 = (inp[8]) ? node1140 : node1127;
								assign node1127 = (inp[4]) ? node1129 : 3'b010;
									assign node1129 = (inp[2]) ? node1135 : node1130;
										assign node1130 = (inp[5]) ? node1132 : 3'b010;
											assign node1132 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1135 = (inp[3]) ? 3'b000 : node1136;
											assign node1136 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1140 = (inp[4]) ? node1146 : node1141;
									assign node1141 = (inp[11]) ? node1143 : 3'b110;
										assign node1143 = (inp[2]) ? 3'b100 : 3'b110;
									assign node1146 = (inp[11]) ? node1150 : node1147;
										assign node1147 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1150 = (inp[2]) ? 3'b100 : 3'b010;
							assign node1153 = (inp[8]) ? node1161 : node1154;
								assign node1154 = (inp[11]) ? node1158 : node1155;
									assign node1155 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1158 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1161 = (inp[11]) ? node1173 : node1162;
									assign node1162 = (inp[2]) ? node1168 : node1163;
										assign node1163 = (inp[3]) ? 3'b010 : node1164;
											assign node1164 = (inp[4]) ? 3'b010 : 3'b000;
										assign node1168 = (inp[4]) ? node1170 : 3'b110;
											assign node1170 = (inp[3]) ? 3'b100 : 3'b110;
									assign node1173 = (inp[2]) ? 3'b000 : node1174;
										assign node1174 = (inp[3]) ? 3'b100 : node1175;
											assign node1175 = (inp[4]) ? 3'b100 : 3'b110;
					assign node1180 = (inp[1]) ? 3'b000 : node1181;
						assign node1181 = (inp[7]) ? node1183 : 3'b000;
							assign node1183 = (inp[8]) ? node1185 : 3'b000;
								assign node1185 = (inp[11]) ? node1193 : node1186;
									assign node1186 = (inp[2]) ? 3'b100 : node1187;
										assign node1187 = (inp[3]) ? 3'b100 : node1188;
											assign node1188 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1193 = (inp[3]) ? 3'b000 : node1194;
										assign node1194 = (inp[2]) ? 3'b000 : 3'b100;

endmodule