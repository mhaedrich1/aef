module dtc_split5_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;

	assign outp = (inp[9]) ? node208 : node1;
		assign node1 = (inp[6]) ? node127 : node2;
			assign node2 = (inp[10]) ? node48 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[3]) ? node8 : 3'b111;
							assign node8 = (inp[11]) ? 3'b011 : 3'b111;
					assign node11 = (inp[11]) ? node27 : node12;
						assign node12 = (inp[3]) ? node20 : node13;
							assign node13 = (inp[1]) ? node15 : 3'b111;
								assign node15 = (inp[8]) ? node17 : 3'b111;
									assign node17 = (inp[2]) ? 3'b111 : 3'b011;
							assign node20 = (inp[8]) ? 3'b011 : node21;
								assign node21 = (inp[5]) ? node23 : 3'b111;
									assign node23 = (inp[4]) ? 3'b011 : 3'b111;
						assign node27 = (inp[3]) ? node41 : node28;
							assign node28 = (inp[1]) ? node36 : node29;
								assign node29 = (inp[8]) ? 3'b011 : node30;
									assign node30 = (inp[4]) ? 3'b011 : node31;
										assign node31 = (inp[2]) ? 3'b011 : 3'b111;
								assign node36 = (inp[2]) ? 3'b011 : node37;
									assign node37 = (inp[8]) ? 3'b001 : 3'b011;
							assign node41 = (inp[8]) ? 3'b101 : node42;
								assign node42 = (inp[4]) ? node44 : 3'b011;
									assign node44 = (inp[5]) ? 3'b101 : 3'b111;
				assign node48 = (inp[11]) ? node98 : node49;
					assign node49 = (inp[8]) ? node71 : node50;
						assign node50 = (inp[3]) ? node60 : node51;
							assign node51 = (inp[4]) ? node57 : node52;
								assign node52 = (inp[2]) ? 3'b111 : node53;
									assign node53 = (inp[7]) ? 3'b011 : 3'b111;
								assign node57 = (inp[7]) ? 3'b101 : 3'b111;
							assign node60 = (inp[4]) ? node68 : node61;
								assign node61 = (inp[7]) ? 3'b111 : node62;
									assign node62 = (inp[2]) ? 3'b011 : node63;
										assign node63 = (inp[1]) ? 3'b011 : 3'b111;
								assign node68 = (inp[7]) ? 3'b001 : 3'b011;
						assign node71 = (inp[3]) ? node87 : node72;
							assign node72 = (inp[7]) ? node74 : 3'b011;
								assign node74 = (inp[2]) ? node82 : node75;
									assign node75 = (inp[4]) ? node77 : 3'b101;
										assign node77 = (inp[0]) ? 3'b010 : node78;
											assign node78 = (inp[5]) ? 3'b001 : 3'b101;
									assign node82 = (inp[0]) ? node84 : 3'b001;
										assign node84 = (inp[5]) ? 3'b010 : 3'b001;
							assign node87 = (inp[7]) ? node91 : node88;
								assign node88 = (inp[4]) ? 3'b101 : 3'b001;
								assign node91 = (inp[1]) ? node93 : 3'b001;
									assign node93 = (inp[0]) ? node95 : 3'b001;
										assign node95 = (inp[2]) ? 3'b001 : 3'b110;
					assign node98 = (inp[7]) ? node108 : node99;
						assign node99 = (inp[3]) ? node103 : node100;
							assign node100 = (inp[8]) ? 3'b101 : 3'b011;
							assign node103 = (inp[8]) ? node105 : 3'b101;
								assign node105 = (inp[4]) ? 3'b001 : 3'b101;
						assign node108 = (inp[8]) ? node116 : node109;
							assign node109 = (inp[4]) ? node111 : 3'b101;
								assign node111 = (inp[3]) ? node113 : 3'b101;
									assign node113 = (inp[5]) ? 3'b110 : 3'b101;
							assign node116 = (inp[3]) ? node122 : node117;
								assign node117 = (inp[2]) ? 3'b101 : node118;
									assign node118 = (inp[1]) ? 3'b110 : 3'b101;
								assign node122 = (inp[5]) ? node124 : 3'b110;
									assign node124 = (inp[4]) ? 3'b010 : 3'b110;
			assign node127 = (inp[10]) ? node187 : node128;
				assign node128 = (inp[11]) ? node168 : node129;
					assign node129 = (inp[7]) ? node147 : node130;
						assign node130 = (inp[8]) ? node136 : node131;
							assign node131 = (inp[4]) ? node133 : 3'b011;
								assign node133 = (inp[3]) ? 3'b101 : 3'b011;
							assign node136 = (inp[5]) ? node140 : node137;
								assign node137 = (inp[4]) ? 3'b001 : 3'b011;
								assign node140 = (inp[1]) ? 3'b001 : node141;
									assign node141 = (inp[2]) ? 3'b001 : node142;
										assign node142 = (inp[0]) ? 3'b001 : 3'b101;
						assign node147 = (inp[4]) ? node157 : node148;
							assign node148 = (inp[8]) ? node154 : node149;
								assign node149 = (inp[3]) ? 3'b001 : node150;
									assign node150 = (inp[2]) ? 3'b001 : 3'b101;
								assign node154 = (inp[3]) ? 3'b110 : 3'b001;
							assign node157 = (inp[3]) ? node161 : node158;
								assign node158 = (inp[8]) ? 3'b110 : 3'b001;
								assign node161 = (inp[8]) ? node163 : 3'b110;
									assign node163 = (inp[0]) ? node165 : 3'b110;
										assign node165 = (inp[5]) ? 3'b010 : 3'b110;
					assign node168 = (inp[8]) ? node176 : node169;
						assign node169 = (inp[7]) ? node171 : 3'b001;
							assign node171 = (inp[4]) ? node173 : 3'b110;
								assign node173 = (inp[3]) ? 3'b010 : 3'b110;
						assign node176 = (inp[7]) ? node178 : 3'b110;
							assign node178 = (inp[4]) ? node180 : 3'b010;
								assign node180 = (inp[0]) ? node182 : 3'b010;
									assign node182 = (inp[5]) ? node184 : 3'b010;
										assign node184 = (inp[3]) ? 3'b100 : 3'b010;
				assign node187 = (inp[7]) ? node195 : node188;
					assign node188 = (inp[8]) ? node192 : node189;
						assign node189 = (inp[11]) ? 3'b010 : 3'b110;
						assign node192 = (inp[11]) ? 3'b100 : 3'b010;
					assign node195 = (inp[11]) ? 3'b000 : node196;
						assign node196 = (inp[5]) ? node198 : 3'b100;
							assign node198 = (inp[8]) ? node200 : 3'b100;
								assign node200 = (inp[2]) ? node202 : 3'b100;
									assign node202 = (inp[4]) ? node204 : 3'b100;
										assign node204 = (inp[3]) ? 3'b000 : 3'b100;
		assign node208 = (inp[6]) ? node272 : node209;
			assign node209 = (inp[10]) ? node257 : node210;
				assign node210 = (inp[8]) ? node232 : node211;
					assign node211 = (inp[7]) ? node229 : node212;
						assign node212 = (inp[3]) ? node218 : node213;
							assign node213 = (inp[4]) ? 3'b101 : node214;
								assign node214 = (inp[11]) ? 3'b001 : 3'b101;
							assign node218 = (inp[11]) ? node226 : node219;
								assign node219 = (inp[2]) ? 3'b001 : node220;
									assign node220 = (inp[5]) ? node222 : 3'b101;
										assign node222 = (inp[0]) ? 3'b001 : 3'b101;
								assign node226 = (inp[4]) ? 3'b110 : 3'b001;
						assign node229 = (inp[11]) ? 3'b100 : 3'b010;
					assign node232 = (inp[7]) ? node244 : node233;
						assign node233 = (inp[11]) ? node235 : 3'b000;
							assign node235 = (inp[0]) ? node237 : 3'b010;
								assign node237 = (inp[5]) ? node239 : 3'b010;
									assign node239 = (inp[4]) ? node241 : 3'b010;
										assign node241 = (inp[3]) ? 3'b101 : 3'b110;
						assign node244 = (inp[11]) ? node254 : node245;
							assign node245 = (inp[3]) ? node247 : 3'b010;
								assign node247 = (inp[2]) ? 3'b100 : node248;
									assign node248 = (inp[0]) ? node250 : 3'b010;
										assign node250 = (inp[5]) ? 3'b100 : 3'b010;
							assign node254 = (inp[4]) ? 3'b000 : 3'b100;
				assign node257 = (inp[7]) ? 3'b000 : node258;
					assign node258 = (inp[11]) ? node262 : node259;
						assign node259 = (inp[8]) ? 3'b100 : 3'b010;
						assign node262 = (inp[8]) ? 3'b000 : node263;
							assign node263 = (inp[5]) ? node265 : 3'b100;
								assign node265 = (inp[4]) ? node267 : 3'b100;
									assign node267 = (inp[0]) ? 3'b000 : 3'b100;
			assign node272 = (inp[10]) ? 3'b000 : node273;
				assign node273 = (inp[11]) ? 3'b000 : node274;
					assign node274 = (inp[7]) ? 3'b000 : node275;
						assign node275 = (inp[8]) ? 3'b000 : 3'b100;

endmodule