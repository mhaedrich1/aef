module dtc_split5_bm23 (
	input  wire [12-1:0] inp,
	output wire [12-1:0] outp
);

	wire [12-1:0] node1;
	wire [12-1:0] node2;
	wire [12-1:0] node3;
	wire [12-1:0] node4;
	wire [12-1:0] node5;
	wire [12-1:0] node6;
	wire [12-1:0] node7;
	wire [12-1:0] node8;
	wire [12-1:0] node9;
	wire [12-1:0] node11;
	wire [12-1:0] node12;
	wire [12-1:0] node16;
	wire [12-1:0] node19;
	wire [12-1:0] node20;
	wire [12-1:0] node21;
	wire [12-1:0] node22;
	wire [12-1:0] node27;
	wire [12-1:0] node28;
	wire [12-1:0] node30;
	wire [12-1:0] node34;
	wire [12-1:0] node35;
	wire [12-1:0] node36;
	wire [12-1:0] node39;
	wire [12-1:0] node40;
	wire [12-1:0] node41;
	wire [12-1:0] node45;
	wire [12-1:0] node46;
	wire [12-1:0] node50;
	wire [12-1:0] node51;
	wire [12-1:0] node53;
	wire [12-1:0] node54;
	wire [12-1:0] node59;
	wire [12-1:0] node60;
	wire [12-1:0] node61;
	wire [12-1:0] node62;
	wire [12-1:0] node63;
	wire [12-1:0] node67;
	wire [12-1:0] node69;
	wire [12-1:0] node72;
	wire [12-1:0] node73;
	wire [12-1:0] node75;
	wire [12-1:0] node76;
	wire [12-1:0] node80;
	wire [12-1:0] node83;
	wire [12-1:0] node84;
	wire [12-1:0] node85;
	wire [12-1:0] node87;
	wire [12-1:0] node90;
	wire [12-1:0] node91;
	wire [12-1:0] node95;
	wire [12-1:0] node97;
	wire [12-1:0] node98;
	wire [12-1:0] node99;
	wire [12-1:0] node103;
	wire [12-1:0] node106;
	wire [12-1:0] node107;
	wire [12-1:0] node108;
	wire [12-1:0] node109;
	wire [12-1:0] node110;
	wire [12-1:0] node111;
	wire [12-1:0] node112;
	wire [12-1:0] node116;
	wire [12-1:0] node119;
	wire [12-1:0] node120;
	wire [12-1:0] node123;
	wire [12-1:0] node124;
	wire [12-1:0] node128;
	wire [12-1:0] node129;
	wire [12-1:0] node130;
	wire [12-1:0] node131;
	wire [12-1:0] node135;
	wire [12-1:0] node136;
	wire [12-1:0] node140;
	wire [12-1:0] node141;
	wire [12-1:0] node143;
	wire [12-1:0] node147;
	wire [12-1:0] node148;
	wire [12-1:0] node149;
	wire [12-1:0] node150;
	wire [12-1:0] node154;
	wire [12-1:0] node157;
	wire [12-1:0] node158;
	wire [12-1:0] node161;
	wire [12-1:0] node162;
	wire [12-1:0] node165;
	wire [12-1:0] node167;
	wire [12-1:0] node170;
	wire [12-1:0] node171;
	wire [12-1:0] node172;
	wire [12-1:0] node173;
	wire [12-1:0] node176;
	wire [12-1:0] node178;
	wire [12-1:0] node181;
	wire [12-1:0] node182;
	wire [12-1:0] node185;
	wire [12-1:0] node188;
	wire [12-1:0] node189;
	wire [12-1:0] node190;
	wire [12-1:0] node194;
	wire [12-1:0] node195;
	wire [12-1:0] node197;
	wire [12-1:0] node198;
	wire [12-1:0] node202;
	wire [12-1:0] node205;
	wire [12-1:0] node206;
	wire [12-1:0] node207;
	wire [12-1:0] node208;
	wire [12-1:0] node209;
	wire [12-1:0] node210;
	wire [12-1:0] node212;
	wire [12-1:0] node215;
	wire [12-1:0] node218;
	wire [12-1:0] node219;
	wire [12-1:0] node221;
	wire [12-1:0] node222;
	wire [12-1:0] node227;
	wire [12-1:0] node228;
	wire [12-1:0] node229;
	wire [12-1:0] node230;
	wire [12-1:0] node232;
	wire [12-1:0] node235;
	wire [12-1:0] node236;
	wire [12-1:0] node240;
	wire [12-1:0] node241;
	wire [12-1:0] node243;
	wire [12-1:0] node247;
	wire [12-1:0] node248;
	wire [12-1:0] node250;
	wire [12-1:0] node253;
	wire [12-1:0] node254;
	wire [12-1:0] node255;
	wire [12-1:0] node259;
	wire [12-1:0] node262;
	wire [12-1:0] node263;
	wire [12-1:0] node264;
	wire [12-1:0] node265;
	wire [12-1:0] node266;
	wire [12-1:0] node268;
	wire [12-1:0] node271;
	wire [12-1:0] node274;
	wire [12-1:0] node276;
	wire [12-1:0] node279;
	wire [12-1:0] node280;
	wire [12-1:0] node282;
	wire [12-1:0] node285;
	wire [12-1:0] node287;
	wire [12-1:0] node290;
	wire [12-1:0] node291;
	wire [12-1:0] node292;
	wire [12-1:0] node295;
	wire [12-1:0] node296;
	wire [12-1:0] node300;
	wire [12-1:0] node301;
	wire [12-1:0] node304;
	wire [12-1:0] node305;
	wire [12-1:0] node309;
	wire [12-1:0] node310;
	wire [12-1:0] node311;
	wire [12-1:0] node312;
	wire [12-1:0] node313;
	wire [12-1:0] node315;
	wire [12-1:0] node316;
	wire [12-1:0] node320;
	wire [12-1:0] node321;
	wire [12-1:0] node322;
	wire [12-1:0] node325;
	wire [12-1:0] node329;
	wire [12-1:0] node330;
	wire [12-1:0] node332;
	wire [12-1:0] node333;
	wire [12-1:0] node338;
	wire [12-1:0] node339;
	wire [12-1:0] node340;
	wire [12-1:0] node344;
	wire [12-1:0] node345;
	wire [12-1:0] node346;
	wire [12-1:0] node348;
	wire [12-1:0] node352;
	wire [12-1:0] node355;
	wire [12-1:0] node356;
	wire [12-1:0] node357;
	wire [12-1:0] node358;
	wire [12-1:0] node359;
	wire [12-1:0] node360;
	wire [12-1:0] node365;
	wire [12-1:0] node368;
	wire [12-1:0] node369;
	wire [12-1:0] node370;
	wire [12-1:0] node373;
	wire [12-1:0] node374;
	wire [12-1:0] node378;
	wire [12-1:0] node380;
	wire [12-1:0] node382;
	wire [12-1:0] node385;
	wire [12-1:0] node386;
	wire [12-1:0] node387;
	wire [12-1:0] node390;
	wire [12-1:0] node392;
	wire [12-1:0] node393;
	wire [12-1:0] node397;
	wire [12-1:0] node398;
	wire [12-1:0] node400;
	wire [12-1:0] node401;
	wire [12-1:0] node405;
	wire [12-1:0] node406;
	wire [12-1:0] node410;
	wire [12-1:0] node411;
	wire [12-1:0] node412;
	wire [12-1:0] node413;
	wire [12-1:0] node414;
	wire [12-1:0] node415;
	wire [12-1:0] node416;
	wire [12-1:0] node418;
	wire [12-1:0] node419;
	wire [12-1:0] node424;
	wire [12-1:0] node425;
	wire [12-1:0] node426;
	wire [12-1:0] node427;
	wire [12-1:0] node432;
	wire [12-1:0] node435;
	wire [12-1:0] node436;
	wire [12-1:0] node437;
	wire [12-1:0] node439;
	wire [12-1:0] node442;
	wire [12-1:0] node443;
	wire [12-1:0] node444;
	wire [12-1:0] node447;
	wire [12-1:0] node450;
	wire [12-1:0] node451;
	wire [12-1:0] node455;
	wire [12-1:0] node456;
	wire [12-1:0] node457;
	wire [12-1:0] node459;
	wire [12-1:0] node463;
	wire [12-1:0] node466;
	wire [12-1:0] node467;
	wire [12-1:0] node468;
	wire [12-1:0] node469;
	wire [12-1:0] node470;
	wire [12-1:0] node472;
	wire [12-1:0] node476;
	wire [12-1:0] node478;
	wire [12-1:0] node479;
	wire [12-1:0] node483;
	wire [12-1:0] node484;
	wire [12-1:0] node487;
	wire [12-1:0] node489;
	wire [12-1:0] node490;
	wire [12-1:0] node494;
	wire [12-1:0] node495;
	wire [12-1:0] node496;
	wire [12-1:0] node497;
	wire [12-1:0] node501;
	wire [12-1:0] node503;
	wire [12-1:0] node506;
	wire [12-1:0] node507;
	wire [12-1:0] node510;
	wire [12-1:0] node513;
	wire [12-1:0] node514;
	wire [12-1:0] node515;
	wire [12-1:0] node516;
	wire [12-1:0] node517;
	wire [12-1:0] node518;
	wire [12-1:0] node520;
	wire [12-1:0] node524;
	wire [12-1:0] node527;
	wire [12-1:0] node528;
	wire [12-1:0] node531;
	wire [12-1:0] node532;
	wire [12-1:0] node533;
	wire [12-1:0] node537;
	wire [12-1:0] node540;
	wire [12-1:0] node541;
	wire [12-1:0] node542;
	wire [12-1:0] node543;
	wire [12-1:0] node545;
	wire [12-1:0] node548;
	wire [12-1:0] node549;
	wire [12-1:0] node553;
	wire [12-1:0] node556;
	wire [12-1:0] node557;
	wire [12-1:0] node560;
	wire [12-1:0] node562;
	wire [12-1:0] node565;
	wire [12-1:0] node566;
	wire [12-1:0] node567;
	wire [12-1:0] node568;
	wire [12-1:0] node569;
	wire [12-1:0] node573;
	wire [12-1:0] node575;
	wire [12-1:0] node578;
	wire [12-1:0] node579;
	wire [12-1:0] node580;
	wire [12-1:0] node581;
	wire [12-1:0] node585;
	wire [12-1:0] node586;
	wire [12-1:0] node590;
	wire [12-1:0] node592;
	wire [12-1:0] node594;
	wire [12-1:0] node597;
	wire [12-1:0] node598;
	wire [12-1:0] node599;
	wire [12-1:0] node600;
	wire [12-1:0] node604;
	wire [12-1:0] node606;
	wire [12-1:0] node609;
	wire [12-1:0] node610;
	wire [12-1:0] node613;
	wire [12-1:0] node614;
	wire [12-1:0] node616;
	wire [12-1:0] node620;
	wire [12-1:0] node621;
	wire [12-1:0] node622;
	wire [12-1:0] node623;
	wire [12-1:0] node624;
	wire [12-1:0] node625;
	wire [12-1:0] node626;
	wire [12-1:0] node628;
	wire [12-1:0] node631;
	wire [12-1:0] node632;
	wire [12-1:0] node636;
	wire [12-1:0] node638;
	wire [12-1:0] node641;
	wire [12-1:0] node642;
	wire [12-1:0] node643;
	wire [12-1:0] node644;
	wire [12-1:0] node648;
	wire [12-1:0] node649;
	wire [12-1:0] node653;
	wire [12-1:0] node655;
	wire [12-1:0] node656;
	wire [12-1:0] node660;
	wire [12-1:0] node661;
	wire [12-1:0] node662;
	wire [12-1:0] node663;
	wire [12-1:0] node667;
	wire [12-1:0] node669;
	wire [12-1:0] node672;
	wire [12-1:0] node673;
	wire [12-1:0] node674;
	wire [12-1:0] node678;
	wire [12-1:0] node680;
	wire [12-1:0] node683;
	wire [12-1:0] node684;
	wire [12-1:0] node685;
	wire [12-1:0] node686;
	wire [12-1:0] node690;
	wire [12-1:0] node691;
	wire [12-1:0] node692;
	wire [12-1:0] node696;
	wire [12-1:0] node697;
	wire [12-1:0] node698;
	wire [12-1:0] node702;
	wire [12-1:0] node703;
	wire [12-1:0] node707;
	wire [12-1:0] node708;
	wire [12-1:0] node709;
	wire [12-1:0] node710;
	wire [12-1:0] node712;
	wire [12-1:0] node715;
	wire [12-1:0] node716;
	wire [12-1:0] node720;
	wire [12-1:0] node722;
	wire [12-1:0] node725;
	wire [12-1:0] node726;
	wire [12-1:0] node729;
	wire [12-1:0] node732;
	wire [12-1:0] node733;
	wire [12-1:0] node734;
	wire [12-1:0] node735;
	wire [12-1:0] node736;
	wire [12-1:0] node737;
	wire [12-1:0] node738;
	wire [12-1:0] node743;
	wire [12-1:0] node745;
	wire [12-1:0] node748;
	wire [12-1:0] node749;
	wire [12-1:0] node752;
	wire [12-1:0] node753;
	wire [12-1:0] node757;
	wire [12-1:0] node758;
	wire [12-1:0] node759;
	wire [12-1:0] node762;
	wire [12-1:0] node763;
	wire [12-1:0] node765;
	wire [12-1:0] node768;
	wire [12-1:0] node769;
	wire [12-1:0] node773;
	wire [12-1:0] node774;
	wire [12-1:0] node775;
	wire [12-1:0] node777;
	wire [12-1:0] node781;
	wire [12-1:0] node782;
	wire [12-1:0] node786;
	wire [12-1:0] node787;
	wire [12-1:0] node788;
	wire [12-1:0] node789;
	wire [12-1:0] node792;
	wire [12-1:0] node793;
	wire [12-1:0] node795;
	wire [12-1:0] node799;
	wire [12-1:0] node800;
	wire [12-1:0] node801;
	wire [12-1:0] node805;
	wire [12-1:0] node807;
	wire [12-1:0] node809;
	wire [12-1:0] node812;
	wire [12-1:0] node813;
	wire [12-1:0] node814;
	wire [12-1:0] node817;
	wire [12-1:0] node819;
	wire [12-1:0] node822;
	wire [12-1:0] node823;
	wire [12-1:0] node825;
	wire [12-1:0] node826;
	wire [12-1:0] node830;
	wire [12-1:0] node832;
	wire [12-1:0] node835;
	wire [12-1:0] node836;
	wire [12-1:0] node837;
	wire [12-1:0] node838;
	wire [12-1:0] node839;
	wire [12-1:0] node840;
	wire [12-1:0] node841;
	wire [12-1:0] node842;
	wire [12-1:0] node843;
	wire [12-1:0] node847;
	wire [12-1:0] node850;
	wire [12-1:0] node851;
	wire [12-1:0] node852;
	wire [12-1:0] node857;
	wire [12-1:0] node858;
	wire [12-1:0] node859;
	wire [12-1:0] node860;
	wire [12-1:0] node861;
	wire [12-1:0] node865;
	wire [12-1:0] node866;
	wire [12-1:0] node869;
	wire [12-1:0] node872;
	wire [12-1:0] node874;
	wire [12-1:0] node875;
	wire [12-1:0] node879;
	wire [12-1:0] node880;
	wire [12-1:0] node882;
	wire [12-1:0] node885;
	wire [12-1:0] node886;
	wire [12-1:0] node889;
	wire [12-1:0] node890;
	wire [12-1:0] node894;
	wire [12-1:0] node895;
	wire [12-1:0] node896;
	wire [12-1:0] node897;
	wire [12-1:0] node898;
	wire [12-1:0] node900;
	wire [12-1:0] node904;
	wire [12-1:0] node907;
	wire [12-1:0] node908;
	wire [12-1:0] node911;
	wire [12-1:0] node912;
	wire [12-1:0] node913;
	wire [12-1:0] node917;
	wire [12-1:0] node918;
	wire [12-1:0] node922;
	wire [12-1:0] node923;
	wire [12-1:0] node924;
	wire [12-1:0] node926;
	wire [12-1:0] node927;
	wire [12-1:0] node931;
	wire [12-1:0] node933;
	wire [12-1:0] node935;
	wire [12-1:0] node938;
	wire [12-1:0] node939;
	wire [12-1:0] node940;
	wire [12-1:0] node944;
	wire [12-1:0] node947;
	wire [12-1:0] node948;
	wire [12-1:0] node949;
	wire [12-1:0] node950;
	wire [12-1:0] node951;
	wire [12-1:0] node952;
	wire [12-1:0] node953;
	wire [12-1:0] node958;
	wire [12-1:0] node960;
	wire [12-1:0] node961;
	wire [12-1:0] node965;
	wire [12-1:0] node966;
	wire [12-1:0] node967;
	wire [12-1:0] node969;
	wire [12-1:0] node974;
	wire [12-1:0] node975;
	wire [12-1:0] node976;
	wire [12-1:0] node977;
	wire [12-1:0] node979;
	wire [12-1:0] node982;
	wire [12-1:0] node984;
	wire [12-1:0] node987;
	wire [12-1:0] node989;
	wire [12-1:0] node992;
	wire [12-1:0] node993;
	wire [12-1:0] node994;
	wire [12-1:0] node997;
	wire [12-1:0] node998;
	wire [12-1:0] node1002;
	wire [12-1:0] node1003;
	wire [12-1:0] node1005;
	wire [12-1:0] node1009;
	wire [12-1:0] node1010;
	wire [12-1:0] node1011;
	wire [12-1:0] node1012;
	wire [12-1:0] node1013;
	wire [12-1:0] node1015;
	wire [12-1:0] node1019;
	wire [12-1:0] node1020;
	wire [12-1:0] node1022;
	wire [12-1:0] node1027;
	wire [12-1:0] node1028;
	wire [12-1:0] node1029;
	wire [12-1:0] node1030;
	wire [12-1:0] node1034;
	wire [12-1:0] node1036;
	wire [12-1:0] node1039;
	wire [12-1:0] node1040;
	wire [12-1:0] node1041;
	wire [12-1:0] node1044;
	wire [12-1:0] node1045;
	wire [12-1:0] node1049;
	wire [12-1:0] node1051;
	wire [12-1:0] node1053;
	wire [12-1:0] node1056;
	wire [12-1:0] node1057;
	wire [12-1:0] node1058;
	wire [12-1:0] node1059;
	wire [12-1:0] node1060;
	wire [12-1:0] node1061;
	wire [12-1:0] node1062;
	wire [12-1:0] node1064;
	wire [12-1:0] node1067;
	wire [12-1:0] node1068;
	wire [12-1:0] node1072;
	wire [12-1:0] node1075;
	wire [12-1:0] node1076;
	wire [12-1:0] node1080;
	wire [12-1:0] node1081;
	wire [12-1:0] node1082;
	wire [12-1:0] node1083;
	wire [12-1:0] node1084;
	wire [12-1:0] node1089;
	wire [12-1:0] node1091;
	wire [12-1:0] node1094;
	wire [12-1:0] node1095;
	wire [12-1:0] node1096;
	wire [12-1:0] node1097;
	wire [12-1:0] node1100;
	wire [12-1:0] node1104;
	wire [12-1:0] node1105;
	wire [12-1:0] node1107;
	wire [12-1:0] node1111;
	wire [12-1:0] node1112;
	wire [12-1:0] node1113;
	wire [12-1:0] node1114;
	wire [12-1:0] node1116;
	wire [12-1:0] node1120;
	wire [12-1:0] node1121;
	wire [12-1:0] node1122;
	wire [12-1:0] node1123;
	wire [12-1:0] node1128;
	wire [12-1:0] node1129;
	wire [12-1:0] node1131;
	wire [12-1:0] node1135;
	wire [12-1:0] node1136;
	wire [12-1:0] node1137;
	wire [12-1:0] node1140;
	wire [12-1:0] node1142;
	wire [12-1:0] node1143;
	wire [12-1:0] node1147;
	wire [12-1:0] node1148;
	wire [12-1:0] node1149;
	wire [12-1:0] node1151;
	wire [12-1:0] node1154;
	wire [12-1:0] node1156;
	wire [12-1:0] node1159;
	wire [12-1:0] node1161;
	wire [12-1:0] node1162;
	wire [12-1:0] node1166;
	wire [12-1:0] node1167;
	wire [12-1:0] node1168;
	wire [12-1:0] node1169;
	wire [12-1:0] node1170;
	wire [12-1:0] node1171;
	wire [12-1:0] node1174;
	wire [12-1:0] node1176;
	wire [12-1:0] node1179;
	wire [12-1:0] node1180;
	wire [12-1:0] node1182;
	wire [12-1:0] node1185;
	wire [12-1:0] node1186;
	wire [12-1:0] node1190;
	wire [12-1:0] node1191;
	wire [12-1:0] node1192;
	wire [12-1:0] node1194;
	wire [12-1:0] node1198;
	wire [12-1:0] node1200;
	wire [12-1:0] node1202;
	wire [12-1:0] node1205;
	wire [12-1:0] node1206;
	wire [12-1:0] node1207;
	wire [12-1:0] node1208;
	wire [12-1:0] node1210;
	wire [12-1:0] node1214;
	wire [12-1:0] node1215;
	wire [12-1:0] node1219;
	wire [12-1:0] node1220;
	wire [12-1:0] node1221;
	wire [12-1:0] node1223;
	wire [12-1:0] node1226;
	wire [12-1:0] node1228;
	wire [12-1:0] node1231;
	wire [12-1:0] node1233;
	wire [12-1:0] node1236;
	wire [12-1:0] node1237;
	wire [12-1:0] node1238;
	wire [12-1:0] node1239;
	wire [12-1:0] node1241;
	wire [12-1:0] node1244;
	wire [12-1:0] node1246;
	wire [12-1:0] node1247;
	wire [12-1:0] node1251;
	wire [12-1:0] node1252;
	wire [12-1:0] node1255;
	wire [12-1:0] node1257;
	wire [12-1:0] node1260;
	wire [12-1:0] node1261;
	wire [12-1:0] node1263;
	wire [12-1:0] node1266;
	wire [12-1:0] node1267;
	wire [12-1:0] node1268;
	wire [12-1:0] node1270;
	wire [12-1:0] node1273;
	wire [12-1:0] node1274;
	wire [12-1:0] node1277;
	wire [12-1:0] node1280;
	wire [12-1:0] node1282;
	wire [12-1:0] node1285;
	wire [12-1:0] node1286;
	wire [12-1:0] node1287;
	wire [12-1:0] node1288;
	wire [12-1:0] node1289;
	wire [12-1:0] node1290;
	wire [12-1:0] node1291;
	wire [12-1:0] node1293;
	wire [12-1:0] node1294;
	wire [12-1:0] node1298;
	wire [12-1:0] node1300;
	wire [12-1:0] node1301;
	wire [12-1:0] node1305;
	wire [12-1:0] node1306;
	wire [12-1:0] node1310;
	wire [12-1:0] node1311;
	wire [12-1:0] node1313;
	wire [12-1:0] node1314;
	wire [12-1:0] node1315;
	wire [12-1:0] node1318;
	wire [12-1:0] node1322;
	wire [12-1:0] node1323;
	wire [12-1:0] node1324;
	wire [12-1:0] node1326;
	wire [12-1:0] node1330;
	wire [12-1:0] node1332;
	wire [12-1:0] node1333;
	wire [12-1:0] node1337;
	wire [12-1:0] node1338;
	wire [12-1:0] node1339;
	wire [12-1:0] node1340;
	wire [12-1:0] node1341;
	wire [12-1:0] node1343;
	wire [12-1:0] node1346;
	wire [12-1:0] node1348;
	wire [12-1:0] node1351;
	wire [12-1:0] node1352;
	wire [12-1:0] node1354;
	wire [12-1:0] node1358;
	wire [12-1:0] node1359;
	wire [12-1:0] node1360;
	wire [12-1:0] node1362;
	wire [12-1:0] node1366;
	wire [12-1:0] node1368;
	wire [12-1:0] node1371;
	wire [12-1:0] node1372;
	wire [12-1:0] node1373;
	wire [12-1:0] node1375;
	wire [12-1:0] node1376;
	wire [12-1:0] node1379;
	wire [12-1:0] node1382;
	wire [12-1:0] node1384;
	wire [12-1:0] node1387;
	wire [12-1:0] node1388;
	wire [12-1:0] node1389;
	wire [12-1:0] node1392;
	wire [12-1:0] node1394;
	wire [12-1:0] node1397;
	wire [12-1:0] node1400;
	wire [12-1:0] node1401;
	wire [12-1:0] node1402;
	wire [12-1:0] node1403;
	wire [12-1:0] node1404;
	wire [12-1:0] node1406;
	wire [12-1:0] node1408;
	wire [12-1:0] node1411;
	wire [12-1:0] node1412;
	wire [12-1:0] node1414;
	wire [12-1:0] node1418;
	wire [12-1:0] node1419;
	wire [12-1:0] node1422;
	wire [12-1:0] node1425;
	wire [12-1:0] node1426;
	wire [12-1:0] node1427;
	wire [12-1:0] node1429;
	wire [12-1:0] node1432;
	wire [12-1:0] node1435;
	wire [12-1:0] node1436;
	wire [12-1:0] node1439;
	wire [12-1:0] node1441;
	wire [12-1:0] node1442;
	wire [12-1:0] node1446;
	wire [12-1:0] node1447;
	wire [12-1:0] node1448;
	wire [12-1:0] node1449;
	wire [12-1:0] node1450;
	wire [12-1:0] node1455;
	wire [12-1:0] node1456;
	wire [12-1:0] node1457;
	wire [12-1:0] node1459;
	wire [12-1:0] node1463;
	wire [12-1:0] node1466;
	wire [12-1:0] node1467;
	wire [12-1:0] node1468;
	wire [12-1:0] node1470;
	wire [12-1:0] node1472;
	wire [12-1:0] node1475;
	wire [12-1:0] node1476;
	wire [12-1:0] node1480;
	wire [12-1:0] node1481;
	wire [12-1:0] node1484;
	wire [12-1:0] node1485;
	wire [12-1:0] node1489;
	wire [12-1:0] node1490;
	wire [12-1:0] node1491;
	wire [12-1:0] node1492;
	wire [12-1:0] node1493;
	wire [12-1:0] node1494;
	wire [12-1:0] node1496;
	wire [12-1:0] node1497;
	wire [12-1:0] node1501;
	wire [12-1:0] node1503;
	wire [12-1:0] node1506;
	wire [12-1:0] node1507;
	wire [12-1:0] node1508;
	wire [12-1:0] node1509;
	wire [12-1:0] node1513;
	wire [12-1:0] node1514;
	wire [12-1:0] node1518;
	wire [12-1:0] node1521;
	wire [12-1:0] node1522;
	wire [12-1:0] node1523;
	wire [12-1:0] node1525;
	wire [12-1:0] node1526;
	wire [12-1:0] node1530;
	wire [12-1:0] node1531;
	wire [12-1:0] node1533;
	wire [12-1:0] node1537;
	wire [12-1:0] node1538;
	wire [12-1:0] node1539;
	wire [12-1:0] node1540;
	wire [12-1:0] node1543;
	wire [12-1:0] node1546;
	wire [12-1:0] node1548;
	wire [12-1:0] node1551;
	wire [12-1:0] node1552;
	wire [12-1:0] node1554;
	wire [12-1:0] node1557;
	wire [12-1:0] node1559;
	wire [12-1:0] node1562;
	wire [12-1:0] node1563;
	wire [12-1:0] node1565;
	wire [12-1:0] node1566;
	wire [12-1:0] node1567;
	wire [12-1:0] node1570;
	wire [12-1:0] node1573;
	wire [12-1:0] node1574;
	wire [12-1:0] node1576;
	wire [12-1:0] node1580;
	wire [12-1:0] node1581;
	wire [12-1:0] node1582;
	wire [12-1:0] node1584;
	wire [12-1:0] node1586;
	wire [12-1:0] node1589;
	wire [12-1:0] node1590;
	wire [12-1:0] node1594;
	wire [12-1:0] node1595;
	wire [12-1:0] node1597;
	wire [12-1:0] node1598;
	wire [12-1:0] node1601;
	wire [12-1:0] node1604;
	wire [12-1:0] node1605;
	wire [12-1:0] node1607;
	wire [12-1:0] node1611;
	wire [12-1:0] node1612;
	wire [12-1:0] node1613;
	wire [12-1:0] node1614;
	wire [12-1:0] node1615;
	wire [12-1:0] node1616;
	wire [12-1:0] node1620;
	wire [12-1:0] node1622;
	wire [12-1:0] node1623;
	wire [12-1:0] node1627;
	wire [12-1:0] node1628;
	wire [12-1:0] node1629;
	wire [12-1:0] node1631;
	wire [12-1:0] node1635;
	wire [12-1:0] node1636;
	wire [12-1:0] node1638;
	wire [12-1:0] node1641;
	wire [12-1:0] node1642;
	wire [12-1:0] node1645;
	wire [12-1:0] node1648;
	wire [12-1:0] node1649;
	wire [12-1:0] node1651;
	wire [12-1:0] node1653;
	wire [12-1:0] node1656;
	wire [12-1:0] node1657;
	wire [12-1:0] node1658;
	wire [12-1:0] node1662;
	wire [12-1:0] node1664;
	wire [12-1:0] node1665;
	wire [12-1:0] node1669;
	wire [12-1:0] node1670;
	wire [12-1:0] node1671;
	wire [12-1:0] node1672;
	wire [12-1:0] node1673;
	wire [12-1:0] node1677;
	wire [12-1:0] node1678;
	wire [12-1:0] node1680;
	wire [12-1:0] node1684;
	wire [12-1:0] node1685;
	wire [12-1:0] node1688;
	wire [12-1:0] node1691;
	wire [12-1:0] node1692;
	wire [12-1:0] node1694;
	wire [12-1:0] node1695;
	wire [12-1:0] node1697;
	wire [12-1:0] node1701;
	wire [12-1:0] node1702;
	wire [12-1:0] node1705;
	wire [12-1:0] node1706;
	wire [12-1:0] node1710;
	wire [12-1:0] node1711;
	wire [12-1:0] node1712;
	wire [12-1:0] node1713;
	wire [12-1:0] node1714;
	wire [12-1:0] node1715;
	wire [12-1:0] node1716;
	wire [12-1:0] node1717;
	wire [12-1:0] node1718;
	wire [12-1:0] node1719;
	wire [12-1:0] node1721;
	wire [12-1:0] node1724;
	wire [12-1:0] node1725;
	wire [12-1:0] node1729;
	wire [12-1:0] node1732;
	wire [12-1:0] node1733;
	wire [12-1:0] node1735;
	wire [12-1:0] node1736;
	wire [12-1:0] node1740;
	wire [12-1:0] node1743;
	wire [12-1:0] node1744;
	wire [12-1:0] node1745;
	wire [12-1:0] node1746;
	wire [12-1:0] node1747;
	wire [12-1:0] node1750;
	wire [12-1:0] node1754;
	wire [12-1:0] node1756;
	wire [12-1:0] node1759;
	wire [12-1:0] node1760;
	wire [12-1:0] node1761;
	wire [12-1:0] node1764;
	wire [12-1:0] node1765;
	wire [12-1:0] node1769;
	wire [12-1:0] node1770;
	wire [12-1:0] node1771;
	wire [12-1:0] node1776;
	wire [12-1:0] node1777;
	wire [12-1:0] node1778;
	wire [12-1:0] node1779;
	wire [12-1:0] node1781;
	wire [12-1:0] node1784;
	wire [12-1:0] node1787;
	wire [12-1:0] node1788;
	wire [12-1:0] node1790;
	wire [12-1:0] node1791;
	wire [12-1:0] node1795;
	wire [12-1:0] node1797;
	wire [12-1:0] node1800;
	wire [12-1:0] node1801;
	wire [12-1:0] node1802;
	wire [12-1:0] node1803;
	wire [12-1:0] node1805;
	wire [12-1:0] node1808;
	wire [12-1:0] node1809;
	wire [12-1:0] node1813;
	wire [12-1:0] node1815;
	wire [12-1:0] node1816;
	wire [12-1:0] node1821;
	wire [12-1:0] node1822;
	wire [12-1:0] node1823;
	wire [12-1:0] node1824;
	wire [12-1:0] node1825;
	wire [12-1:0] node1826;
	wire [12-1:0] node1827;
	wire [12-1:0] node1831;
	wire [12-1:0] node1832;
	wire [12-1:0] node1836;
	wire [12-1:0] node1837;
	wire [12-1:0] node1839;
	wire [12-1:0] node1842;
	wire [12-1:0] node1843;
	wire [12-1:0] node1847;
	wire [12-1:0] node1848;
	wire [12-1:0] node1849;
	wire [12-1:0] node1853;
	wire [12-1:0] node1854;
	wire [12-1:0] node1855;
	wire [12-1:0] node1859;
	wire [12-1:0] node1860;
	wire [12-1:0] node1864;
	wire [12-1:0] node1865;
	wire [12-1:0] node1866;
	wire [12-1:0] node1867;
	wire [12-1:0] node1868;
	wire [12-1:0] node1873;
	wire [12-1:0] node1875;
	wire [12-1:0] node1878;
	wire [12-1:0] node1879;
	wire [12-1:0] node1880;
	wire [12-1:0] node1884;
	wire [12-1:0] node1885;
	wire [12-1:0] node1887;
	wire [12-1:0] node1891;
	wire [12-1:0] node1892;
	wire [12-1:0] node1893;
	wire [12-1:0] node1894;
	wire [12-1:0] node1896;
	wire [12-1:0] node1899;
	wire [12-1:0] node1900;
	wire [12-1:0] node1904;
	wire [12-1:0] node1905;
	wire [12-1:0] node1906;
	wire [12-1:0] node1908;
	wire [12-1:0] node1912;
	wire [12-1:0] node1914;
	wire [12-1:0] node1917;
	wire [12-1:0] node1918;
	wire [12-1:0] node1919;
	wire [12-1:0] node1920;
	wire [12-1:0] node1921;
	wire [12-1:0] node1926;
	wire [12-1:0] node1929;
	wire [12-1:0] node1930;
	wire [12-1:0] node1931;
	wire [12-1:0] node1933;
	wire [12-1:0] node1937;
	wire [12-1:0] node1938;
	wire [12-1:0] node1940;
	wire [12-1:0] node1943;
	wire [12-1:0] node1946;
	wire [12-1:0] node1947;
	wire [12-1:0] node1948;
	wire [12-1:0] node1949;
	wire [12-1:0] node1950;
	wire [12-1:0] node1951;
	wire [12-1:0] node1953;
	wire [12-1:0] node1954;
	wire [12-1:0] node1958;
	wire [12-1:0] node1961;
	wire [12-1:0] node1962;
	wire [12-1:0] node1964;
	wire [12-1:0] node1965;
	wire [12-1:0] node1969;
	wire [12-1:0] node1971;
	wire [12-1:0] node1972;
	wire [12-1:0] node1976;
	wire [12-1:0] node1977;
	wire [12-1:0] node1978;
	wire [12-1:0] node1980;
	wire [12-1:0] node1983;
	wire [12-1:0] node1985;
	wire [12-1:0] node1988;
	wire [12-1:0] node1989;
	wire [12-1:0] node1992;
	wire [12-1:0] node1993;
	wire [12-1:0] node1995;
	wire [12-1:0] node1999;
	wire [12-1:0] node2000;
	wire [12-1:0] node2001;
	wire [12-1:0] node2002;
	wire [12-1:0] node2004;
	wire [12-1:0] node2005;
	wire [12-1:0] node2010;
	wire [12-1:0] node2011;
	wire [12-1:0] node2012;
	wire [12-1:0] node2014;
	wire [12-1:0] node2017;
	wire [12-1:0] node2018;
	wire [12-1:0] node2022;
	wire [12-1:0] node2025;
	wire [12-1:0] node2026;
	wire [12-1:0] node2027;
	wire [12-1:0] node2028;
	wire [12-1:0] node2032;
	wire [12-1:0] node2033;
	wire [12-1:0] node2035;
	wire [12-1:0] node2039;
	wire [12-1:0] node2040;
	wire [12-1:0] node2042;
	wire [12-1:0] node2043;
	wire [12-1:0] node2046;
	wire [12-1:0] node2049;
	wire [12-1:0] node2050;
	wire [12-1:0] node2054;
	wire [12-1:0] node2055;
	wire [12-1:0] node2056;
	wire [12-1:0] node2057;
	wire [12-1:0] node2058;
	wire [12-1:0] node2059;
	wire [12-1:0] node2061;
	wire [12-1:0] node2064;
	wire [12-1:0] node2065;
	wire [12-1:0] node2069;
	wire [12-1:0] node2072;
	wire [12-1:0] node2073;
	wire [12-1:0] node2076;
	wire [12-1:0] node2077;
	wire [12-1:0] node2079;
	wire [12-1:0] node2083;
	wire [12-1:0] node2084;
	wire [12-1:0] node2085;
	wire [12-1:0] node2086;
	wire [12-1:0] node2088;
	wire [12-1:0] node2092;
	wire [12-1:0] node2094;
	wire [12-1:0] node2095;
	wire [12-1:0] node2099;
	wire [12-1:0] node2100;
	wire [12-1:0] node2101;
	wire [12-1:0] node2102;
	wire [12-1:0] node2106;
	wire [12-1:0] node2108;
	wire [12-1:0] node2111;
	wire [12-1:0] node2112;
	wire [12-1:0] node2114;
	wire [12-1:0] node2117;
	wire [12-1:0] node2120;
	wire [12-1:0] node2121;
	wire [12-1:0] node2122;
	wire [12-1:0] node2123;
	wire [12-1:0] node2124;
	wire [12-1:0] node2126;
	wire [12-1:0] node2130;
	wire [12-1:0] node2133;
	wire [12-1:0] node2134;
	wire [12-1:0] node2135;
	wire [12-1:0] node2137;
	wire [12-1:0] node2140;
	wire [12-1:0] node2141;
	wire [12-1:0] node2144;
	wire [12-1:0] node2148;
	wire [12-1:0] node2149;
	wire [12-1:0] node2150;
	wire [12-1:0] node2152;
	wire [12-1:0] node2154;
	wire [12-1:0] node2157;
	wire [12-1:0] node2158;
	wire [12-1:0] node2160;
	wire [12-1:0] node2164;
	wire [12-1:0] node2165;
	wire [12-1:0] node2167;
	wire [12-1:0] node2169;
	wire [12-1:0] node2172;
	wire [12-1:0] node2173;
	wire [12-1:0] node2176;
	wire [12-1:0] node2178;
	wire [12-1:0] node2181;
	wire [12-1:0] node2182;
	wire [12-1:0] node2183;
	wire [12-1:0] node2184;
	wire [12-1:0] node2185;
	wire [12-1:0] node2186;
	wire [12-1:0] node2188;
	wire [12-1:0] node2189;
	wire [12-1:0] node2190;
	wire [12-1:0] node2195;
	wire [12-1:0] node2196;
	wire [12-1:0] node2199;
	wire [12-1:0] node2201;
	wire [12-1:0] node2204;
	wire [12-1:0] node2205;
	wire [12-1:0] node2206;
	wire [12-1:0] node2207;
	wire [12-1:0] node2211;
	wire [12-1:0] node2212;
	wire [12-1:0] node2214;
	wire [12-1:0] node2218;
	wire [12-1:0] node2219;
	wire [12-1:0] node2220;
	wire [12-1:0] node2222;
	wire [12-1:0] node2227;
	wire [12-1:0] node2228;
	wire [12-1:0] node2229;
	wire [12-1:0] node2230;
	wire [12-1:0] node2231;
	wire [12-1:0] node2232;
	wire [12-1:0] node2236;
	wire [12-1:0] node2237;
	wire [12-1:0] node2241;
	wire [12-1:0] node2244;
	wire [12-1:0] node2245;
	wire [12-1:0] node2246;
	wire [12-1:0] node2248;
	wire [12-1:0] node2252;
	wire [12-1:0] node2255;
	wire [12-1:0] node2256;
	wire [12-1:0] node2257;
	wire [12-1:0] node2258;
	wire [12-1:0] node2262;
	wire [12-1:0] node2264;
	wire [12-1:0] node2267;
	wire [12-1:0] node2268;
	wire [12-1:0] node2269;
	wire [12-1:0] node2272;
	wire [12-1:0] node2273;
	wire [12-1:0] node2277;
	wire [12-1:0] node2279;
	wire [12-1:0] node2280;
	wire [12-1:0] node2284;
	wire [12-1:0] node2285;
	wire [12-1:0] node2286;
	wire [12-1:0] node2287;
	wire [12-1:0] node2288;
	wire [12-1:0] node2290;
	wire [12-1:0] node2291;
	wire [12-1:0] node2295;
	wire [12-1:0] node2297;
	wire [12-1:0] node2300;
	wire [12-1:0] node2303;
	wire [12-1:0] node2304;
	wire [12-1:0] node2306;
	wire [12-1:0] node2308;
	wire [12-1:0] node2311;
	wire [12-1:0] node2312;
	wire [12-1:0] node2313;
	wire [12-1:0] node2314;
	wire [12-1:0] node2319;
	wire [12-1:0] node2320;
	wire [12-1:0] node2323;
	wire [12-1:0] node2325;
	wire [12-1:0] node2328;
	wire [12-1:0] node2329;
	wire [12-1:0] node2330;
	wire [12-1:0] node2332;
	wire [12-1:0] node2333;
	wire [12-1:0] node2335;
	wire [12-1:0] node2339;
	wire [12-1:0] node2340;
	wire [12-1:0] node2341;
	wire [12-1:0] node2345;
	wire [12-1:0] node2347;
	wire [12-1:0] node2350;
	wire [12-1:0] node2351;
	wire [12-1:0] node2352;
	wire [12-1:0] node2353;
	wire [12-1:0] node2357;
	wire [12-1:0] node2359;
	wire [12-1:0] node2362;
	wire [12-1:0] node2363;
	wire [12-1:0] node2366;
	wire [12-1:0] node2367;
	wire [12-1:0] node2371;
	wire [12-1:0] node2372;
	wire [12-1:0] node2373;
	wire [12-1:0] node2374;
	wire [12-1:0] node2375;
	wire [12-1:0] node2377;
	wire [12-1:0] node2378;
	wire [12-1:0] node2379;
	wire [12-1:0] node2382;
	wire [12-1:0] node2385;
	wire [12-1:0] node2386;
	wire [12-1:0] node2390;
	wire [12-1:0] node2391;
	wire [12-1:0] node2392;
	wire [12-1:0] node2396;
	wire [12-1:0] node2398;
	wire [12-1:0] node2399;
	wire [12-1:0] node2403;
	wire [12-1:0] node2404;
	wire [12-1:0] node2405;
	wire [12-1:0] node2406;
	wire [12-1:0] node2408;
	wire [12-1:0] node2411;
	wire [12-1:0] node2413;
	wire [12-1:0] node2416;
	wire [12-1:0] node2417;
	wire [12-1:0] node2419;
	wire [12-1:0] node2422;
	wire [12-1:0] node2423;
	wire [12-1:0] node2427;
	wire [12-1:0] node2428;
	wire [12-1:0] node2429;
	wire [12-1:0] node2431;
	wire [12-1:0] node2434;
	wire [12-1:0] node2436;
	wire [12-1:0] node2439;
	wire [12-1:0] node2440;
	wire [12-1:0] node2444;
	wire [12-1:0] node2445;
	wire [12-1:0] node2446;
	wire [12-1:0] node2447;
	wire [12-1:0] node2448;
	wire [12-1:0] node2453;
	wire [12-1:0] node2454;
	wire [12-1:0] node2455;
	wire [12-1:0] node2459;
	wire [12-1:0] node2460;
	wire [12-1:0] node2463;
	wire [12-1:0] node2465;
	wire [12-1:0] node2468;
	wire [12-1:0] node2469;
	wire [12-1:0] node2470;
	wire [12-1:0] node2473;
	wire [12-1:0] node2474;
	wire [12-1:0] node2476;
	wire [12-1:0] node2479;
	wire [12-1:0] node2480;
	wire [12-1:0] node2484;
	wire [12-1:0] node2485;
	wire [12-1:0] node2488;
	wire [12-1:0] node2491;
	wire [12-1:0] node2492;
	wire [12-1:0] node2493;
	wire [12-1:0] node2494;
	wire [12-1:0] node2496;
	wire [12-1:0] node2497;
	wire [12-1:0] node2499;
	wire [12-1:0] node2503;
	wire [12-1:0] node2504;
	wire [12-1:0] node2505;
	wire [12-1:0] node2507;
	wire [12-1:0] node2510;
	wire [12-1:0] node2513;
	wire [12-1:0] node2515;
	wire [12-1:0] node2518;
	wire [12-1:0] node2519;
	wire [12-1:0] node2520;
	wire [12-1:0] node2521;
	wire [12-1:0] node2525;
	wire [12-1:0] node2526;
	wire [12-1:0] node2527;
	wire [12-1:0] node2530;
	wire [12-1:0] node2534;
	wire [12-1:0] node2535;
	wire [12-1:0] node2537;
	wire [12-1:0] node2538;
	wire [12-1:0] node2542;
	wire [12-1:0] node2545;
	wire [12-1:0] node2546;
	wire [12-1:0] node2547;
	wire [12-1:0] node2548;
	wire [12-1:0] node2550;
	wire [12-1:0] node2551;
	wire [12-1:0] node2555;
	wire [12-1:0] node2557;
	wire [12-1:0] node2560;
	wire [12-1:0] node2561;
	wire [12-1:0] node2562;
	wire [12-1:0] node2565;
	wire [12-1:0] node2568;
	wire [12-1:0] node2569;
	wire [12-1:0] node2571;
	wire [12-1:0] node2574;
	wire [12-1:0] node2577;
	wire [12-1:0] node2578;
	wire [12-1:0] node2579;
	wire [12-1:0] node2582;
	wire [12-1:0] node2583;
	wire [12-1:0] node2584;
	wire [12-1:0] node2588;
	wire [12-1:0] node2589;
	wire [12-1:0] node2593;
	wire [12-1:0] node2594;
	wire [12-1:0] node2595;
	wire [12-1:0] node2599;
	wire [12-1:0] node2602;
	wire [12-1:0] node2603;
	wire [12-1:0] node2604;
	wire [12-1:0] node2605;
	wire [12-1:0] node2606;
	wire [12-1:0] node2607;
	wire [12-1:0] node2608;
	wire [12-1:0] node2609;
	wire [12-1:0] node2610;
	wire [12-1:0] node2611;
	wire [12-1:0] node2616;
	wire [12-1:0] node2617;
	wire [12-1:0] node2620;
	wire [12-1:0] node2621;
	wire [12-1:0] node2625;
	wire [12-1:0] node2626;
	wire [12-1:0] node2628;
	wire [12-1:0] node2632;
	wire [12-1:0] node2633;
	wire [12-1:0] node2634;
	wire [12-1:0] node2636;
	wire [12-1:0] node2637;
	wire [12-1:0] node2640;
	wire [12-1:0] node2643;
	wire [12-1:0] node2646;
	wire [12-1:0] node2647;
	wire [12-1:0] node2650;
	wire [12-1:0] node2652;
	wire [12-1:0] node2655;
	wire [12-1:0] node2656;
	wire [12-1:0] node2657;
	wire [12-1:0] node2658;
	wire [12-1:0] node2659;
	wire [12-1:0] node2661;
	wire [12-1:0] node2665;
	wire [12-1:0] node2666;
	wire [12-1:0] node2668;
	wire [12-1:0] node2672;
	wire [12-1:0] node2673;
	wire [12-1:0] node2676;
	wire [12-1:0] node2678;
	wire [12-1:0] node2681;
	wire [12-1:0] node2682;
	wire [12-1:0] node2683;
	wire [12-1:0] node2686;
	wire [12-1:0] node2688;
	wire [12-1:0] node2691;
	wire [12-1:0] node2692;
	wire [12-1:0] node2693;
	wire [12-1:0] node2695;
	wire [12-1:0] node2699;
	wire [12-1:0] node2702;
	wire [12-1:0] node2703;
	wire [12-1:0] node2704;
	wire [12-1:0] node2705;
	wire [12-1:0] node2706;
	wire [12-1:0] node2707;
	wire [12-1:0] node2709;
	wire [12-1:0] node2713;
	wire [12-1:0] node2716;
	wire [12-1:0] node2717;
	wire [12-1:0] node2718;
	wire [12-1:0] node2722;
	wire [12-1:0] node2724;
	wire [12-1:0] node2725;
	wire [12-1:0] node2729;
	wire [12-1:0] node2730;
	wire [12-1:0] node2732;
	wire [12-1:0] node2735;
	wire [12-1:0] node2736;
	wire [12-1:0] node2740;
	wire [12-1:0] node2741;
	wire [12-1:0] node2742;
	wire [12-1:0] node2743;
	wire [12-1:0] node2744;
	wire [12-1:0] node2746;
	wire [12-1:0] node2750;
	wire [12-1:0] node2753;
	wire [12-1:0] node2754;
	wire [12-1:0] node2757;
	wire [12-1:0] node2760;
	wire [12-1:0] node2761;
	wire [12-1:0] node2762;
	wire [12-1:0] node2763;
	wire [12-1:0] node2765;
	wire [12-1:0] node2769;
	wire [12-1:0] node2771;
	wire [12-1:0] node2774;
	wire [12-1:0] node2775;
	wire [12-1:0] node2776;
	wire [12-1:0] node2780;
	wire [12-1:0] node2782;
	wire [12-1:0] node2785;
	wire [12-1:0] node2786;
	wire [12-1:0] node2787;
	wire [12-1:0] node2788;
	wire [12-1:0] node2789;
	wire [12-1:0] node2790;
	wire [12-1:0] node2791;
	wire [12-1:0] node2792;
	wire [12-1:0] node2797;
	wire [12-1:0] node2798;
	wire [12-1:0] node2799;
	wire [12-1:0] node2802;
	wire [12-1:0] node2805;
	wire [12-1:0] node2807;
	wire [12-1:0] node2810;
	wire [12-1:0] node2811;
	wire [12-1:0] node2812;
	wire [12-1:0] node2814;
	wire [12-1:0] node2818;
	wire [12-1:0] node2820;
	wire [12-1:0] node2823;
	wire [12-1:0] node2824;
	wire [12-1:0] node2825;
	wire [12-1:0] node2828;
	wire [12-1:0] node2829;
	wire [12-1:0] node2833;
	wire [12-1:0] node2834;
	wire [12-1:0] node2837;
	wire [12-1:0] node2840;
	wire [12-1:0] node2841;
	wire [12-1:0] node2842;
	wire [12-1:0] node2843;
	wire [12-1:0] node2844;
	wire [12-1:0] node2848;
	wire [12-1:0] node2850;
	wire [12-1:0] node2853;
	wire [12-1:0] node2854;
	wire [12-1:0] node2855;
	wire [12-1:0] node2857;
	wire [12-1:0] node2861;
	wire [12-1:0] node2862;
	wire [12-1:0] node2863;
	wire [12-1:0] node2867;
	wire [12-1:0] node2868;
	wire [12-1:0] node2872;
	wire [12-1:0] node2873;
	wire [12-1:0] node2874;
	wire [12-1:0] node2875;
	wire [12-1:0] node2876;
	wire [12-1:0] node2881;
	wire [12-1:0] node2882;
	wire [12-1:0] node2883;
	wire [12-1:0] node2886;
	wire [12-1:0] node2889;
	wire [12-1:0] node2890;
	wire [12-1:0] node2894;
	wire [12-1:0] node2895;
	wire [12-1:0] node2896;
	wire [12-1:0] node2898;
	wire [12-1:0] node2901;
	wire [12-1:0] node2902;
	wire [12-1:0] node2906;
	wire [12-1:0] node2909;
	wire [12-1:0] node2910;
	wire [12-1:0] node2911;
	wire [12-1:0] node2912;
	wire [12-1:0] node2913;
	wire [12-1:0] node2915;
	wire [12-1:0] node2918;
	wire [12-1:0] node2921;
	wire [12-1:0] node2922;
	wire [12-1:0] node2926;
	wire [12-1:0] node2927;
	wire [12-1:0] node2929;
	wire [12-1:0] node2930;
	wire [12-1:0] node2931;
	wire [12-1:0] node2935;
	wire [12-1:0] node2936;
	wire [12-1:0] node2940;
	wire [12-1:0] node2941;
	wire [12-1:0] node2944;
	wire [12-1:0] node2946;
	wire [12-1:0] node2947;
	wire [12-1:0] node2951;
	wire [12-1:0] node2952;
	wire [12-1:0] node2953;
	wire [12-1:0] node2954;
	wire [12-1:0] node2956;
	wire [12-1:0] node2958;
	wire [12-1:0] node2961;
	wire [12-1:0] node2962;
	wire [12-1:0] node2964;
	wire [12-1:0] node2968;
	wire [12-1:0] node2969;
	wire [12-1:0] node2972;
	wire [12-1:0] node2975;
	wire [12-1:0] node2976;
	wire [12-1:0] node2977;
	wire [12-1:0] node2979;
	wire [12-1:0] node2980;
	wire [12-1:0] node2984;
	wire [12-1:0] node2987;
	wire [12-1:0] node2988;
	wire [12-1:0] node2989;
	wire [12-1:0] node2991;
	wire [12-1:0] node2995;
	wire [12-1:0] node2997;
	wire [12-1:0] node2998;
	wire [12-1:0] node3002;
	wire [12-1:0] node3003;
	wire [12-1:0] node3004;
	wire [12-1:0] node3005;
	wire [12-1:0] node3006;
	wire [12-1:0] node3007;
	wire [12-1:0] node3010;
	wire [12-1:0] node3011;
	wire [12-1:0] node3013;
	wire [12-1:0] node3016;
	wire [12-1:0] node3019;
	wire [12-1:0] node3020;
	wire [12-1:0] node3021;
	wire [12-1:0] node3023;
	wire [12-1:0] node3024;
	wire [12-1:0] node3027;
	wire [12-1:0] node3030;
	wire [12-1:0] node3032;
	wire [12-1:0] node3033;
	wire [12-1:0] node3037;
	wire [12-1:0] node3038;
	wire [12-1:0] node3039;
	wire [12-1:0] node3041;
	wire [12-1:0] node3045;
	wire [12-1:0] node3048;
	wire [12-1:0] node3049;
	wire [12-1:0] node3050;
	wire [12-1:0] node3051;
	wire [12-1:0] node3052;
	wire [12-1:0] node3054;
	wire [12-1:0] node3058;
	wire [12-1:0] node3060;
	wire [12-1:0] node3061;
	wire [12-1:0] node3065;
	wire [12-1:0] node3066;
	wire [12-1:0] node3068;
	wire [12-1:0] node3069;
	wire [12-1:0] node3072;
	wire [12-1:0] node3076;
	wire [12-1:0] node3077;
	wire [12-1:0] node3078;
	wire [12-1:0] node3079;
	wire [12-1:0] node3081;
	wire [12-1:0] node3085;
	wire [12-1:0] node3086;
	wire [12-1:0] node3087;
	wire [12-1:0] node3090;
	wire [12-1:0] node3094;
	wire [12-1:0] node3095;
	wire [12-1:0] node3096;
	wire [12-1:0] node3100;
	wire [12-1:0] node3101;
	wire [12-1:0] node3103;
	wire [12-1:0] node3107;
	wire [12-1:0] node3108;
	wire [12-1:0] node3109;
	wire [12-1:0] node3110;
	wire [12-1:0] node3111;
	wire [12-1:0] node3113;
	wire [12-1:0] node3114;
	wire [12-1:0] node3118;
	wire [12-1:0] node3119;
	wire [12-1:0] node3121;
	wire [12-1:0] node3125;
	wire [12-1:0] node3126;
	wire [12-1:0] node3127;
	wire [12-1:0] node3131;
	wire [12-1:0] node3132;
	wire [12-1:0] node3136;
	wire [12-1:0] node3137;
	wire [12-1:0] node3139;
	wire [12-1:0] node3140;
	wire [12-1:0] node3144;
	wire [12-1:0] node3146;
	wire [12-1:0] node3148;
	wire [12-1:0] node3151;
	wire [12-1:0] node3152;
	wire [12-1:0] node3153;
	wire [12-1:0] node3155;
	wire [12-1:0] node3158;
	wire [12-1:0] node3159;
	wire [12-1:0] node3160;
	wire [12-1:0] node3162;
	wire [12-1:0] node3165;
	wire [12-1:0] node3166;
	wire [12-1:0] node3170;
	wire [12-1:0] node3171;
	wire [12-1:0] node3173;
	wire [12-1:0] node3176;
	wire [12-1:0] node3177;
	wire [12-1:0] node3181;
	wire [12-1:0] node3182;
	wire [12-1:0] node3184;
	wire [12-1:0] node3187;
	wire [12-1:0] node3188;
	wire [12-1:0] node3191;
	wire [12-1:0] node3193;
	wire [12-1:0] node3194;
	wire [12-1:0] node3198;
	wire [12-1:0] node3199;
	wire [12-1:0] node3200;
	wire [12-1:0] node3201;
	wire [12-1:0] node3202;
	wire [12-1:0] node3204;
	wire [12-1:0] node3205;
	wire [12-1:0] node3206;
	wire [12-1:0] node3210;
	wire [12-1:0] node3211;
	wire [12-1:0] node3215;
	wire [12-1:0] node3216;
	wire [12-1:0] node3217;
	wire [12-1:0] node3218;
	wire [12-1:0] node3222;
	wire [12-1:0] node3224;
	wire [12-1:0] node3227;
	wire [12-1:0] node3229;
	wire [12-1:0] node3232;
	wire [12-1:0] node3233;
	wire [12-1:0] node3234;
	wire [12-1:0] node3236;
	wire [12-1:0] node3237;
	wire [12-1:0] node3241;
	wire [12-1:0] node3242;
	wire [12-1:0] node3243;
	wire [12-1:0] node3248;
	wire [12-1:0] node3249;
	wire [12-1:0] node3251;
	wire [12-1:0] node3252;
	wire [12-1:0] node3255;
	wire [12-1:0] node3258;
	wire [12-1:0] node3261;
	wire [12-1:0] node3262;
	wire [12-1:0] node3263;
	wire [12-1:0] node3264;
	wire [12-1:0] node3266;
	wire [12-1:0] node3268;
	wire [12-1:0] node3271;
	wire [12-1:0] node3272;
	wire [12-1:0] node3276;
	wire [12-1:0] node3277;
	wire [12-1:0] node3280;
	wire [12-1:0] node3283;
	wire [12-1:0] node3284;
	wire [12-1:0] node3285;
	wire [12-1:0] node3286;
	wire [12-1:0] node3290;
	wire [12-1:0] node3291;
	wire [12-1:0] node3293;
	wire [12-1:0] node3297;
	wire [12-1:0] node3298;
	wire [12-1:0] node3299;
	wire [12-1:0] node3301;
	wire [12-1:0] node3304;
	wire [12-1:0] node3305;
	wire [12-1:0] node3308;
	wire [12-1:0] node3311;
	wire [12-1:0] node3313;
	wire [12-1:0] node3316;
	wire [12-1:0] node3317;
	wire [12-1:0] node3318;
	wire [12-1:0] node3319;
	wire [12-1:0] node3320;
	wire [12-1:0] node3323;
	wire [12-1:0] node3324;
	wire [12-1:0] node3326;
	wire [12-1:0] node3330;
	wire [12-1:0] node3331;
	wire [12-1:0] node3332;
	wire [12-1:0] node3336;
	wire [12-1:0] node3338;
	wire [12-1:0] node3339;
	wire [12-1:0] node3343;
	wire [12-1:0] node3344;
	wire [12-1:0] node3345;
	wire [12-1:0] node3346;
	wire [12-1:0] node3348;
	wire [12-1:0] node3352;
	wire [12-1:0] node3353;
	wire [12-1:0] node3357;
	wire [12-1:0] node3358;
	wire [12-1:0] node3360;
	wire [12-1:0] node3361;
	wire [12-1:0] node3365;
	wire [12-1:0] node3367;
	wire [12-1:0] node3370;
	wire [12-1:0] node3371;
	wire [12-1:0] node3372;
	wire [12-1:0] node3373;
	wire [12-1:0] node3374;
	wire [12-1:0] node3378;
	wire [12-1:0] node3379;
	wire [12-1:0] node3381;
	wire [12-1:0] node3384;
	wire [12-1:0] node3387;
	wire [12-1:0] node3388;
	wire [12-1:0] node3389;
	wire [12-1:0] node3391;
	wire [12-1:0] node3395;
	wire [12-1:0] node3396;
	wire [12-1:0] node3398;
	wire [12-1:0] node3401;
	wire [12-1:0] node3402;
	wire [12-1:0] node3406;
	wire [12-1:0] node3407;
	wire [12-1:0] node3408;
	wire [12-1:0] node3410;
	wire [12-1:0] node3411;
	wire [12-1:0] node3415;
	wire [12-1:0] node3417;
	wire [12-1:0] node3419;
	wire [12-1:0] node3422;
	wire [12-1:0] node3424;
	wire [12-1:0] node3425;
	wire [12-1:0] node3427;

	assign outp = (inp[3]) ? node1710 : node1;
		assign node1 = (inp[2]) ? node835 : node2;
			assign node2 = (inp[7]) ? node410 : node3;
				assign node3 = (inp[8]) ? node205 : node4;
					assign node4 = (inp[9]) ? node106 : node5;
						assign node5 = (inp[0]) ? node59 : node6;
							assign node6 = (inp[4]) ? node34 : node7;
								assign node7 = (inp[5]) ? node19 : node8;
									assign node8 = (inp[6]) ? node16 : node9;
										assign node9 = (inp[11]) ? node11 : 12'b011111111111;
											assign node11 = (inp[10]) ? 12'b001111111111 : node12;
												assign node12 = (inp[1]) ? 12'b001111111111 : 12'b011111111111;
										assign node16 = (inp[11]) ? 12'b000111111111 : 12'b001111111111;
									assign node19 = (inp[11]) ? node27 : node20;
										assign node20 = (inp[10]) ? 12'b000111111111 : node21;
											assign node21 = (inp[1]) ? 12'b001111111111 : node22;
												assign node22 = (inp[6]) ? 12'b001111111111 : 12'b011111111111;
										assign node27 = (inp[6]) ? 12'b000011111111 : node28;
											assign node28 = (inp[10]) ? node30 : 12'b000111111111;
												assign node30 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
								assign node34 = (inp[11]) ? node50 : node35;
									assign node35 = (inp[5]) ? node39 : node36;
										assign node36 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
										assign node39 = (inp[6]) ? node45 : node40;
											assign node40 = (inp[10]) ? 12'b000111111111 : node41;
												assign node41 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
											assign node45 = (inp[10]) ? 12'b000011111111 : node46;
												assign node46 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
									assign node50 = (inp[1]) ? 12'b000011111111 : node51;
										assign node51 = (inp[10]) ? node53 : 12'b000111111111;
											assign node53 = (inp[5]) ? 12'b000011111111 : node54;
												assign node54 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
							assign node59 = (inp[5]) ? node83 : node60;
								assign node60 = (inp[1]) ? node72 : node61;
									assign node61 = (inp[4]) ? node67 : node62;
										assign node62 = (inp[6]) ? 12'b000111111111 : node63;
											assign node63 = (inp[10]) ? 12'b001111111111 : 12'b011111111111;
										assign node67 = (inp[6]) ? node69 : 12'b000111111111;
											assign node69 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
									assign node72 = (inp[11]) ? node80 : node73;
										assign node73 = (inp[10]) ? node75 : 12'b000111111111;
											assign node75 = (inp[4]) ? 12'b000011111111 : node76;
												assign node76 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
										assign node80 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
								assign node83 = (inp[4]) ? node95 : node84;
									assign node84 = (inp[11]) ? node90 : node85;
										assign node85 = (inp[10]) ? node87 : 12'b000111111111;
											assign node87 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
										assign node90 = (inp[6]) ? 12'b000001111111 : node91;
											assign node91 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
									assign node95 = (inp[10]) ? node97 : 12'b000011111111;
										assign node97 = (inp[1]) ? node103 : node98;
											assign node98 = (inp[11]) ? 12'b000001111111 : node99;
												assign node99 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
											assign node103 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
						assign node106 = (inp[11]) ? node170 : node107;
							assign node107 = (inp[4]) ? node147 : node108;
								assign node108 = (inp[0]) ? node128 : node109;
									assign node109 = (inp[10]) ? node119 : node110;
										assign node110 = (inp[5]) ? node116 : node111;
											assign node111 = (inp[1]) ? 12'b001111111111 : node112;
												assign node112 = (inp[6]) ? 12'b001111111111 : 12'b011111111111;
											assign node116 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
										assign node119 = (inp[1]) ? node123 : node120;
											assign node120 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
											assign node123 = (inp[6]) ? 12'b000011111111 : node124;
												assign node124 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node128 = (inp[5]) ? node140 : node129;
										assign node129 = (inp[6]) ? node135 : node130;
											assign node130 = (inp[1]) ? 12'b000111111111 : node131;
												assign node131 = (inp[10]) ? 12'b000111111111 : 12'b001111111111;
											assign node135 = (inp[1]) ? 12'b000011111111 : node136;
												assign node136 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
										assign node140 = (inp[6]) ? 12'b000001111111 : node141;
											assign node141 = (inp[1]) ? node143 : 12'b000011111111;
												assign node143 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
								assign node147 = (inp[10]) ? node157 : node148;
									assign node148 = (inp[1]) ? node154 : node149;
										assign node149 = (inp[0]) ? 12'b000011111111 : node150;
											assign node150 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
										assign node154 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node157 = (inp[1]) ? node161 : node158;
										assign node158 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
										assign node161 = (inp[5]) ? node165 : node162;
											assign node162 = (inp[0]) ? 12'b000000111111 : 12'b000011111111;
											assign node165 = (inp[6]) ? node167 : 12'b000000111111;
												assign node167 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
							assign node170 = (inp[5]) ? node188 : node171;
								assign node171 = (inp[0]) ? node181 : node172;
									assign node172 = (inp[6]) ? node176 : node173;
										assign node173 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
										assign node176 = (inp[10]) ? node178 : 12'b000011111111;
											assign node178 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node181 = (inp[4]) ? node185 : node182;
										assign node182 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
										assign node185 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
								assign node188 = (inp[1]) ? node194 : node189;
									assign node189 = (inp[10]) ? 12'b000001111111 : node190;
										assign node190 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node194 = (inp[6]) ? node202 : node195;
										assign node195 = (inp[4]) ? node197 : 12'b000001111111;
											assign node197 = (inp[10]) ? 12'b000000111111 : node198;
												assign node198 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node202 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
					assign node205 = (inp[5]) ? node309 : node206;
						assign node206 = (inp[9]) ? node262 : node207;
							assign node207 = (inp[0]) ? node227 : node208;
								assign node208 = (inp[1]) ? node218 : node209;
									assign node209 = (inp[4]) ? node215 : node210;
										assign node210 = (inp[11]) ? node212 : 12'b001111111111;
											assign node212 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
										assign node215 = (inp[11]) ? 12'b000011111111 : 12'b000111111111;
									assign node218 = (inp[10]) ? 12'b000011111111 : node219;
										assign node219 = (inp[4]) ? node221 : 12'b000111111111;
											assign node221 = (inp[11]) ? 12'b000011111111 : node222;
												assign node222 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
								assign node227 = (inp[11]) ? node247 : node228;
									assign node228 = (inp[1]) ? node240 : node229;
										assign node229 = (inp[10]) ? node235 : node230;
											assign node230 = (inp[4]) ? node232 : 12'b000111111111;
												assign node232 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
											assign node235 = (inp[4]) ? 12'b000011111111 : node236;
												assign node236 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
										assign node240 = (inp[4]) ? 12'b000001111111 : node241;
											assign node241 = (inp[6]) ? node243 : 12'b000011111111;
												assign node243 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
									assign node247 = (inp[4]) ? node253 : node248;
										assign node248 = (inp[10]) ? node250 : 12'b000011111111;
											assign node250 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
										assign node253 = (inp[6]) ? node259 : node254;
											assign node254 = (inp[10]) ? 12'b000001111111 : node255;
												assign node255 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
											assign node259 = (inp[1]) ? 12'b000000011111 : 12'b000001111111;
							assign node262 = (inp[1]) ? node290 : node263;
								assign node263 = (inp[11]) ? node279 : node264;
									assign node264 = (inp[0]) ? node274 : node265;
										assign node265 = (inp[10]) ? node271 : node266;
											assign node266 = (inp[6]) ? node268 : 12'b000111111111;
												assign node268 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
											assign node271 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node274 = (inp[6]) ? node276 : 12'b000011111111;
											assign node276 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node279 = (inp[6]) ? node285 : node280;
										assign node280 = (inp[10]) ? node282 : 12'b000011111111;
											assign node282 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node285 = (inp[0]) ? node287 : 12'b000001111111;
											assign node287 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
								assign node290 = (inp[0]) ? node300 : node291;
									assign node291 = (inp[6]) ? node295 : node292;
										assign node292 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node295 = (inp[10]) ? 12'b000000111111 : node296;
											assign node296 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node300 = (inp[4]) ? node304 : node301;
										assign node301 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node304 = (inp[11]) ? 12'b000000011111 : node305;
											assign node305 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
						assign node309 = (inp[11]) ? node355 : node310;
							assign node310 = (inp[4]) ? node338 : node311;
								assign node311 = (inp[1]) ? node329 : node312;
									assign node312 = (inp[0]) ? node320 : node313;
										assign node313 = (inp[6]) ? node315 : 12'b001111111111;
											assign node315 = (inp[9]) ? 12'b000011111111 : node316;
												assign node316 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
										assign node320 = (inp[6]) ? 12'b000001111111 : node321;
											assign node321 = (inp[9]) ? node325 : node322;
												assign node322 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
												assign node325 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
									assign node329 = (inp[6]) ? 12'b000001111111 : node330;
										assign node330 = (inp[0]) ? node332 : 12'b000011111111;
											assign node332 = (inp[10]) ? 12'b000001111111 : node333;
												assign node333 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node338 = (inp[0]) ? node344 : node339;
									assign node339 = (inp[9]) ? 12'b000001111111 : node340;
										assign node340 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
									assign node344 = (inp[10]) ? node352 : node345;
										assign node345 = (inp[6]) ? 12'b000000111111 : node346;
											assign node346 = (inp[9]) ? node348 : 12'b000001111111;
												assign node348 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node352 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
							assign node355 = (inp[10]) ? node385 : node356;
								assign node356 = (inp[0]) ? node368 : node357;
									assign node357 = (inp[1]) ? node365 : node358;
										assign node358 = (inp[9]) ? 12'b000011111111 : node359;
											assign node359 = (inp[6]) ? 12'b000011111111 : node360;
												assign node360 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
										assign node365 = (inp[4]) ? 12'b000000111111 : 12'b000011111111;
									assign node368 = (inp[9]) ? node378 : node369;
										assign node369 = (inp[4]) ? node373 : node370;
											assign node370 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
											assign node373 = (inp[1]) ? 12'b000000111111 : node374;
												assign node374 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node378 = (inp[1]) ? node380 : 12'b000000111111;
											assign node380 = (inp[4]) ? node382 : 12'b000000111111;
												assign node382 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
								assign node385 = (inp[6]) ? node397 : node386;
									assign node386 = (inp[9]) ? node390 : node387;
										assign node387 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node390 = (inp[0]) ? node392 : 12'b000000111111;
											assign node392 = (inp[1]) ? 12'b000000011111 : node393;
												assign node393 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
									assign node397 = (inp[1]) ? node405 : node398;
										assign node398 = (inp[0]) ? node400 : 12'b000000111111;
											assign node400 = (inp[4]) ? 12'b000000011111 : node401;
												assign node401 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
										assign node405 = (inp[4]) ? 12'b000000001111 : node406;
											assign node406 = (inp[0]) ? 12'b000000001111 : 12'b000000111111;
				assign node410 = (inp[11]) ? node620 : node411;
					assign node411 = (inp[6]) ? node513 : node412;
						assign node412 = (inp[9]) ? node466 : node413;
							assign node413 = (inp[0]) ? node435 : node414;
								assign node414 = (inp[1]) ? node424 : node415;
									assign node415 = (inp[4]) ? 12'b000111111111 : node416;
										assign node416 = (inp[5]) ? node418 : 12'b001111111111;
											assign node418 = (inp[10]) ? 12'b000111111111 : node419;
												assign node419 = (inp[8]) ? 12'b000111111111 : 12'b001111111111;
									assign node424 = (inp[8]) ? node432 : node425;
										assign node425 = (inp[10]) ? 12'b000011111111 : node426;
											assign node426 = (inp[4]) ? 12'b000111111111 : node427;
												assign node427 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
										assign node432 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
								assign node435 = (inp[8]) ? node455 : node436;
									assign node436 = (inp[4]) ? node442 : node437;
										assign node437 = (inp[5]) ? node439 : 12'b001111111111;
											assign node439 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
										assign node442 = (inp[10]) ? node450 : node443;
											assign node443 = (inp[1]) ? node447 : node444;
												assign node444 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
												assign node447 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
											assign node450 = (inp[5]) ? 12'b000001111111 : node451;
												assign node451 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
									assign node455 = (inp[4]) ? node463 : node456;
										assign node456 = (inp[5]) ? 12'b000001111111 : node457;
											assign node457 = (inp[10]) ? node459 : 12'b000011111111;
												assign node459 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
										assign node463 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
							assign node466 = (inp[1]) ? node494 : node467;
								assign node467 = (inp[10]) ? node483 : node468;
									assign node468 = (inp[0]) ? node476 : node469;
										assign node469 = (inp[8]) ? 12'b000011111111 : node470;
											assign node470 = (inp[4]) ? node472 : 12'b000111111111;
												assign node472 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
										assign node476 = (inp[8]) ? node478 : 12'b000011111111;
											assign node478 = (inp[5]) ? 12'b000001111111 : node479;
												assign node479 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node483 = (inp[4]) ? node487 : node484;
										assign node484 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
										assign node487 = (inp[0]) ? node489 : 12'b000001111111;
											assign node489 = (inp[8]) ? 12'b000000111111 : node490;
												assign node490 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
								assign node494 = (inp[0]) ? node506 : node495;
									assign node495 = (inp[4]) ? node501 : node496;
										assign node496 = (inp[5]) ? 12'b000001111111 : node497;
											assign node497 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
										assign node501 = (inp[5]) ? node503 : 12'b000001111111;
											assign node503 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
									assign node506 = (inp[5]) ? node510 : node507;
										assign node507 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node510 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
						assign node513 = (inp[10]) ? node565 : node514;
							assign node514 = (inp[0]) ? node540 : node515;
								assign node515 = (inp[1]) ? node527 : node516;
									assign node516 = (inp[5]) ? node524 : node517;
										assign node517 = (inp[9]) ? 12'b000011111111 : node518;
											assign node518 = (inp[8]) ? node520 : 12'b000111111111;
												assign node520 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
										assign node524 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node527 = (inp[5]) ? node531 : node528;
										assign node528 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node531 = (inp[9]) ? node537 : node532;
											assign node532 = (inp[8]) ? 12'b000001111111 : node533;
												assign node533 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
											assign node537 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node540 = (inp[9]) ? node556 : node541;
									assign node541 = (inp[5]) ? node553 : node542;
										assign node542 = (inp[4]) ? node548 : node543;
											assign node543 = (inp[1]) ? node545 : 12'b000011111111;
												assign node545 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
											assign node548 = (inp[1]) ? 12'b000001111111 : node549;
												assign node549 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
										assign node553 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
									assign node556 = (inp[4]) ? node560 : node557;
										assign node557 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node560 = (inp[8]) ? node562 : 12'b000000111111;
											assign node562 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
							assign node565 = (inp[4]) ? node597 : node566;
								assign node566 = (inp[5]) ? node578 : node567;
									assign node567 = (inp[1]) ? node573 : node568;
										assign node568 = (inp[8]) ? 12'b000001111111 : node569;
											assign node569 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node573 = (inp[0]) ? node575 : 12'b000001111111;
											assign node575 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node578 = (inp[9]) ? node590 : node579;
										assign node579 = (inp[8]) ? node585 : node580;
											assign node580 = (inp[0]) ? 12'b000001111111 : node581;
												assign node581 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
											assign node585 = (inp[0]) ? 12'b000000111111 : node586;
												assign node586 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node590 = (inp[8]) ? node592 : 12'b000000111111;
											assign node592 = (inp[0]) ? node594 : 12'b000000111111;
												assign node594 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
								assign node597 = (inp[5]) ? node609 : node598;
									assign node598 = (inp[9]) ? node604 : node599;
										assign node599 = (inp[1]) ? 12'b000000111111 : node600;
											assign node600 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node604 = (inp[1]) ? node606 : 12'b000000111111;
											assign node606 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
									assign node609 = (inp[0]) ? node613 : node610;
										assign node610 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node613 = (inp[8]) ? 12'b000000001111 : node614;
											assign node614 = (inp[1]) ? node616 : 12'b000000011111;
												assign node616 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
					assign node620 = (inp[9]) ? node732 : node621;
						assign node621 = (inp[6]) ? node683 : node622;
							assign node622 = (inp[5]) ? node660 : node623;
								assign node623 = (inp[0]) ? node641 : node624;
									assign node624 = (inp[8]) ? node636 : node625;
										assign node625 = (inp[10]) ? node631 : node626;
											assign node626 = (inp[1]) ? node628 : 12'b000111111111;
												assign node628 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
											assign node631 = (inp[1]) ? 12'b000011111111 : node632;
												assign node632 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
										assign node636 = (inp[1]) ? node638 : 12'b000011111111;
											assign node638 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node641 = (inp[4]) ? node653 : node642;
										assign node642 = (inp[8]) ? node648 : node643;
											assign node643 = (inp[1]) ? 12'b000011111111 : node644;
												assign node644 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
											assign node648 = (inp[1]) ? 12'b000001111111 : node649;
												assign node649 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
										assign node653 = (inp[1]) ? node655 : 12'b000001111111;
											assign node655 = (inp[10]) ? 12'b000000111111 : node656;
												assign node656 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node660 = (inp[8]) ? node672 : node661;
									assign node661 = (inp[4]) ? node667 : node662;
										assign node662 = (inp[1]) ? 12'b000001111111 : node663;
											assign node663 = (inp[0]) ? 12'b000011111111 : 12'b000111111111;
										assign node667 = (inp[1]) ? node669 : 12'b000001111111;
											assign node669 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
									assign node672 = (inp[1]) ? node678 : node673;
										assign node673 = (inp[10]) ? 12'b000000111111 : node674;
											assign node674 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node678 = (inp[10]) ? node680 : 12'b000000111111;
											assign node680 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
							assign node683 = (inp[10]) ? node707 : node684;
								assign node684 = (inp[0]) ? node690 : node685;
									assign node685 = (inp[1]) ? 12'b000001111111 : node686;
										assign node686 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node690 = (inp[5]) ? node696 : node691;
										assign node691 = (inp[8]) ? 12'b000000111111 : node692;
											assign node692 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node696 = (inp[4]) ? node702 : node697;
											assign node697 = (inp[1]) ? 12'b000000111111 : node698;
												assign node698 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
											assign node702 = (inp[1]) ? 12'b000000011111 : node703;
												assign node703 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
								assign node707 = (inp[0]) ? node725 : node708;
									assign node708 = (inp[5]) ? node720 : node709;
										assign node709 = (inp[1]) ? node715 : node710;
											assign node710 = (inp[8]) ? node712 : 12'b000001111111;
												assign node712 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
											assign node715 = (inp[4]) ? 12'b000000111111 : node716;
												assign node716 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
										assign node720 = (inp[8]) ? node722 : 12'b000000111111;
											assign node722 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
									assign node725 = (inp[8]) ? node729 : node726;
										assign node726 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
										assign node729 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
						assign node732 = (inp[8]) ? node786 : node733;
							assign node733 = (inp[1]) ? node757 : node734;
								assign node734 = (inp[10]) ? node748 : node735;
									assign node735 = (inp[4]) ? node743 : node736;
										assign node736 = (inp[0]) ? 12'b000001111111 : node737;
											assign node737 = (inp[6]) ? 12'b000011111111 : node738;
												assign node738 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
										assign node743 = (inp[5]) ? node745 : 12'b000001111111;
											assign node745 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
									assign node748 = (inp[5]) ? node752 : node749;
										assign node749 = (inp[6]) ? 12'b000000111111 : 12'b000011111111;
										assign node752 = (inp[6]) ? 12'b000000011111 : node753;
											assign node753 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
								assign node757 = (inp[6]) ? node773 : node758;
									assign node758 = (inp[4]) ? node762 : node759;
										assign node759 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node762 = (inp[5]) ? node768 : node763;
											assign node763 = (inp[10]) ? node765 : 12'b000000111111;
												assign node765 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
											assign node768 = (inp[10]) ? 12'b000000011111 : node769;
												assign node769 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node773 = (inp[10]) ? node781 : node774;
										assign node774 = (inp[4]) ? 12'b000000011111 : node775;
											assign node775 = (inp[0]) ? node777 : 12'b000000111111;
												assign node777 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node781 = (inp[5]) ? 12'b000000001111 : node782;
											assign node782 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
							assign node786 = (inp[5]) ? node812 : node787;
								assign node787 = (inp[6]) ? node799 : node788;
									assign node788 = (inp[4]) ? node792 : node789;
										assign node789 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node792 = (inp[10]) ? 12'b000000011111 : node793;
											assign node793 = (inp[1]) ? node795 : 12'b000000111111;
												assign node795 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node799 = (inp[0]) ? node805 : node800;
										assign node800 = (inp[4]) ? 12'b000000011111 : node801;
											assign node801 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
										assign node805 = (inp[10]) ? node807 : 12'b000000011111;
											assign node807 = (inp[1]) ? node809 : 12'b000000011111;
												assign node809 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
								assign node812 = (inp[0]) ? node822 : node813;
									assign node813 = (inp[4]) ? node817 : node814;
										assign node814 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
										assign node817 = (inp[1]) ? node819 : 12'b000000011111;
											assign node819 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
									assign node822 = (inp[10]) ? node830 : node823;
										assign node823 = (inp[4]) ? node825 : 12'b000000011111;
											assign node825 = (inp[6]) ? 12'b000000001111 : node826;
												assign node826 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
										assign node830 = (inp[4]) ? node832 : 12'b000000001111;
											assign node832 = (inp[6]) ? 12'b000000000011 : 12'b000000000111;
			assign node835 = (inp[10]) ? node1285 : node836;
				assign node836 = (inp[6]) ? node1056 : node837;
					assign node837 = (inp[7]) ? node947 : node838;
						assign node838 = (inp[4]) ? node894 : node839;
							assign node839 = (inp[5]) ? node857 : node840;
								assign node840 = (inp[0]) ? node850 : node841;
									assign node841 = (inp[8]) ? node847 : node842;
										assign node842 = (inp[9]) ? 12'b000111111111 : node843;
											assign node843 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
										assign node847 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
									assign node850 = (inp[9]) ? 12'b000001111111 : node851;
										assign node851 = (inp[1]) ? 12'b000011111111 : node852;
											assign node852 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
								assign node857 = (inp[1]) ? node879 : node858;
									assign node858 = (inp[9]) ? node872 : node859;
										assign node859 = (inp[11]) ? node865 : node860;
											assign node860 = (inp[0]) ? 12'b000111111111 : node861;
												assign node861 = (inp[8]) ? 12'b000111111111 : 12'b001111111111;
											assign node865 = (inp[8]) ? node869 : node866;
												assign node866 = (inp[0]) ? 12'b000011111111 : 12'b000111111111;
												assign node869 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node872 = (inp[0]) ? node874 : 12'b000011111111;
											assign node874 = (inp[8]) ? 12'b000001111111 : node875;
												assign node875 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
									assign node879 = (inp[11]) ? node885 : node880;
										assign node880 = (inp[9]) ? node882 : 12'b000011111111;
											assign node882 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node885 = (inp[8]) ? node889 : node886;
											assign node886 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
											assign node889 = (inp[9]) ? 12'b000000111111 : node890;
												assign node890 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
							assign node894 = (inp[11]) ? node922 : node895;
								assign node895 = (inp[0]) ? node907 : node896;
									assign node896 = (inp[8]) ? node904 : node897;
										assign node897 = (inp[5]) ? 12'b000011111111 : node898;
											assign node898 = (inp[1]) ? node900 : 12'b000111111111;
												assign node900 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node904 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node907 = (inp[9]) ? node911 : node908;
										assign node908 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
										assign node911 = (inp[1]) ? node917 : node912;
											assign node912 = (inp[8]) ? 12'b000001111111 : node913;
												assign node913 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
											assign node917 = (inp[5]) ? 12'b000000111111 : node918;
												assign node918 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node922 = (inp[1]) ? node938 : node923;
									assign node923 = (inp[8]) ? node931 : node924;
										assign node924 = (inp[5]) ? node926 : 12'b000011111111;
											assign node926 = (inp[0]) ? 12'b000001111111 : node927;
												assign node927 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node931 = (inp[0]) ? node933 : 12'b000001111111;
											assign node933 = (inp[9]) ? node935 : 12'b000001111111;
												assign node935 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node938 = (inp[0]) ? node944 : node939;
										assign node939 = (inp[8]) ? 12'b000000111111 : node940;
											assign node940 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node944 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
						assign node947 = (inp[8]) ? node1009 : node948;
							assign node948 = (inp[9]) ? node974 : node949;
								assign node949 = (inp[1]) ? node965 : node950;
									assign node950 = (inp[5]) ? node958 : node951;
										assign node951 = (inp[4]) ? 12'b000011111111 : node952;
											assign node952 = (inp[11]) ? 12'b000111111111 : node953;
												assign node953 = (inp[0]) ? 12'b000111111111 : 12'b001111111111;
										assign node958 = (inp[11]) ? node960 : 12'b000011111111;
											assign node960 = (inp[4]) ? 12'b000001111111 : node961;
												assign node961 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
									assign node965 = (inp[11]) ? 12'b000000111111 : node966;
										assign node966 = (inp[5]) ? 12'b000001111111 : node967;
											assign node967 = (inp[4]) ? node969 : 12'b000011111111;
												assign node969 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node974 = (inp[5]) ? node992 : node975;
									assign node975 = (inp[0]) ? node987 : node976;
										assign node976 = (inp[1]) ? node982 : node977;
											assign node977 = (inp[11]) ? node979 : 12'b000011111111;
												assign node979 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
											assign node982 = (inp[4]) ? node984 : 12'b000001111111;
												assign node984 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node987 = (inp[11]) ? node989 : 12'b000001111111;
											assign node989 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
									assign node992 = (inp[0]) ? node1002 : node993;
										assign node993 = (inp[4]) ? node997 : node994;
											assign node994 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
											assign node997 = (inp[1]) ? 12'b000000111111 : node998;
												assign node998 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1002 = (inp[11]) ? 12'b000000011111 : node1003;
											assign node1003 = (inp[4]) ? node1005 : 12'b000000111111;
												assign node1005 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
							assign node1009 = (inp[0]) ? node1027 : node1010;
								assign node1010 = (inp[9]) ? 12'b000000111111 : node1011;
									assign node1011 = (inp[11]) ? node1019 : node1012;
										assign node1012 = (inp[1]) ? 12'b000001111111 : node1013;
											assign node1013 = (inp[5]) ? node1015 : 12'b000011111111;
												assign node1015 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node1019 = (inp[5]) ? 12'b000000011111 : node1020;
											assign node1020 = (inp[4]) ? node1022 : 12'b000001111111;
												assign node1022 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node1027 = (inp[1]) ? node1039 : node1028;
									assign node1028 = (inp[5]) ? node1034 : node1029;
										assign node1029 = (inp[4]) ? 12'b000000111111 : node1030;
											assign node1030 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node1034 = (inp[11]) ? node1036 : 12'b000000111111;
											assign node1036 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node1039 = (inp[4]) ? node1049 : node1040;
										assign node1040 = (inp[5]) ? node1044 : node1041;
											assign node1041 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
											assign node1044 = (inp[9]) ? 12'b000000011111 : node1045;
												assign node1045 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node1049 = (inp[5]) ? node1051 : 12'b000000011111;
											assign node1051 = (inp[11]) ? node1053 : 12'b000000011111;
												assign node1053 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
					assign node1056 = (inp[5]) ? node1166 : node1057;
						assign node1057 = (inp[8]) ? node1111 : node1058;
							assign node1058 = (inp[4]) ? node1080 : node1059;
								assign node1059 = (inp[0]) ? node1075 : node1060;
									assign node1060 = (inp[7]) ? node1072 : node1061;
										assign node1061 = (inp[11]) ? node1067 : node1062;
											assign node1062 = (inp[9]) ? node1064 : 12'b000111111111;
												assign node1064 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
											assign node1067 = (inp[1]) ? 12'b000011111111 : node1068;
												assign node1068 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node1072 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
									assign node1075 = (inp[11]) ? 12'b000001111111 : node1076;
										assign node1076 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
								assign node1080 = (inp[11]) ? node1094 : node1081;
									assign node1081 = (inp[7]) ? node1089 : node1082;
										assign node1082 = (inp[0]) ? 12'b000001111111 : node1083;
											assign node1083 = (inp[1]) ? 12'b000011111111 : node1084;
												assign node1084 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node1089 = (inp[9]) ? node1091 : 12'b000001111111;
											assign node1091 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node1094 = (inp[0]) ? node1104 : node1095;
										assign node1095 = (inp[9]) ? 12'b000000111111 : node1096;
											assign node1096 = (inp[7]) ? node1100 : node1097;
												assign node1097 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
												assign node1100 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node1104 = (inp[7]) ? 12'b000000011111 : node1105;
											assign node1105 = (inp[9]) ? node1107 : 12'b000000111111;
												assign node1107 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
							assign node1111 = (inp[9]) ? node1135 : node1112;
								assign node1112 = (inp[0]) ? node1120 : node1113;
									assign node1113 = (inp[4]) ? 12'b000001111111 : node1114;
										assign node1114 = (inp[1]) ? node1116 : 12'b000011111111;
											assign node1116 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
									assign node1120 = (inp[7]) ? node1128 : node1121;
										assign node1121 = (inp[1]) ? 12'b000000111111 : node1122;
											assign node1122 = (inp[4]) ? 12'b000001111111 : node1123;
												assign node1123 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node1128 = (inp[4]) ? 12'b000000011111 : node1129;
											assign node1129 = (inp[11]) ? node1131 : 12'b000001111111;
												assign node1131 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
								assign node1135 = (inp[7]) ? node1147 : node1136;
									assign node1136 = (inp[4]) ? node1140 : node1137;
										assign node1137 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node1140 = (inp[11]) ? node1142 : 12'b000000111111;
											assign node1142 = (inp[0]) ? 12'b000000011111 : node1143;
												assign node1143 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node1147 = (inp[0]) ? node1159 : node1148;
										assign node1148 = (inp[4]) ? node1154 : node1149;
											assign node1149 = (inp[11]) ? node1151 : 12'b000000111111;
												assign node1151 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
											assign node1154 = (inp[11]) ? node1156 : 12'b000000011111;
												assign node1156 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
										assign node1159 = (inp[11]) ? node1161 : 12'b000000011111;
											assign node1161 = (inp[4]) ? 12'b000000001111 : node1162;
												assign node1162 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
						assign node1166 = (inp[1]) ? node1236 : node1167;
							assign node1167 = (inp[8]) ? node1205 : node1168;
								assign node1168 = (inp[11]) ? node1190 : node1169;
									assign node1169 = (inp[4]) ? node1179 : node1170;
										assign node1170 = (inp[7]) ? node1174 : node1171;
											assign node1171 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
											assign node1174 = (inp[9]) ? node1176 : 12'b000001111111;
												assign node1176 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node1179 = (inp[9]) ? node1185 : node1180;
											assign node1180 = (inp[7]) ? node1182 : 12'b000001111111;
												assign node1182 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
											assign node1185 = (inp[0]) ? 12'b000000111111 : node1186;
												assign node1186 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
									assign node1190 = (inp[0]) ? node1198 : node1191;
										assign node1191 = (inp[7]) ? 12'b000000111111 : node1192;
											assign node1192 = (inp[9]) ? node1194 : 12'b000001111111;
												assign node1194 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1198 = (inp[9]) ? node1200 : 12'b000000111111;
											assign node1200 = (inp[4]) ? node1202 : 12'b000000011111;
												assign node1202 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
								assign node1205 = (inp[9]) ? node1219 : node1206;
									assign node1206 = (inp[4]) ? node1214 : node1207;
										assign node1207 = (inp[11]) ? 12'b000000111111 : node1208;
											assign node1208 = (inp[0]) ? node1210 : 12'b000001111111;
												assign node1210 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
										assign node1214 = (inp[0]) ? 12'b000000001111 : node1215;
											assign node1215 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node1219 = (inp[0]) ? node1231 : node1220;
										assign node1220 = (inp[11]) ? node1226 : node1221;
											assign node1221 = (inp[7]) ? node1223 : 12'b000000111111;
												assign node1223 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
											assign node1226 = (inp[7]) ? node1228 : 12'b000000011111;
												assign node1228 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node1231 = (inp[7]) ? node1233 : 12'b000000011111;
											assign node1233 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
							assign node1236 = (inp[4]) ? node1260 : node1237;
								assign node1237 = (inp[9]) ? node1251 : node1238;
									assign node1238 = (inp[8]) ? node1244 : node1239;
										assign node1239 = (inp[0]) ? node1241 : 12'b000001111111;
											assign node1241 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node1244 = (inp[11]) ? node1246 : 12'b000000111111;
											assign node1246 = (inp[0]) ? 12'b000000011111 : node1247;
												assign node1247 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node1251 = (inp[11]) ? node1255 : node1252;
										assign node1252 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node1255 = (inp[0]) ? node1257 : 12'b000000011111;
											assign node1257 = (inp[8]) ? 12'b000000000111 : 12'b000000001111;
								assign node1260 = (inp[9]) ? node1266 : node1261;
									assign node1261 = (inp[8]) ? node1263 : 12'b000000011111;
										assign node1263 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node1266 = (inp[11]) ? node1280 : node1267;
										assign node1267 = (inp[0]) ? node1273 : node1268;
											assign node1268 = (inp[8]) ? node1270 : 12'b000000011111;
												assign node1270 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
											assign node1273 = (inp[7]) ? node1277 : node1274;
												assign node1274 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
												assign node1277 = (inp[8]) ? 12'b000000000111 : 12'b000000001111;
										assign node1280 = (inp[8]) ? node1282 : 12'b000000001111;
											assign node1282 = (inp[7]) ? 12'b000000000011 : 12'b000000000111;
				assign node1285 = (inp[9]) ? node1489 : node1286;
					assign node1286 = (inp[5]) ? node1400 : node1287;
						assign node1287 = (inp[1]) ? node1337 : node1288;
							assign node1288 = (inp[4]) ? node1310 : node1289;
								assign node1289 = (inp[6]) ? node1305 : node1290;
									assign node1290 = (inp[8]) ? node1298 : node1291;
										assign node1291 = (inp[0]) ? node1293 : 12'b000111111111;
											assign node1293 = (inp[11]) ? 12'b000011111111 : node1294;
												assign node1294 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
										assign node1298 = (inp[0]) ? node1300 : 12'b000011111111;
											assign node1300 = (inp[11]) ? 12'b000001111111 : node1301;
												assign node1301 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
									assign node1305 = (inp[8]) ? 12'b000001111111 : node1306;
										assign node1306 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node1310 = (inp[8]) ? node1322 : node1311;
									assign node1311 = (inp[7]) ? node1313 : 12'b000011111111;
										assign node1313 = (inp[0]) ? 12'b000000111111 : node1314;
											assign node1314 = (inp[6]) ? node1318 : node1315;
												assign node1315 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
												assign node1318 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node1322 = (inp[0]) ? node1330 : node1323;
										assign node1323 = (inp[6]) ? 12'b000000111111 : node1324;
											assign node1324 = (inp[11]) ? node1326 : 12'b000001111111;
												assign node1326 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
										assign node1330 = (inp[7]) ? node1332 : 12'b000000111111;
											assign node1332 = (inp[6]) ? 12'b000000011111 : node1333;
												assign node1333 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node1337 = (inp[6]) ? node1371 : node1338;
								assign node1338 = (inp[7]) ? node1358 : node1339;
									assign node1339 = (inp[11]) ? node1351 : node1340;
										assign node1340 = (inp[0]) ? node1346 : node1341;
											assign node1341 = (inp[4]) ? node1343 : 12'b000011111111;
												assign node1343 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
											assign node1346 = (inp[8]) ? node1348 : 12'b000001111111;
												assign node1348 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1351 = (inp[4]) ? 12'b000000111111 : node1352;
											assign node1352 = (inp[0]) ? node1354 : 12'b000001111111;
												assign node1354 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
									assign node1358 = (inp[0]) ? node1366 : node1359;
										assign node1359 = (inp[8]) ? 12'b000000111111 : node1360;
											assign node1360 = (inp[11]) ? node1362 : 12'b000001111111;
												assign node1362 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1366 = (inp[11]) ? node1368 : 12'b000000111111;
											assign node1368 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node1371 = (inp[7]) ? node1387 : node1372;
									assign node1372 = (inp[4]) ? node1382 : node1373;
										assign node1373 = (inp[11]) ? node1375 : 12'b000001111111;
											assign node1375 = (inp[8]) ? node1379 : node1376;
												assign node1376 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
												assign node1379 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node1382 = (inp[0]) ? node1384 : 12'b000000111111;
											assign node1384 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1387 = (inp[4]) ? node1397 : node1388;
										assign node1388 = (inp[11]) ? node1392 : node1389;
											assign node1389 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
											assign node1392 = (inp[8]) ? node1394 : 12'b000000011111;
												assign node1394 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
										assign node1397 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
						assign node1400 = (inp[0]) ? node1446 : node1401;
							assign node1401 = (inp[11]) ? node1425 : node1402;
								assign node1402 = (inp[1]) ? node1418 : node1403;
									assign node1403 = (inp[7]) ? node1411 : node1404;
										assign node1404 = (inp[4]) ? node1406 : 12'b000011111111;
											assign node1406 = (inp[6]) ? node1408 : 12'b000001111111;
												assign node1408 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
										assign node1411 = (inp[4]) ? 12'b000000111111 : node1412;
											assign node1412 = (inp[8]) ? node1414 : 12'b000001111111;
												assign node1414 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
									assign node1418 = (inp[8]) ? node1422 : node1419;
										assign node1419 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node1422 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
								assign node1425 = (inp[7]) ? node1435 : node1426;
									assign node1426 = (inp[8]) ? node1432 : node1427;
										assign node1427 = (inp[6]) ? node1429 : 12'b000011111111;
											assign node1429 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node1432 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node1435 = (inp[6]) ? node1439 : node1436;
										assign node1436 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node1439 = (inp[4]) ? node1441 : 12'b000000011111;
											assign node1441 = (inp[1]) ? 12'b000000001111 : node1442;
												assign node1442 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
							assign node1446 = (inp[8]) ? node1466 : node1447;
								assign node1447 = (inp[1]) ? node1455 : node1448;
									assign node1448 = (inp[11]) ? 12'b000000111111 : node1449;
										assign node1449 = (inp[6]) ? 12'b000000111111 : node1450;
											assign node1450 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
									assign node1455 = (inp[11]) ? node1463 : node1456;
										assign node1456 = (inp[6]) ? 12'b000000011111 : node1457;
											assign node1457 = (inp[4]) ? node1459 : 12'b000000111111;
												assign node1459 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node1463 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
								assign node1466 = (inp[11]) ? node1480 : node1467;
									assign node1467 = (inp[1]) ? node1475 : node1468;
										assign node1468 = (inp[6]) ? node1470 : 12'b000000011111;
											assign node1470 = (inp[4]) ? node1472 : 12'b000000011111;
												assign node1472 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node1475 = (inp[4]) ? 12'b000000001111 : node1476;
											assign node1476 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
									assign node1480 = (inp[4]) ? node1484 : node1481;
										assign node1481 = (inp[6]) ? 12'b000000001111 : 12'b000000111111;
										assign node1484 = (inp[6]) ? 12'b000000000111 : node1485;
											assign node1485 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
					assign node1489 = (inp[0]) ? node1611 : node1490;
						assign node1490 = (inp[1]) ? node1562 : node1491;
							assign node1491 = (inp[6]) ? node1521 : node1492;
								assign node1492 = (inp[7]) ? node1506 : node1493;
									assign node1493 = (inp[8]) ? node1501 : node1494;
										assign node1494 = (inp[4]) ? node1496 : 12'b000011111111;
											assign node1496 = (inp[5]) ? 12'b000001111111 : node1497;
												assign node1497 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node1501 = (inp[5]) ? node1503 : 12'b000001111111;
											assign node1503 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node1506 = (inp[5]) ? node1518 : node1507;
										assign node1507 = (inp[4]) ? node1513 : node1508;
											assign node1508 = (inp[11]) ? 12'b000001111111 : node1509;
												assign node1509 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
											assign node1513 = (inp[11]) ? 12'b000000111111 : node1514;
												assign node1514 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
										assign node1518 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
								assign node1521 = (inp[7]) ? node1537 : node1522;
									assign node1522 = (inp[4]) ? node1530 : node1523;
										assign node1523 = (inp[5]) ? node1525 : 12'b000001111111;
											assign node1525 = (inp[8]) ? 12'b000000111111 : node1526;
												assign node1526 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1530 = (inp[8]) ? 12'b000000011111 : node1531;
											assign node1531 = (inp[5]) ? node1533 : 12'b000000111111;
												assign node1533 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node1537 = (inp[8]) ? node1551 : node1538;
										assign node1538 = (inp[5]) ? node1546 : node1539;
											assign node1539 = (inp[4]) ? node1543 : node1540;
												assign node1540 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
												assign node1543 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
											assign node1546 = (inp[11]) ? node1548 : 12'b000000011111;
												assign node1548 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node1551 = (inp[4]) ? node1557 : node1552;
											assign node1552 = (inp[5]) ? node1554 : 12'b000000011111;
												assign node1554 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
											assign node1557 = (inp[5]) ? node1559 : 12'b000000001111;
												assign node1559 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
							assign node1562 = (inp[4]) ? node1580 : node1563;
								assign node1563 = (inp[6]) ? node1565 : 12'b000000111111;
									assign node1565 = (inp[11]) ? node1573 : node1566;
										assign node1566 = (inp[8]) ? node1570 : node1567;
											assign node1567 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
											assign node1570 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node1573 = (inp[5]) ? 12'b000000001111 : node1574;
											assign node1574 = (inp[7]) ? node1576 : 12'b000000011111;
												assign node1576 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
								assign node1580 = (inp[5]) ? node1594 : node1581;
									assign node1581 = (inp[6]) ? node1589 : node1582;
										assign node1582 = (inp[8]) ? node1584 : 12'b000000111111;
											assign node1584 = (inp[11]) ? node1586 : 12'b000000011111;
												assign node1586 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node1589 = (inp[8]) ? 12'b000000001111 : node1590;
											assign node1590 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1594 = (inp[7]) ? node1604 : node1595;
										assign node1595 = (inp[6]) ? node1597 : 12'b000000011111;
											assign node1597 = (inp[11]) ? node1601 : node1598;
												assign node1598 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
												assign node1601 = (inp[8]) ? 12'b000000000111 : 12'b000000001111;
										assign node1604 = (inp[6]) ? 12'b000000000111 : node1605;
											assign node1605 = (inp[8]) ? node1607 : 12'b000000001111;
												assign node1607 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
						assign node1611 = (inp[6]) ? node1669 : node1612;
							assign node1612 = (inp[8]) ? node1648 : node1613;
								assign node1613 = (inp[5]) ? node1627 : node1614;
									assign node1614 = (inp[1]) ? node1620 : node1615;
										assign node1615 = (inp[11]) ? 12'b000000111111 : node1616;
											assign node1616 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
										assign node1620 = (inp[11]) ? node1622 : 12'b000000111111;
											assign node1622 = (inp[4]) ? 12'b000000001111 : node1623;
												assign node1623 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node1627 = (inp[1]) ? node1635 : node1628;
										assign node1628 = (inp[7]) ? 12'b000000011111 : node1629;
											assign node1629 = (inp[4]) ? node1631 : 12'b000000111111;
												assign node1631 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node1635 = (inp[11]) ? node1641 : node1636;
											assign node1636 = (inp[7]) ? node1638 : 12'b000000011111;
												assign node1638 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
											assign node1641 = (inp[7]) ? node1645 : node1642;
												assign node1642 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
												assign node1645 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
								assign node1648 = (inp[4]) ? node1656 : node1649;
									assign node1649 = (inp[7]) ? node1651 : 12'b000000011111;
										assign node1651 = (inp[11]) ? node1653 : 12'b000000011111;
											assign node1653 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
									assign node1656 = (inp[5]) ? node1662 : node1657;
										assign node1657 = (inp[7]) ? 12'b000000001111 : node1658;
											assign node1658 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
										assign node1662 = (inp[11]) ? node1664 : 12'b000000011111;
											assign node1664 = (inp[7]) ? 12'b000000000111 : node1665;
												assign node1665 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
							assign node1669 = (inp[7]) ? node1691 : node1670;
								assign node1670 = (inp[1]) ? node1684 : node1671;
									assign node1671 = (inp[11]) ? node1677 : node1672;
										assign node1672 = (inp[4]) ? 12'b000000011111 : node1673;
											assign node1673 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node1677 = (inp[4]) ? 12'b000000001111 : node1678;
											assign node1678 = (inp[5]) ? node1680 : 12'b000000011111;
												assign node1680 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
									assign node1684 = (inp[5]) ? node1688 : node1685;
										assign node1685 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node1688 = (inp[8]) ? 12'b000000000111 : 12'b000000001111;
								assign node1691 = (inp[4]) ? node1701 : node1692;
									assign node1692 = (inp[1]) ? node1694 : 12'b000000001111;
										assign node1694 = (inp[8]) ? 12'b000000000111 : node1695;
											assign node1695 = (inp[5]) ? node1697 : 12'b000000001111;
												assign node1697 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
									assign node1701 = (inp[8]) ? node1705 : node1702;
										assign node1702 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
										assign node1705 = (inp[1]) ? 12'b000000000011 : node1706;
											assign node1706 = (inp[11]) ? 12'b000000000011 : 12'b000000000111;
		assign node1710 = (inp[8]) ? node2602 : node1711;
			assign node1711 = (inp[10]) ? node2181 : node1712;
				assign node1712 = (inp[11]) ? node1946 : node1713;
					assign node1713 = (inp[4]) ? node1821 : node1714;
						assign node1714 = (inp[7]) ? node1776 : node1715;
							assign node1715 = (inp[1]) ? node1743 : node1716;
								assign node1716 = (inp[9]) ? node1732 : node1717;
									assign node1717 = (inp[5]) ? node1729 : node1718;
										assign node1718 = (inp[2]) ? node1724 : node1719;
											assign node1719 = (inp[6]) ? node1721 : 12'b001111111111;
												assign node1721 = (inp[0]) ? 12'b000111111111 : 12'b001111111111;
											assign node1724 = (inp[0]) ? 12'b000111111111 : node1725;
												assign node1725 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
										assign node1729 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
									assign node1732 = (inp[0]) ? node1740 : node1733;
										assign node1733 = (inp[5]) ? node1735 : 12'b000111111111;
											assign node1735 = (inp[6]) ? 12'b000011111111 : node1736;
												assign node1736 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
										assign node1740 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
								assign node1743 = (inp[2]) ? node1759 : node1744;
									assign node1744 = (inp[0]) ? node1754 : node1745;
										assign node1745 = (inp[6]) ? 12'b000011111111 : node1746;
											assign node1746 = (inp[5]) ? node1750 : node1747;
												assign node1747 = (inp[9]) ? 12'b000111111111 : 12'b001111111111;
												assign node1750 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node1754 = (inp[9]) ? node1756 : 12'b000011111111;
											assign node1756 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node1759 = (inp[9]) ? node1769 : node1760;
										assign node1760 = (inp[0]) ? node1764 : node1761;
											assign node1761 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
											assign node1764 = (inp[5]) ? 12'b000001111111 : node1765;
												assign node1765 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
										assign node1769 = (inp[6]) ? 12'b000000111111 : node1770;
											assign node1770 = (inp[0]) ? 12'b000001111111 : node1771;
												assign node1771 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
							assign node1776 = (inp[9]) ? node1800 : node1777;
								assign node1777 = (inp[0]) ? node1787 : node1778;
									assign node1778 = (inp[1]) ? node1784 : node1779;
										assign node1779 = (inp[6]) ? node1781 : 12'b000111111111;
											assign node1781 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node1784 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node1787 = (inp[5]) ? node1795 : node1788;
										assign node1788 = (inp[6]) ? node1790 : 12'b000011111111;
											assign node1790 = (inp[1]) ? 12'b000001111111 : node1791;
												assign node1791 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node1795 = (inp[1]) ? node1797 : 12'b000001111111;
											assign node1797 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
								assign node1800 = (inp[2]) ? 12'b000000111111 : node1801;
									assign node1801 = (inp[1]) ? node1813 : node1802;
										assign node1802 = (inp[6]) ? node1808 : node1803;
											assign node1803 = (inp[5]) ? node1805 : 12'b000011111111;
												assign node1805 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
											assign node1808 = (inp[5]) ? 12'b000001111111 : node1809;
												assign node1809 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node1813 = (inp[0]) ? node1815 : 12'b000001111111;
											assign node1815 = (inp[6]) ? 12'b000000111111 : node1816;
												assign node1816 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
						assign node1821 = (inp[0]) ? node1891 : node1822;
							assign node1822 = (inp[6]) ? node1864 : node1823;
								assign node1823 = (inp[5]) ? node1847 : node1824;
									assign node1824 = (inp[7]) ? node1836 : node1825;
										assign node1825 = (inp[2]) ? node1831 : node1826;
											assign node1826 = (inp[9]) ? 12'b000111111111 : node1827;
												assign node1827 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
											assign node1831 = (inp[9]) ? 12'b000001111111 : node1832;
												assign node1832 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
										assign node1836 = (inp[1]) ? node1842 : node1837;
											assign node1837 = (inp[2]) ? node1839 : 12'b000011111111;
												assign node1839 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
											assign node1842 = (inp[2]) ? 12'b000001111111 : node1843;
												assign node1843 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node1847 = (inp[2]) ? node1853 : node1848;
										assign node1848 = (inp[9]) ? 12'b000001111111 : node1849;
											assign node1849 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
										assign node1853 = (inp[1]) ? node1859 : node1854;
											assign node1854 = (inp[7]) ? 12'b000001111111 : node1855;
												assign node1855 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
											assign node1859 = (inp[7]) ? 12'b000000111111 : node1860;
												assign node1860 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
								assign node1864 = (inp[1]) ? node1878 : node1865;
									assign node1865 = (inp[9]) ? node1873 : node1866;
										assign node1866 = (inp[2]) ? 12'b000001111111 : node1867;
											assign node1867 = (inp[5]) ? 12'b000011111111 : node1868;
												assign node1868 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
										assign node1873 = (inp[7]) ? node1875 : 12'b000001111111;
											assign node1875 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
									assign node1878 = (inp[9]) ? node1884 : node1879;
										assign node1879 = (inp[5]) ? 12'b000000111111 : node1880;
											assign node1880 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node1884 = (inp[2]) ? 12'b000000011111 : node1885;
											assign node1885 = (inp[5]) ? node1887 : 12'b000000111111;
												assign node1887 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
							assign node1891 = (inp[6]) ? node1917 : node1892;
								assign node1892 = (inp[9]) ? node1904 : node1893;
									assign node1893 = (inp[2]) ? node1899 : node1894;
										assign node1894 = (inp[5]) ? node1896 : 12'b000011111111;
											assign node1896 = (inp[7]) ? 12'b000000111111 : 12'b000011111111;
										assign node1899 = (inp[5]) ? 12'b000000111111 : node1900;
											assign node1900 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node1904 = (inp[7]) ? node1912 : node1905;
										assign node1905 = (inp[5]) ? 12'b000000111111 : node1906;
											assign node1906 = (inp[2]) ? node1908 : 12'b000001111111;
												assign node1908 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node1912 = (inp[1]) ? node1914 : 12'b000000111111;
											assign node1914 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
								assign node1917 = (inp[1]) ? node1929 : node1918;
									assign node1918 = (inp[9]) ? node1926 : node1919;
										assign node1919 = (inp[2]) ? 12'b000000111111 : node1920;
											assign node1920 = (inp[5]) ? 12'b000000111111 : node1921;
												assign node1921 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
										assign node1926 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node1929 = (inp[5]) ? node1937 : node1930;
										assign node1930 = (inp[9]) ? 12'b000000011111 : node1931;
											assign node1931 = (inp[7]) ? node1933 : 12'b000000111111;
												assign node1933 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
										assign node1937 = (inp[9]) ? node1943 : node1938;
											assign node1938 = (inp[2]) ? node1940 : 12'b000000011111;
												assign node1940 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
											assign node1943 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
					assign node1946 = (inp[7]) ? node2054 : node1947;
						assign node1947 = (inp[2]) ? node1999 : node1948;
							assign node1948 = (inp[1]) ? node1976 : node1949;
								assign node1949 = (inp[0]) ? node1961 : node1950;
									assign node1950 = (inp[9]) ? node1958 : node1951;
										assign node1951 = (inp[4]) ? node1953 : 12'b000111111111;
											assign node1953 = (inp[6]) ? 12'b000011111111 : node1954;
												assign node1954 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
										assign node1958 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node1961 = (inp[5]) ? node1969 : node1962;
										assign node1962 = (inp[9]) ? node1964 : 12'b000011111111;
											assign node1964 = (inp[6]) ? 12'b000001111111 : node1965;
												assign node1965 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node1969 = (inp[6]) ? node1971 : 12'b000001111111;
											assign node1971 = (inp[9]) ? 12'b000000111111 : node1972;
												assign node1972 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
								assign node1976 = (inp[0]) ? node1988 : node1977;
									assign node1977 = (inp[6]) ? node1983 : node1978;
										assign node1978 = (inp[4]) ? node1980 : 12'b000011111111;
											assign node1980 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node1983 = (inp[5]) ? node1985 : 12'b000001111111;
											assign node1985 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node1988 = (inp[9]) ? node1992 : node1989;
										assign node1989 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1992 = (inp[5]) ? 12'b000000011111 : node1993;
											assign node1993 = (inp[6]) ? node1995 : 12'b000000111111;
												assign node1995 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
							assign node1999 = (inp[5]) ? node2025 : node2000;
								assign node2000 = (inp[6]) ? node2010 : node2001;
									assign node2001 = (inp[9]) ? 12'b000001111111 : node2002;
										assign node2002 = (inp[4]) ? node2004 : 12'b000011111111;
											assign node2004 = (inp[0]) ? 12'b000000111111 : node2005;
												assign node2005 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
									assign node2010 = (inp[9]) ? node2022 : node2011;
										assign node2011 = (inp[1]) ? node2017 : node2012;
											assign node2012 = (inp[0]) ? node2014 : 12'b000001111111;
												assign node2014 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
											assign node2017 = (inp[4]) ? 12'b000000111111 : node2018;
												assign node2018 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
										assign node2022 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node2025 = (inp[1]) ? node2039 : node2026;
									assign node2026 = (inp[4]) ? node2032 : node2027;
										assign node2027 = (inp[0]) ? 12'b000000111111 : node2028;
											assign node2028 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node2032 = (inp[0]) ? 12'b000000011111 : node2033;
											assign node2033 = (inp[6]) ? node2035 : 12'b000000111111;
												assign node2035 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node2039 = (inp[6]) ? node2049 : node2040;
										assign node2040 = (inp[4]) ? node2042 : 12'b000000111111;
											assign node2042 = (inp[9]) ? node2046 : node2043;
												assign node2043 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
												assign node2046 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
										assign node2049 = (inp[0]) ? 12'b000000001111 : node2050;
											assign node2050 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
						assign node2054 = (inp[9]) ? node2120 : node2055;
							assign node2055 = (inp[6]) ? node2083 : node2056;
								assign node2056 = (inp[5]) ? node2072 : node2057;
									assign node2057 = (inp[4]) ? node2069 : node2058;
										assign node2058 = (inp[0]) ? node2064 : node2059;
											assign node2059 = (inp[1]) ? node2061 : 12'b000011111111;
												assign node2061 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
											assign node2064 = (inp[2]) ? 12'b000001111111 : node2065;
												assign node2065 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
										assign node2069 = (inp[1]) ? 12'b000001111111 : 12'b000000111111;
									assign node2072 = (inp[0]) ? node2076 : node2073;
										assign node2073 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node2076 = (inp[4]) ? 12'b000000011111 : node2077;
											assign node2077 = (inp[1]) ? node2079 : 12'b000000111111;
												assign node2079 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
								assign node2083 = (inp[1]) ? node2099 : node2084;
									assign node2084 = (inp[0]) ? node2092 : node2085;
										assign node2085 = (inp[2]) ? 12'b000000111111 : node2086;
											assign node2086 = (inp[4]) ? node2088 : 12'b000001111111;
												assign node2088 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node2092 = (inp[2]) ? node2094 : 12'b000000111111;
											assign node2094 = (inp[5]) ? 12'b000000011111 : node2095;
												assign node2095 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
									assign node2099 = (inp[2]) ? node2111 : node2100;
										assign node2100 = (inp[0]) ? node2106 : node2101;
											assign node2101 = (inp[5]) ? 12'b000000111111 : node2102;
												assign node2102 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
											assign node2106 = (inp[5]) ? node2108 : 12'b000000011111;
												assign node2108 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node2111 = (inp[0]) ? node2117 : node2112;
											assign node2112 = (inp[5]) ? node2114 : 12'b000000011111;
												assign node2114 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
											assign node2117 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
							assign node2120 = (inp[0]) ? node2148 : node2121;
								assign node2121 = (inp[1]) ? node2133 : node2122;
									assign node2122 = (inp[4]) ? node2130 : node2123;
										assign node2123 = (inp[6]) ? 12'b000000111111 : node2124;
											assign node2124 = (inp[5]) ? node2126 : 12'b000001111111;
												assign node2126 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node2130 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node2133 = (inp[4]) ? 12'b000000001111 : node2134;
										assign node2134 = (inp[2]) ? node2140 : node2135;
											assign node2135 = (inp[5]) ? node2137 : 12'b000000111111;
												assign node2137 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
											assign node2140 = (inp[6]) ? node2144 : node2141;
												assign node2141 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
												assign node2144 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node2148 = (inp[6]) ? node2164 : node2149;
									assign node2149 = (inp[4]) ? node2157 : node2150;
										assign node2150 = (inp[2]) ? node2152 : 12'b000000111111;
											assign node2152 = (inp[5]) ? node2154 : 12'b000000111111;
												assign node2154 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
										assign node2157 = (inp[1]) ? 12'b000000001111 : node2158;
											assign node2158 = (inp[2]) ? node2160 : 12'b000000011111;
												assign node2160 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
									assign node2164 = (inp[4]) ? node2172 : node2165;
										assign node2165 = (inp[5]) ? node2167 : 12'b000000001111;
											assign node2167 = (inp[2]) ? node2169 : 12'b000000001111;
												assign node2169 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
										assign node2172 = (inp[2]) ? node2176 : node2173;
											assign node2173 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
											assign node2176 = (inp[1]) ? node2178 : 12'b000000000111;
												assign node2178 = (inp[5]) ? 12'b000000000011 : 12'b000000000111;
				assign node2181 = (inp[9]) ? node2371 : node2182;
					assign node2182 = (inp[1]) ? node2284 : node2183;
						assign node2183 = (inp[4]) ? node2227 : node2184;
							assign node2184 = (inp[6]) ? node2204 : node2185;
								assign node2185 = (inp[11]) ? node2195 : node2186;
									assign node2186 = (inp[7]) ? node2188 : 12'b000111111111;
										assign node2188 = (inp[5]) ? 12'b000001111111 : node2189;
											assign node2189 = (inp[0]) ? 12'b000001111111 : node2190;
												assign node2190 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
									assign node2195 = (inp[7]) ? node2199 : node2196;
										assign node2196 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node2199 = (inp[0]) ? node2201 : 12'b000001111111;
											assign node2201 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
								assign node2204 = (inp[0]) ? node2218 : node2205;
									assign node2205 = (inp[5]) ? node2211 : node2206;
										assign node2206 = (inp[11]) ? 12'b000001111111 : node2207;
											assign node2207 = (inp[7]) ? 12'b000001111111 : 12'b000111111111;
										assign node2211 = (inp[11]) ? 12'b000000011111 : node2212;
											assign node2212 = (inp[2]) ? node2214 : 12'b000001111111;
												assign node2214 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
									assign node2218 = (inp[7]) ? 12'b000000111111 : node2219;
										assign node2219 = (inp[11]) ? 12'b000000111111 : node2220;
											assign node2220 = (inp[5]) ? node2222 : 12'b000001111111;
												assign node2222 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
							assign node2227 = (inp[5]) ? node2255 : node2228;
								assign node2228 = (inp[6]) ? node2244 : node2229;
									assign node2229 = (inp[2]) ? node2241 : node2230;
										assign node2230 = (inp[7]) ? node2236 : node2231;
											assign node2231 = (inp[11]) ? 12'b000011111111 : node2232;
												assign node2232 = (inp[0]) ? 12'b000011111111 : 12'b000111111111;
											assign node2236 = (inp[11]) ? 12'b000001111111 : node2237;
												assign node2237 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
										assign node2241 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node2244 = (inp[7]) ? node2252 : node2245;
										assign node2245 = (inp[11]) ? 12'b000000111111 : node2246;
											assign node2246 = (inp[0]) ? node2248 : 12'b000001111111;
												assign node2248 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node2252 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node2255 = (inp[2]) ? node2267 : node2256;
									assign node2256 = (inp[0]) ? node2262 : node2257;
										assign node2257 = (inp[6]) ? 12'b000000111111 : node2258;
											assign node2258 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node2262 = (inp[7]) ? node2264 : 12'b000000111111;
											assign node2264 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
									assign node2267 = (inp[0]) ? node2277 : node2268;
										assign node2268 = (inp[7]) ? node2272 : node2269;
											assign node2269 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
											assign node2272 = (inp[11]) ? 12'b000000011111 : node2273;
												assign node2273 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
										assign node2277 = (inp[11]) ? node2279 : 12'b000000011111;
											assign node2279 = (inp[6]) ? 12'b000000001111 : node2280;
												assign node2280 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
						assign node2284 = (inp[0]) ? node2328 : node2285;
							assign node2285 = (inp[6]) ? node2303 : node2286;
								assign node2286 = (inp[2]) ? node2300 : node2287;
									assign node2287 = (inp[7]) ? node2295 : node2288;
										assign node2288 = (inp[11]) ? node2290 : 12'b000011111111;
											assign node2290 = (inp[5]) ? 12'b000001111111 : node2291;
												assign node2291 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node2295 = (inp[5]) ? node2297 : 12'b000001111111;
											assign node2297 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node2300 = (inp[4]) ? 12'b000000111111 : 12'b000011111111;
								assign node2303 = (inp[4]) ? node2311 : node2304;
									assign node2304 = (inp[11]) ? node2306 : 12'b000001111111;
										assign node2306 = (inp[2]) ? node2308 : 12'b000000111111;
											assign node2308 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node2311 = (inp[11]) ? node2319 : node2312;
										assign node2312 = (inp[2]) ? 12'b000000011111 : node2313;
											assign node2313 = (inp[7]) ? 12'b000000011111 : node2314;
												assign node2314 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node2319 = (inp[7]) ? node2323 : node2320;
											assign node2320 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
											assign node2323 = (inp[2]) ? node2325 : 12'b000000001111;
												assign node2325 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
							assign node2328 = (inp[5]) ? node2350 : node2329;
								assign node2329 = (inp[7]) ? node2339 : node2330;
									assign node2330 = (inp[11]) ? node2332 : 12'b000000111111;
										assign node2332 = (inp[6]) ? 12'b000000011111 : node2333;
											assign node2333 = (inp[4]) ? node2335 : 12'b000000111111;
												assign node2335 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
									assign node2339 = (inp[11]) ? node2345 : node2340;
										assign node2340 = (inp[2]) ? 12'b000000011111 : node2341;
											assign node2341 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
										assign node2345 = (inp[4]) ? node2347 : 12'b000000011111;
											assign node2347 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
								assign node2350 = (inp[7]) ? node2362 : node2351;
									assign node2351 = (inp[2]) ? node2357 : node2352;
										assign node2352 = (inp[6]) ? 12'b000000011111 : node2353;
											assign node2353 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node2357 = (inp[6]) ? node2359 : 12'b000000011111;
											assign node2359 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node2362 = (inp[6]) ? node2366 : node2363;
										assign node2363 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
										assign node2366 = (inp[4]) ? 12'b000000000011 : node2367;
											assign node2367 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
					assign node2371 = (inp[7]) ? node2491 : node2372;
						assign node2372 = (inp[1]) ? node2444 : node2373;
							assign node2373 = (inp[4]) ? node2403 : node2374;
								assign node2374 = (inp[2]) ? node2390 : node2375;
									assign node2375 = (inp[6]) ? node2377 : 12'b000001111111;
										assign node2377 = (inp[11]) ? node2385 : node2378;
											assign node2378 = (inp[0]) ? node2382 : node2379;
												assign node2379 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
												assign node2382 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
											assign node2385 = (inp[0]) ? 12'b000000111111 : node2386;
												assign node2386 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
									assign node2390 = (inp[6]) ? node2396 : node2391;
										assign node2391 = (inp[0]) ? 12'b000000111111 : node2392;
											assign node2392 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node2396 = (inp[5]) ? node2398 : 12'b000000111111;
											assign node2398 = (inp[0]) ? 12'b000000011111 : node2399;
												assign node2399 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node2403 = (inp[0]) ? node2427 : node2404;
									assign node2404 = (inp[11]) ? node2416 : node2405;
										assign node2405 = (inp[5]) ? node2411 : node2406;
											assign node2406 = (inp[6]) ? node2408 : 12'b000001111111;
												assign node2408 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
											assign node2411 = (inp[6]) ? node2413 : 12'b000000111111;
												assign node2413 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
										assign node2416 = (inp[6]) ? node2422 : node2417;
											assign node2417 = (inp[2]) ? node2419 : 12'b000000111111;
												assign node2419 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
											assign node2422 = (inp[5]) ? 12'b000000011111 : node2423;
												assign node2423 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
									assign node2427 = (inp[6]) ? node2439 : node2428;
										assign node2428 = (inp[2]) ? node2434 : node2429;
											assign node2429 = (inp[5]) ? node2431 : 12'b000000111111;
												assign node2431 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
											assign node2434 = (inp[5]) ? node2436 : 12'b000000011111;
												assign node2436 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node2439 = (inp[11]) ? 12'b000000001111 : node2440;
											assign node2440 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
							assign node2444 = (inp[4]) ? node2468 : node2445;
								assign node2445 = (inp[6]) ? node2453 : node2446;
									assign node2446 = (inp[0]) ? 12'b000000111111 : node2447;
										assign node2447 = (inp[11]) ? 12'b000000111111 : node2448;
											assign node2448 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
									assign node2453 = (inp[11]) ? node2459 : node2454;
										assign node2454 = (inp[5]) ? 12'b000000011111 : node2455;
											assign node2455 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node2459 = (inp[2]) ? node2463 : node2460;
											assign node2460 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
											assign node2463 = (inp[5]) ? node2465 : 12'b000000001111;
												assign node2465 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
								assign node2468 = (inp[2]) ? node2484 : node2469;
									assign node2469 = (inp[11]) ? node2473 : node2470;
										assign node2470 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
										assign node2473 = (inp[5]) ? node2479 : node2474;
											assign node2474 = (inp[0]) ? node2476 : 12'b000000011111;
												assign node2476 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
											assign node2479 = (inp[6]) ? 12'b000000001111 : node2480;
												assign node2480 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node2484 = (inp[0]) ? node2488 : node2485;
										assign node2485 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node2488 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
						assign node2491 = (inp[0]) ? node2545 : node2492;
							assign node2492 = (inp[5]) ? node2518 : node2493;
								assign node2493 = (inp[4]) ? node2503 : node2494;
									assign node2494 = (inp[2]) ? node2496 : 12'b000001111111;
										assign node2496 = (inp[1]) ? 12'b000000011111 : node2497;
											assign node2497 = (inp[11]) ? node2499 : 12'b000000111111;
												assign node2499 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
									assign node2503 = (inp[6]) ? node2513 : node2504;
										assign node2504 = (inp[1]) ? node2510 : node2505;
											assign node2505 = (inp[2]) ? node2507 : 12'b000000111111;
												assign node2507 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
											assign node2510 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
										assign node2513 = (inp[11]) ? node2515 : 12'b000000011111;
											assign node2515 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
								assign node2518 = (inp[11]) ? node2534 : node2519;
									assign node2519 = (inp[6]) ? node2525 : node2520;
										assign node2520 = (inp[1]) ? 12'b000000011111 : node2521;
											assign node2521 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
										assign node2525 = (inp[1]) ? 12'b000000001111 : node2526;
											assign node2526 = (inp[2]) ? node2530 : node2527;
												assign node2527 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
												assign node2530 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
									assign node2534 = (inp[6]) ? node2542 : node2535;
										assign node2535 = (inp[2]) ? node2537 : 12'b000000011111;
											assign node2537 = (inp[1]) ? 12'b000000001111 : node2538;
												assign node2538 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node2542 = (inp[1]) ? 12'b000000001111 : 12'b000000000111;
							assign node2545 = (inp[6]) ? node2577 : node2546;
								assign node2546 = (inp[5]) ? node2560 : node2547;
									assign node2547 = (inp[2]) ? node2555 : node2548;
										assign node2548 = (inp[11]) ? node2550 : 12'b000000111111;
											assign node2550 = (inp[1]) ? 12'b000000011111 : node2551;
												assign node2551 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
										assign node2555 = (inp[1]) ? node2557 : 12'b000000011111;
											assign node2557 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node2560 = (inp[4]) ? node2568 : node2561;
										assign node2561 = (inp[1]) ? node2565 : node2562;
											assign node2562 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
											assign node2565 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node2568 = (inp[2]) ? node2574 : node2569;
											assign node2569 = (inp[11]) ? node2571 : 12'b000000001111;
												assign node2571 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
											assign node2574 = (inp[1]) ? 12'b000000000011 : 12'b000000000111;
								assign node2577 = (inp[1]) ? node2593 : node2578;
									assign node2578 = (inp[2]) ? node2582 : node2579;
										assign node2579 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node2582 = (inp[5]) ? node2588 : node2583;
											assign node2583 = (inp[11]) ? 12'b000000001111 : node2584;
												assign node2584 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
											assign node2588 = (inp[11]) ? 12'b000000000111 : node2589;
												assign node2589 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
									assign node2593 = (inp[2]) ? node2599 : node2594;
										assign node2594 = (inp[11]) ? 12'b000000000111 : node2595;
											assign node2595 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
										assign node2599 = (inp[4]) ? 12'b000000000001 : 12'b000000000111;
			assign node2602 = (inp[6]) ? node3002 : node2603;
				assign node2603 = (inp[10]) ? node2785 : node2604;
					assign node2604 = (inp[5]) ? node2702 : node2605;
						assign node2605 = (inp[1]) ? node2655 : node2606;
							assign node2606 = (inp[0]) ? node2632 : node2607;
								assign node2607 = (inp[11]) ? node2625 : node2608;
									assign node2608 = (inp[2]) ? node2616 : node2609;
										assign node2609 = (inp[4]) ? 12'b000011111111 : node2610;
											assign node2610 = (inp[7]) ? 12'b000111111111 : node2611;
												assign node2611 = (inp[9]) ? 12'b000111111111 : 12'b001111111111;
										assign node2616 = (inp[9]) ? node2620 : node2617;
											assign node2617 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
											assign node2620 = (inp[7]) ? 12'b000001111111 : node2621;
												assign node2621 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node2625 = (inp[9]) ? 12'b000000111111 : node2626;
										assign node2626 = (inp[2]) ? node2628 : 12'b000011111111;
											assign node2628 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
								assign node2632 = (inp[9]) ? node2646 : node2633;
									assign node2633 = (inp[7]) ? node2643 : node2634;
										assign node2634 = (inp[4]) ? node2636 : 12'b000011111111;
											assign node2636 = (inp[2]) ? node2640 : node2637;
												assign node2637 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
												assign node2640 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node2643 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
									assign node2646 = (inp[4]) ? node2650 : node2647;
										assign node2647 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node2650 = (inp[7]) ? node2652 : 12'b000000111111;
											assign node2652 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
							assign node2655 = (inp[4]) ? node2681 : node2656;
								assign node2656 = (inp[9]) ? node2672 : node2657;
									assign node2657 = (inp[0]) ? node2665 : node2658;
										assign node2658 = (inp[2]) ? 12'b000001111111 : node2659;
											assign node2659 = (inp[11]) ? node2661 : 12'b000111111111;
												assign node2661 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
										assign node2665 = (inp[2]) ? 12'b000000111111 : node2666;
											assign node2666 = (inp[11]) ? node2668 : 12'b000011111111;
												assign node2668 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
									assign node2672 = (inp[11]) ? node2676 : node2673;
										assign node2673 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node2676 = (inp[7]) ? node2678 : 12'b000000111111;
											assign node2678 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
								assign node2681 = (inp[2]) ? node2691 : node2682;
									assign node2682 = (inp[9]) ? node2686 : node2683;
										assign node2683 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
										assign node2686 = (inp[0]) ? node2688 : 12'b000000111111;
											assign node2688 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node2691 = (inp[7]) ? node2699 : node2692;
										assign node2692 = (inp[9]) ? 12'b000000011111 : node2693;
											assign node2693 = (inp[11]) ? node2695 : 12'b000000111111;
												assign node2695 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node2699 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
						assign node2702 = (inp[11]) ? node2740 : node2703;
							assign node2703 = (inp[2]) ? node2729 : node2704;
								assign node2704 = (inp[1]) ? node2716 : node2705;
									assign node2705 = (inp[9]) ? node2713 : node2706;
										assign node2706 = (inp[4]) ? 12'b000001111111 : node2707;
											assign node2707 = (inp[0]) ? node2709 : 12'b000011111111;
												assign node2709 = (inp[7]) ? 12'b000001111111 : 12'b000011111111;
										assign node2713 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
									assign node2716 = (inp[0]) ? node2722 : node2717;
										assign node2717 = (inp[4]) ? 12'b000000111111 : node2718;
											assign node2718 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node2722 = (inp[7]) ? node2724 : 12'b000000111111;
											assign node2724 = (inp[9]) ? 12'b000000011111 : node2725;
												assign node2725 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
								assign node2729 = (inp[4]) ? node2735 : node2730;
									assign node2730 = (inp[7]) ? node2732 : 12'b000000111111;
										assign node2732 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node2735 = (inp[1]) ? 12'b000000001111 : node2736;
										assign node2736 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
							assign node2740 = (inp[1]) ? node2760 : node2741;
								assign node2741 = (inp[7]) ? node2753 : node2742;
									assign node2742 = (inp[9]) ? node2750 : node2743;
										assign node2743 = (inp[4]) ? 12'b000000111111 : node2744;
											assign node2744 = (inp[0]) ? node2746 : 12'b000001111111;
												assign node2746 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
										assign node2750 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node2753 = (inp[2]) ? node2757 : node2754;
										assign node2754 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
										assign node2757 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
								assign node2760 = (inp[4]) ? node2774 : node2761;
									assign node2761 = (inp[2]) ? node2769 : node2762;
										assign node2762 = (inp[0]) ? 12'b000000011111 : node2763;
											assign node2763 = (inp[9]) ? node2765 : 12'b000000111111;
												assign node2765 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
										assign node2769 = (inp[9]) ? node2771 : 12'b000000011111;
											assign node2771 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
									assign node2774 = (inp[9]) ? node2780 : node2775;
										assign node2775 = (inp[2]) ? 12'b000000001111 : node2776;
											assign node2776 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node2780 = (inp[0]) ? node2782 : 12'b000000001111;
											assign node2782 = (inp[2]) ? 12'b000000000011 : 12'b000000000111;
					assign node2785 = (inp[1]) ? node2909 : node2786;
						assign node2786 = (inp[0]) ? node2840 : node2787;
							assign node2787 = (inp[11]) ? node2823 : node2788;
								assign node2788 = (inp[5]) ? node2810 : node2789;
									assign node2789 = (inp[7]) ? node2797 : node2790;
										assign node2790 = (inp[2]) ? 12'b000001111111 : node2791;
											assign node2791 = (inp[9]) ? 12'b000011111111 : node2792;
												assign node2792 = (inp[4]) ? 12'b000011111111 : 12'b000111111111;
										assign node2797 = (inp[9]) ? node2805 : node2798;
											assign node2798 = (inp[4]) ? node2802 : node2799;
												assign node2799 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
												assign node2802 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
											assign node2805 = (inp[2]) ? node2807 : 12'b000000111111;
												assign node2807 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
									assign node2810 = (inp[9]) ? node2818 : node2811;
										assign node2811 = (inp[7]) ? 12'b000000111111 : node2812;
											assign node2812 = (inp[2]) ? node2814 : 12'b000001111111;
												assign node2814 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node2818 = (inp[7]) ? node2820 : 12'b000000111111;
											assign node2820 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
								assign node2823 = (inp[7]) ? node2833 : node2824;
									assign node2824 = (inp[2]) ? node2828 : node2825;
										assign node2825 = (inp[5]) ? 12'b000000111111 : 12'b000011111111;
										assign node2828 = (inp[5]) ? 12'b000000011111 : node2829;
											assign node2829 = (inp[9]) ? 12'b000000011111 : 12'b000001111111;
									assign node2833 = (inp[5]) ? node2837 : node2834;
										assign node2834 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
										assign node2837 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
							assign node2840 = (inp[9]) ? node2872 : node2841;
								assign node2841 = (inp[7]) ? node2853 : node2842;
									assign node2842 = (inp[2]) ? node2848 : node2843;
										assign node2843 = (inp[4]) ? 12'b000000111111 : node2844;
											assign node2844 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node2848 = (inp[5]) ? node2850 : 12'b000000111111;
											assign node2850 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
									assign node2853 = (inp[2]) ? node2861 : node2854;
										assign node2854 = (inp[4]) ? 12'b000000011111 : node2855;
											assign node2855 = (inp[11]) ? node2857 : 12'b000000111111;
												assign node2857 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node2861 = (inp[5]) ? node2867 : node2862;
											assign node2862 = (inp[4]) ? 12'b000000011111 : node2863;
												assign node2863 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
											assign node2867 = (inp[11]) ? 12'b000000001111 : node2868;
												assign node2868 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node2872 = (inp[2]) ? node2894 : node2873;
									assign node2873 = (inp[4]) ? node2881 : node2874;
										assign node2874 = (inp[11]) ? 12'b000000011111 : node2875;
											assign node2875 = (inp[7]) ? 12'b000000111111 : node2876;
												assign node2876 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node2881 = (inp[11]) ? node2889 : node2882;
											assign node2882 = (inp[5]) ? node2886 : node2883;
												assign node2883 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
												assign node2886 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
											assign node2889 = (inp[7]) ? 12'b000000001111 : node2890;
												assign node2890 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
									assign node2894 = (inp[4]) ? node2906 : node2895;
										assign node2895 = (inp[11]) ? node2901 : node2896;
											assign node2896 = (inp[5]) ? node2898 : 12'b000000011111;
												assign node2898 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
											assign node2901 = (inp[5]) ? 12'b000000001111 : node2902;
												assign node2902 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node2906 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
						assign node2909 = (inp[0]) ? node2951 : node2910;
							assign node2910 = (inp[7]) ? node2926 : node2911;
								assign node2911 = (inp[2]) ? node2921 : node2912;
									assign node2912 = (inp[4]) ? node2918 : node2913;
										assign node2913 = (inp[5]) ? node2915 : 12'b000001111111;
											assign node2915 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node2918 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node2921 = (inp[11]) ? 12'b000000011111 : node2922;
										assign node2922 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
								assign node2926 = (inp[9]) ? node2940 : node2927;
									assign node2927 = (inp[5]) ? node2929 : 12'b000000111111;
										assign node2929 = (inp[11]) ? node2935 : node2930;
											assign node2930 = (inp[4]) ? 12'b000000011111 : node2931;
												assign node2931 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
											assign node2935 = (inp[2]) ? 12'b000000001111 : node2936;
												assign node2936 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
									assign node2940 = (inp[5]) ? node2944 : node2941;
										assign node2941 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
										assign node2944 = (inp[11]) ? node2946 : 12'b000000001111;
											assign node2946 = (inp[2]) ? 12'b000000000111 : node2947;
												assign node2947 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
							assign node2951 = (inp[9]) ? node2975 : node2952;
								assign node2952 = (inp[5]) ? node2968 : node2953;
									assign node2953 = (inp[2]) ? node2961 : node2954;
										assign node2954 = (inp[7]) ? node2956 : 12'b000000011111;
											assign node2956 = (inp[4]) ? node2958 : 12'b000000011111;
												assign node2958 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node2961 = (inp[11]) ? 12'b000000001111 : node2962;
											assign node2962 = (inp[4]) ? node2964 : 12'b000000011111;
												assign node2964 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
									assign node2968 = (inp[2]) ? node2972 : node2969;
										assign node2969 = (inp[4]) ? 12'b000000001111 : 12'b000000111111;
										assign node2972 = (inp[11]) ? 12'b000000000011 : 12'b000000001111;
								assign node2975 = (inp[4]) ? node2987 : node2976;
									assign node2976 = (inp[5]) ? node2984 : node2977;
										assign node2977 = (inp[2]) ? node2979 : 12'b000000111111;
											assign node2979 = (inp[11]) ? 12'b000000001111 : node2980;
												assign node2980 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node2984 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
									assign node2987 = (inp[2]) ? node2995 : node2988;
										assign node2988 = (inp[11]) ? 12'b000000000111 : node2989;
											assign node2989 = (inp[5]) ? node2991 : 12'b000000001111;
												assign node2991 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
										assign node2995 = (inp[5]) ? node2997 : 12'b000000000111;
											assign node2997 = (inp[7]) ? 12'b000000000011 : node2998;
												assign node2998 = (inp[11]) ? 12'b000000000011 : 12'b000000000111;
				assign node3002 = (inp[4]) ? node3198 : node3003;
					assign node3003 = (inp[2]) ? node3107 : node3004;
						assign node3004 = (inp[0]) ? node3048 : node3005;
							assign node3005 = (inp[1]) ? node3019 : node3006;
								assign node3006 = (inp[11]) ? node3010 : node3007;
									assign node3007 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
									assign node3010 = (inp[9]) ? node3016 : node3011;
										assign node3011 = (inp[10]) ? node3013 : 12'b000001111111;
											assign node3013 = (inp[7]) ? 12'b000000011111 : 12'b000001111111;
										assign node3016 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
								assign node3019 = (inp[7]) ? node3037 : node3020;
									assign node3020 = (inp[11]) ? node3030 : node3021;
										assign node3021 = (inp[10]) ? node3023 : 12'b000001111111;
											assign node3023 = (inp[9]) ? node3027 : node3024;
												assign node3024 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
												assign node3027 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node3030 = (inp[10]) ? node3032 : 12'b000000111111;
											assign node3032 = (inp[5]) ? 12'b000000011111 : node3033;
												assign node3033 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node3037 = (inp[9]) ? node3045 : node3038;
										assign node3038 = (inp[10]) ? 12'b000000011111 : node3039;
											assign node3039 = (inp[11]) ? node3041 : 12'b000000111111;
												assign node3041 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node3045 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
							assign node3048 = (inp[5]) ? node3076 : node3049;
								assign node3049 = (inp[9]) ? node3065 : node3050;
									assign node3050 = (inp[11]) ? node3058 : node3051;
										assign node3051 = (inp[10]) ? 12'b000000111111 : node3052;
											assign node3052 = (inp[7]) ? node3054 : 12'b000001111111;
												assign node3054 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node3058 = (inp[1]) ? node3060 : 12'b000000111111;
											assign node3060 = (inp[10]) ? 12'b000000011111 : node3061;
												assign node3061 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
									assign node3065 = (inp[1]) ? 12'b000000001111 : node3066;
										assign node3066 = (inp[11]) ? node3068 : 12'b000000111111;
											assign node3068 = (inp[7]) ? node3072 : node3069;
												assign node3069 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
												assign node3072 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
								assign node3076 = (inp[1]) ? node3094 : node3077;
									assign node3077 = (inp[7]) ? node3085 : node3078;
										assign node3078 = (inp[9]) ? 12'b000000011111 : node3079;
											assign node3079 = (inp[10]) ? node3081 : 12'b000000111111;
												assign node3081 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node3085 = (inp[9]) ? 12'b000000001111 : node3086;
											assign node3086 = (inp[10]) ? node3090 : node3087;
												assign node3087 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
												assign node3090 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node3094 = (inp[9]) ? node3100 : node3095;
										assign node3095 = (inp[11]) ? 12'b000000001111 : node3096;
											assign node3096 = (inp[7]) ? 12'b000000001111 : 12'b000000011111;
										assign node3100 = (inp[10]) ? 12'b000000000111 : node3101;
											assign node3101 = (inp[7]) ? node3103 : 12'b000000001111;
												assign node3103 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
						assign node3107 = (inp[11]) ? node3151 : node3108;
							assign node3108 = (inp[1]) ? node3136 : node3109;
								assign node3109 = (inp[9]) ? node3125 : node3110;
									assign node3110 = (inp[0]) ? node3118 : node3111;
										assign node3111 = (inp[10]) ? node3113 : 12'b000001111111;
											assign node3113 = (inp[5]) ? 12'b000000111111 : node3114;
												assign node3114 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
										assign node3118 = (inp[10]) ? 12'b000000011111 : node3119;
											assign node3119 = (inp[7]) ? node3121 : 12'b000000111111;
												assign node3121 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node3125 = (inp[5]) ? node3131 : node3126;
										assign node3126 = (inp[7]) ? 12'b000000011111 : node3127;
											assign node3127 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node3131 = (inp[10]) ? 12'b000000001111 : node3132;
											assign node3132 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
								assign node3136 = (inp[7]) ? node3144 : node3137;
									assign node3137 = (inp[9]) ? node3139 : 12'b000000011111;
										assign node3139 = (inp[0]) ? 12'b000000011111 : node3140;
											assign node3140 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node3144 = (inp[5]) ? node3146 : 12'b000000001111;
										assign node3146 = (inp[10]) ? node3148 : 12'b000000001111;
											assign node3148 = (inp[9]) ? 12'b000000000011 : 12'b000000000111;
							assign node3151 = (inp[1]) ? node3181 : node3152;
								assign node3152 = (inp[5]) ? node3158 : node3153;
									assign node3153 = (inp[10]) ? node3155 : 12'b000000011111;
										assign node3155 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
									assign node3158 = (inp[7]) ? node3170 : node3159;
										assign node3159 = (inp[9]) ? node3165 : node3160;
											assign node3160 = (inp[10]) ? node3162 : 12'b000000011111;
												assign node3162 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
											assign node3165 = (inp[10]) ? 12'b000000001111 : node3166;
												assign node3166 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
										assign node3170 = (inp[0]) ? node3176 : node3171;
											assign node3171 = (inp[9]) ? node3173 : 12'b000000001111;
												assign node3173 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
											assign node3176 = (inp[9]) ? 12'b000000000111 : node3177;
												assign node3177 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
								assign node3181 = (inp[5]) ? node3187 : node3182;
									assign node3182 = (inp[0]) ? node3184 : 12'b000000001111;
										assign node3184 = (inp[9]) ? 12'b000000000011 : 12'b000000001111;
									assign node3187 = (inp[10]) ? node3191 : node3188;
										assign node3188 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
										assign node3191 = (inp[7]) ? node3193 : 12'b000000000111;
											assign node3193 = (inp[9]) ? 12'b000000000011 : node3194;
												assign node3194 = (inp[0]) ? 12'b000000000011 : 12'b000000000111;
					assign node3198 = (inp[7]) ? node3316 : node3199;
						assign node3199 = (inp[5]) ? node3261 : node3200;
							assign node3200 = (inp[2]) ? node3232 : node3201;
								assign node3201 = (inp[10]) ? node3215 : node3202;
									assign node3202 = (inp[9]) ? node3204 : 12'b000001111111;
										assign node3204 = (inp[1]) ? node3210 : node3205;
											assign node3205 = (inp[11]) ? 12'b000000111111 : node3206;
												assign node3206 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
											assign node3210 = (inp[0]) ? 12'b000000011111 : node3211;
												assign node3211 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node3215 = (inp[1]) ? node3227 : node3216;
										assign node3216 = (inp[0]) ? node3222 : node3217;
											assign node3217 = (inp[11]) ? 12'b000000111111 : node3218;
												assign node3218 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
											assign node3222 = (inp[9]) ? node3224 : 12'b000000011111;
												assign node3224 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
										assign node3227 = (inp[9]) ? node3229 : 12'b000000011111;
											assign node3229 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
								assign node3232 = (inp[11]) ? node3248 : node3233;
									assign node3233 = (inp[0]) ? node3241 : node3234;
										assign node3234 = (inp[10]) ? node3236 : 12'b000000111111;
											assign node3236 = (inp[9]) ? 12'b000000011111 : node3237;
												assign node3237 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
										assign node3241 = (inp[10]) ? 12'b000000001111 : node3242;
											assign node3242 = (inp[1]) ? 12'b000000001111 : node3243;
												assign node3243 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node3248 = (inp[0]) ? node3258 : node3249;
										assign node3249 = (inp[1]) ? node3251 : 12'b000000011111;
											assign node3251 = (inp[9]) ? node3255 : node3252;
												assign node3252 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
												assign node3255 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
										assign node3258 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
							assign node3261 = (inp[0]) ? node3283 : node3262;
								assign node3262 = (inp[10]) ? node3276 : node3263;
									assign node3263 = (inp[11]) ? node3271 : node3264;
										assign node3264 = (inp[9]) ? node3266 : 12'b000000111111;
											assign node3266 = (inp[2]) ? node3268 : 12'b000000011111;
												assign node3268 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
										assign node3271 = (inp[9]) ? 12'b000000001111 : node3272;
											assign node3272 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
									assign node3276 = (inp[1]) ? node3280 : node3277;
										assign node3277 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
										assign node3280 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
								assign node3283 = (inp[2]) ? node3297 : node3284;
									assign node3284 = (inp[11]) ? node3290 : node3285;
										assign node3285 = (inp[1]) ? 12'b000000001111 : node3286;
											assign node3286 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
										assign node3290 = (inp[10]) ? 12'b000000000111 : node3291;
											assign node3291 = (inp[9]) ? node3293 : 12'b000000001111;
												assign node3293 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
									assign node3297 = (inp[1]) ? node3311 : node3298;
										assign node3298 = (inp[11]) ? node3304 : node3299;
											assign node3299 = (inp[10]) ? node3301 : 12'b000000001111;
												assign node3301 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
											assign node3304 = (inp[9]) ? node3308 : node3305;
												assign node3305 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
												assign node3308 = (inp[10]) ? 12'b000000000011 : 12'b000000000111;
										assign node3311 = (inp[9]) ? node3313 : 12'b000000000111;
											assign node3313 = (inp[11]) ? 12'b000000000001 : 12'b000000000111;
						assign node3316 = (inp[11]) ? node3370 : node3317;
							assign node3317 = (inp[5]) ? node3343 : node3318;
								assign node3318 = (inp[9]) ? node3330 : node3319;
									assign node3319 = (inp[1]) ? node3323 : node3320;
										assign node3320 = (inp[10]) ? 12'b000000011111 : 12'b000001111111;
										assign node3323 = (inp[10]) ? 12'b000000001111 : node3324;
											assign node3324 = (inp[2]) ? node3326 : 12'b000000011111;
												assign node3326 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node3330 = (inp[10]) ? node3336 : node3331;
										assign node3331 = (inp[0]) ? 12'b000000001111 : node3332;
											assign node3332 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
										assign node3336 = (inp[2]) ? node3338 : 12'b000000001111;
											assign node3338 = (inp[0]) ? 12'b000000000111 : node3339;
												assign node3339 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
								assign node3343 = (inp[1]) ? node3357 : node3344;
									assign node3344 = (inp[0]) ? node3352 : node3345;
										assign node3345 = (inp[9]) ? 12'b000000001111 : node3346;
											assign node3346 = (inp[2]) ? node3348 : 12'b000000011111;
												assign node3348 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
										assign node3352 = (inp[2]) ? 12'b000000000111 : node3353;
											assign node3353 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
									assign node3357 = (inp[10]) ? node3365 : node3358;
										assign node3358 = (inp[0]) ? node3360 : 12'b000000001111;
											assign node3360 = (inp[9]) ? 12'b000000000111 : node3361;
												assign node3361 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
										assign node3365 = (inp[2]) ? node3367 : 12'b000000000111;
											assign node3367 = (inp[9]) ? 12'b000000000011 : 12'b000000000111;
							assign node3370 = (inp[5]) ? node3406 : node3371;
								assign node3371 = (inp[2]) ? node3387 : node3372;
									assign node3372 = (inp[1]) ? node3378 : node3373;
										assign node3373 = (inp[0]) ? 12'b000000001111 : node3374;
											assign node3374 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
										assign node3378 = (inp[0]) ? node3384 : node3379;
											assign node3379 = (inp[10]) ? node3381 : 12'b000000001111;
												assign node3381 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
											assign node3384 = (inp[9]) ? 12'b000000000011 : 12'b000000000111;
									assign node3387 = (inp[9]) ? node3395 : node3388;
										assign node3388 = (inp[0]) ? 12'b000000000111 : node3389;
											assign node3389 = (inp[10]) ? node3391 : 12'b000000001111;
												assign node3391 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
										assign node3395 = (inp[10]) ? node3401 : node3396;
											assign node3396 = (inp[0]) ? node3398 : 12'b000000000111;
												assign node3398 = (inp[1]) ? 12'b000000000011 : 12'b000000000111;
											assign node3401 = (inp[1]) ? 12'b000000000011 : node3402;
												assign node3402 = (inp[0]) ? 12'b000000000011 : 12'b000000000111;
								assign node3406 = (inp[1]) ? node3422 : node3407;
									assign node3407 = (inp[10]) ? node3415 : node3408;
										assign node3408 = (inp[2]) ? node3410 : 12'b000000001111;
											assign node3410 = (inp[9]) ? 12'b000000000111 : node3411;
												assign node3411 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
										assign node3415 = (inp[2]) ? node3417 : 12'b000000000111;
											assign node3417 = (inp[0]) ? node3419 : 12'b000000000011;
												assign node3419 = (inp[9]) ? 12'b000000000001 : 12'b000000000011;
									assign node3422 = (inp[9]) ? node3424 : 12'b000000000011;
										assign node3424 = (inp[0]) ? 12'b000000000001 : node3425;
											assign node3425 = (inp[10]) ? node3427 : 12'b000000000011;
												assign node3427 = (inp[2]) ? 12'b000000000001 : 12'b000000000011;

endmodule