module dtc_split33_bm22 (
	input  wire [11-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node12;
	wire [11-1:0] node13;
	wire [11-1:0] node17;
	wire [11-1:0] node18;
	wire [11-1:0] node20;
	wire [11-1:0] node23;
	wire [11-1:0] node24;
	wire [11-1:0] node27;
	wire [11-1:0] node30;
	wire [11-1:0] node31;
	wire [11-1:0] node32;
	wire [11-1:0] node35;
	wire [11-1:0] node36;
	wire [11-1:0] node40;
	wire [11-1:0] node41;
	wire [11-1:0] node42;
	wire [11-1:0] node45;
	wire [11-1:0] node48;
	wire [11-1:0] node49;
	wire [11-1:0] node53;
	wire [11-1:0] node54;
	wire [11-1:0] node55;
	wire [11-1:0] node56;
	wire [11-1:0] node57;
	wire [11-1:0] node60;
	wire [11-1:0] node63;
	wire [11-1:0] node64;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node70;
	wire [11-1:0] node73;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node83;
	wire [11-1:0] node86;
	wire [11-1:0] node87;
	wire [11-1:0] node91;
	wire [11-1:0] node92;
	wire [11-1:0] node93;
	wire [11-1:0] node96;
	wire [11-1:0] node99;
	wire [11-1:0] node101;
	wire [11-1:0] node104;
	wire [11-1:0] node105;
	wire [11-1:0] node106;
	wire [11-1:0] node107;
	wire [11-1:0] node108;
	wire [11-1:0] node109;
	wire [11-1:0] node113;
	wire [11-1:0] node114;
	wire [11-1:0] node118;
	wire [11-1:0] node119;
	wire [11-1:0] node120;
	wire [11-1:0] node124;
	wire [11-1:0] node125;
	wire [11-1:0] node128;
	wire [11-1:0] node131;
	wire [11-1:0] node132;
	wire [11-1:0] node133;
	wire [11-1:0] node134;
	wire [11-1:0] node137;
	wire [11-1:0] node140;
	wire [11-1:0] node141;
	wire [11-1:0] node145;
	wire [11-1:0] node146;
	wire [11-1:0] node149;
	wire [11-1:0] node150;
	wire [11-1:0] node153;
	wire [11-1:0] node156;
	wire [11-1:0] node157;
	wire [11-1:0] node158;
	wire [11-1:0] node159;
	wire [11-1:0] node160;
	wire [11-1:0] node164;
	wire [11-1:0] node165;
	wire [11-1:0] node169;
	wire [11-1:0] node170;
	wire [11-1:0] node171;
	wire [11-1:0] node174;
	wire [11-1:0] node177;
	wire [11-1:0] node178;
	wire [11-1:0] node182;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node185;
	wire [11-1:0] node188;
	wire [11-1:0] node191;
	wire [11-1:0] node192;
	wire [11-1:0] node195;
	wire [11-1:0] node198;
	wire [11-1:0] node199;
	wire [11-1:0] node203;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node206;
	wire [11-1:0] node207;
	wire [11-1:0] node208;
	wire [11-1:0] node209;
	wire [11-1:0] node212;
	wire [11-1:0] node215;
	wire [11-1:0] node216;
	wire [11-1:0] node219;
	wire [11-1:0] node222;
	wire [11-1:0] node223;
	wire [11-1:0] node225;
	wire [11-1:0] node228;
	wire [11-1:0] node229;
	wire [11-1:0] node233;
	wire [11-1:0] node234;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node241;
	wire [11-1:0] node242;
	wire [11-1:0] node244;
	wire [11-1:0] node247;
	wire [11-1:0] node248;
	wire [11-1:0] node252;
	wire [11-1:0] node253;
	wire [11-1:0] node254;
	wire [11-1:0] node255;
	wire [11-1:0] node256;
	wire [11-1:0] node259;
	wire [11-1:0] node262;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node269;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node274;
	wire [11-1:0] node277;
	wire [11-1:0] node278;
	wire [11-1:0] node281;
	wire [11-1:0] node284;
	wire [11-1:0] node285;
	wire [11-1:0] node286;
	wire [11-1:0] node287;
	wire [11-1:0] node290;
	wire [11-1:0] node293;
	wire [11-1:0] node294;
	wire [11-1:0] node298;
	wire [11-1:0] node299;
	wire [11-1:0] node301;
	wire [11-1:0] node304;
	wire [11-1:0] node305;
	wire [11-1:0] node308;
	wire [11-1:0] node311;
	wire [11-1:0] node312;
	wire [11-1:0] node313;
	wire [11-1:0] node314;
	wire [11-1:0] node316;
	wire [11-1:0] node317;
	wire [11-1:0] node321;
	wire [11-1:0] node323;
	wire [11-1:0] node326;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node336;
	wire [11-1:0] node337;
	wire [11-1:0] node339;
	wire [11-1:0] node342;
	wire [11-1:0] node343;
	wire [11-1:0] node346;
	wire [11-1:0] node349;
	wire [11-1:0] node350;
	wire [11-1:0] node351;
	wire [11-1:0] node352;
	wire [11-1:0] node353;
	wire [11-1:0] node356;
	wire [11-1:0] node359;
	wire [11-1:0] node360;
	wire [11-1:0] node364;
	wire [11-1:0] node365;
	wire [11-1:0] node366;
	wire [11-1:0] node369;
	wire [11-1:0] node372;
	wire [11-1:0] node373;
	wire [11-1:0] node376;
	wire [11-1:0] node379;
	wire [11-1:0] node380;
	wire [11-1:0] node381;
	wire [11-1:0] node384;
	wire [11-1:0] node385;
	wire [11-1:0] node389;
	wire [11-1:0] node390;
	wire [11-1:0] node393;
	wire [11-1:0] node394;
	wire [11-1:0] node397;
	wire [11-1:0] node400;
	wire [11-1:0] node401;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node404;
	wire [11-1:0] node405;
	wire [11-1:0] node406;
	wire [11-1:0] node407;
	wire [11-1:0] node411;
	wire [11-1:0] node413;
	wire [11-1:0] node416;
	wire [11-1:0] node417;
	wire [11-1:0] node418;
	wire [11-1:0] node421;
	wire [11-1:0] node424;
	wire [11-1:0] node425;
	wire [11-1:0] node428;
	wire [11-1:0] node431;
	wire [11-1:0] node432;
	wire [11-1:0] node433;
	wire [11-1:0] node435;
	wire [11-1:0] node438;
	wire [11-1:0] node439;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node445;
	wire [11-1:0] node448;
	wire [11-1:0] node451;
	wire [11-1:0] node454;
	wire [11-1:0] node455;
	wire [11-1:0] node456;
	wire [11-1:0] node457;
	wire [11-1:0] node459;
	wire [11-1:0] node462;
	wire [11-1:0] node463;
	wire [11-1:0] node466;
	wire [11-1:0] node469;
	wire [11-1:0] node470;
	wire [11-1:0] node471;
	wire [11-1:0] node474;
	wire [11-1:0] node477;
	wire [11-1:0] node479;
	wire [11-1:0] node482;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node485;
	wire [11-1:0] node488;
	wire [11-1:0] node491;
	wire [11-1:0] node494;
	wire [11-1:0] node495;
	wire [11-1:0] node496;
	wire [11-1:0] node499;
	wire [11-1:0] node502;
	wire [11-1:0] node503;
	wire [11-1:0] node506;
	wire [11-1:0] node509;
	wire [11-1:0] node510;
	wire [11-1:0] node511;
	wire [11-1:0] node512;
	wire [11-1:0] node513;
	wire [11-1:0] node516;
	wire [11-1:0] node517;
	wire [11-1:0] node520;
	wire [11-1:0] node523;
	wire [11-1:0] node524;
	wire [11-1:0] node527;
	wire [11-1:0] node528;
	wire [11-1:0] node532;
	wire [11-1:0] node533;
	wire [11-1:0] node534;
	wire [11-1:0] node535;
	wire [11-1:0] node538;
	wire [11-1:0] node541;
	wire [11-1:0] node542;
	wire [11-1:0] node545;
	wire [11-1:0] node548;
	wire [11-1:0] node549;
	wire [11-1:0] node553;
	wire [11-1:0] node554;
	wire [11-1:0] node555;
	wire [11-1:0] node556;
	wire [11-1:0] node557;
	wire [11-1:0] node561;
	wire [11-1:0] node562;
	wire [11-1:0] node565;
	wire [11-1:0] node568;
	wire [11-1:0] node569;
	wire [11-1:0] node571;
	wire [11-1:0] node575;
	wire [11-1:0] node576;
	wire [11-1:0] node577;
	wire [11-1:0] node580;
	wire [11-1:0] node582;
	wire [11-1:0] node585;
	wire [11-1:0] node586;
	wire [11-1:0] node587;
	wire [11-1:0] node590;
	wire [11-1:0] node593;
	wire [11-1:0] node594;
	wire [11-1:0] node597;
	wire [11-1:0] node600;
	wire [11-1:0] node601;
	wire [11-1:0] node602;
	wire [11-1:0] node603;
	wire [11-1:0] node604;
	wire [11-1:0] node605;
	wire [11-1:0] node606;
	wire [11-1:0] node609;
	wire [11-1:0] node612;
	wire [11-1:0] node615;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node620;
	wire [11-1:0] node624;
	wire [11-1:0] node625;
	wire [11-1:0] node626;
	wire [11-1:0] node627;
	wire [11-1:0] node630;
	wire [11-1:0] node634;
	wire [11-1:0] node635;
	wire [11-1:0] node636;
	wire [11-1:0] node639;
	wire [11-1:0] node642;
	wire [11-1:0] node644;
	wire [11-1:0] node647;
	wire [11-1:0] node648;
	wire [11-1:0] node649;
	wire [11-1:0] node650;
	wire [11-1:0] node651;
	wire [11-1:0] node655;
	wire [11-1:0] node656;
	wire [11-1:0] node660;
	wire [11-1:0] node661;
	wire [11-1:0] node662;
	wire [11-1:0] node665;
	wire [11-1:0] node668;
	wire [11-1:0] node670;
	wire [11-1:0] node673;
	wire [11-1:0] node674;
	wire [11-1:0] node676;
	wire [11-1:0] node677;
	wire [11-1:0] node680;
	wire [11-1:0] node683;
	wire [11-1:0] node684;
	wire [11-1:0] node685;
	wire [11-1:0] node688;
	wire [11-1:0] node691;
	wire [11-1:0] node692;
	wire [11-1:0] node695;
	wire [11-1:0] node698;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node701;
	wire [11-1:0] node702;
	wire [11-1:0] node704;
	wire [11-1:0] node707;
	wire [11-1:0] node710;
	wire [11-1:0] node711;
	wire [11-1:0] node714;
	wire [11-1:0] node715;
	wire [11-1:0] node718;
	wire [11-1:0] node721;
	wire [11-1:0] node722;
	wire [11-1:0] node723;
	wire [11-1:0] node724;
	wire [11-1:0] node727;
	wire [11-1:0] node730;
	wire [11-1:0] node731;
	wire [11-1:0] node734;
	wire [11-1:0] node737;
	wire [11-1:0] node738;
	wire [11-1:0] node740;
	wire [11-1:0] node743;
	wire [11-1:0] node744;
	wire [11-1:0] node747;
	wire [11-1:0] node750;
	wire [11-1:0] node751;
	wire [11-1:0] node752;
	wire [11-1:0] node753;
	wire [11-1:0] node755;
	wire [11-1:0] node758;
	wire [11-1:0] node759;
	wire [11-1:0] node762;
	wire [11-1:0] node765;
	wire [11-1:0] node766;
	wire [11-1:0] node767;
	wire [11-1:0] node770;
	wire [11-1:0] node773;
	wire [11-1:0] node774;
	wire [11-1:0] node777;
	wire [11-1:0] node780;
	wire [11-1:0] node781;
	wire [11-1:0] node782;
	wire [11-1:0] node783;
	wire [11-1:0] node786;
	wire [11-1:0] node789;
	wire [11-1:0] node790;
	wire [11-1:0] node793;
	wire [11-1:0] node796;
	wire [11-1:0] node797;
	wire [11-1:0] node798;
	wire [11-1:0] node801;
	wire [11-1:0] node804;
	wire [11-1:0] node805;
	wire [11-1:0] node808;

	assign outp = (inp[6]) ? node400 : node1;
		assign node1 = (inp[5]) ? node203 : node2;
			assign node2 = (inp[9]) ? node104 : node3;
				assign node3 = (inp[10]) ? node53 : node4;
					assign node4 = (inp[8]) ? node30 : node5;
						assign node5 = (inp[0]) ? node17 : node6;
							assign node6 = (inp[2]) ? node12 : node7;
								assign node7 = (inp[1]) ? 11'b00011111111 : node8;
									assign node8 = (inp[7]) ? 11'b00111111111 : 11'b01111111111;
								assign node12 = (inp[7]) ? 11'b00011111111 : node13;
									assign node13 = (inp[3]) ? 11'b00011111111 : 11'b00111111111;
							assign node17 = (inp[4]) ? node23 : node18;
								assign node18 = (inp[3]) ? node20 : 11'b00111111111;
									assign node20 = (inp[1]) ? 11'b00001111111 : 11'b00011111111;
								assign node23 = (inp[3]) ? node27 : node24;
									assign node24 = (inp[2]) ? 11'b00001111111 : 11'b00011111111;
									assign node27 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
						assign node30 = (inp[0]) ? node40 : node31;
							assign node31 = (inp[4]) ? node35 : node32;
								assign node32 = (inp[7]) ? 11'b00001111111 : 11'b00111111111;
								assign node35 = (inp[2]) ? 11'b00001111111 : node36;
									assign node36 = (inp[1]) ? 11'b00001111111 : 11'b00001111111;
							assign node40 = (inp[3]) ? node48 : node41;
								assign node41 = (inp[1]) ? node45 : node42;
									assign node42 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
									assign node45 = (inp[2]) ? 11'b00000111111 : 11'b00011111111;
								assign node48 = (inp[7]) ? 11'b00000111111 : node49;
									assign node49 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
					assign node53 = (inp[2]) ? node81 : node54;
						assign node54 = (inp[4]) ? node68 : node55;
							assign node55 = (inp[1]) ? node63 : node56;
								assign node56 = (inp[8]) ? node60 : node57;
									assign node57 = (inp[3]) ? 11'b00011111111 : 11'b00111111111;
									assign node60 = (inp[3]) ? 11'b00001111111 : 11'b00011111111;
								assign node63 = (inp[3]) ? 11'b00001111111 : node64;
									assign node64 = (inp[0]) ? 11'b00001111111 : 11'b00001111111;
							assign node68 = (inp[3]) ? node76 : node69;
								assign node69 = (inp[1]) ? node73 : node70;
									assign node70 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node73 = (inp[7]) ? 11'b00000111111 : 11'b00000111111;
								assign node76 = (inp[8]) ? 11'b00000111111 : node77;
									assign node77 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
						assign node81 = (inp[7]) ? node91 : node82;
							assign node82 = (inp[1]) ? node86 : node83;
								assign node83 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
								assign node86 = (inp[8]) ? 11'b00000111111 : node87;
									assign node87 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
							assign node91 = (inp[1]) ? node99 : node92;
								assign node92 = (inp[0]) ? node96 : node93;
									assign node93 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node96 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node99 = (inp[8]) ? node101 : 11'b00000111111;
									assign node101 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
				assign node104 = (inp[3]) ? node156 : node105;
					assign node105 = (inp[4]) ? node131 : node106;
						assign node106 = (inp[1]) ? node118 : node107;
							assign node107 = (inp[10]) ? node113 : node108;
								assign node108 = (inp[2]) ? 11'b00011111111 : node109;
									assign node109 = (inp[8]) ? 11'b00011111111 : 11'b00011111111;
								assign node113 = (inp[7]) ? 11'b00000111111 : node114;
									assign node114 = (inp[0]) ? 11'b00001111111 : 11'b00011111111;
							assign node118 = (inp[0]) ? node124 : node119;
								assign node119 = (inp[8]) ? 11'b00001111111 : node120;
									assign node120 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
								assign node124 = (inp[7]) ? node128 : node125;
									assign node125 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node128 = (inp[8]) ? 11'b00000111111 : 11'b00000111111;
						assign node131 = (inp[2]) ? node145 : node132;
							assign node132 = (inp[10]) ? node140 : node133;
								assign node133 = (inp[1]) ? node137 : node134;
									assign node134 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
									assign node137 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node140 = (inp[0]) ? 11'b00000111111 : node141;
									assign node141 = (inp[8]) ? 11'b00000111111 : 11'b00000111111;
							assign node145 = (inp[7]) ? node149 : node146;
								assign node146 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node149 = (inp[8]) ? node153 : node150;
									assign node150 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
									assign node153 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
					assign node156 = (inp[8]) ? node182 : node157;
						assign node157 = (inp[0]) ? node169 : node158;
							assign node158 = (inp[4]) ? node164 : node159;
								assign node159 = (inp[7]) ? 11'b00001111111 : node160;
									assign node160 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
								assign node164 = (inp[2]) ? 11'b00000111111 : node165;
									assign node165 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
							assign node169 = (inp[1]) ? node177 : node170;
								assign node170 = (inp[10]) ? node174 : node171;
									assign node171 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
									assign node174 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node177 = (inp[10]) ? 11'b00000001111 : node178;
									assign node178 = (inp[7]) ? 11'b00000011111 : 11'b00000011111;
						assign node182 = (inp[7]) ? node198 : node183;
							assign node183 = (inp[2]) ? node191 : node184;
								assign node184 = (inp[1]) ? node188 : node185;
									assign node185 = (inp[4]) ? 11'b00000111111 : 11'b00000111111;
									assign node188 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node191 = (inp[4]) ? node195 : node192;
									assign node192 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
									assign node195 = (inp[0]) ? 11'b00000000111 : 11'b00000011111;
							assign node198 = (inp[10]) ? 11'b00000001111 : node199;
								assign node199 = (inp[1]) ? 11'b00000000111 : 11'b00000001111;
			assign node203 = (inp[4]) ? node311 : node204;
				assign node204 = (inp[2]) ? node252 : node205;
					assign node205 = (inp[1]) ? node233 : node206;
						assign node206 = (inp[9]) ? node222 : node207;
							assign node207 = (inp[0]) ? node215 : node208;
								assign node208 = (inp[7]) ? node212 : node209;
									assign node209 = (inp[3]) ? 11'b00011111111 : 11'b00111111111;
									assign node212 = (inp[3]) ? 11'b00001111111 : 11'b00011111111;
								assign node215 = (inp[3]) ? node219 : node216;
									assign node216 = (inp[10]) ? 11'b00001111111 : 11'b00011111111;
									assign node219 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node222 = (inp[3]) ? node228 : node223;
								assign node223 = (inp[10]) ? node225 : 11'b00001111111;
									assign node225 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node228 = (inp[0]) ? 11'b00000111111 : node229;
									assign node229 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
						assign node233 = (inp[9]) ? node241 : node234;
							assign node234 = (inp[10]) ? 11'b00000111111 : node235;
								assign node235 = (inp[7]) ? 11'b00001111111 : node236;
									assign node236 = (inp[8]) ? 11'b00000111111 : 11'b00011111111;
							assign node241 = (inp[7]) ? node247 : node242;
								assign node242 = (inp[10]) ? node244 : 11'b00000111111;
									assign node244 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
								assign node247 = (inp[8]) ? 11'b00000001111 : node248;
									assign node248 = (inp[10]) ? 11'b00000001111 : 11'b00000111111;
					assign node252 = (inp[10]) ? node284 : node253;
						assign node253 = (inp[0]) ? node269 : node254;
							assign node254 = (inp[9]) ? node262 : node255;
								assign node255 = (inp[3]) ? node259 : node256;
									assign node256 = (inp[8]) ? 11'b00001111111 : 11'b00001111111;
									assign node259 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node262 = (inp[1]) ? node266 : node263;
									assign node263 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node266 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
							assign node269 = (inp[1]) ? node277 : node270;
								assign node270 = (inp[9]) ? node274 : node271;
									assign node271 = (inp[8]) ? 11'b00000111111 : 11'b00000111111;
									assign node274 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node277 = (inp[3]) ? node281 : node278;
									assign node278 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node281 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
						assign node284 = (inp[8]) ? node298 : node285;
							assign node285 = (inp[3]) ? node293 : node286;
								assign node286 = (inp[1]) ? node290 : node287;
									assign node287 = (inp[0]) ? 11'b00000111111 : 11'b00001111111;
									assign node290 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node293 = (inp[1]) ? 11'b00000000111 : node294;
									assign node294 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node298 = (inp[7]) ? node304 : node299;
								assign node299 = (inp[3]) ? node301 : 11'b00000011111;
									assign node301 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node304 = (inp[3]) ? node308 : node305;
									assign node305 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
									assign node308 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
				assign node311 = (inp[9]) ? node349 : node312;
					assign node312 = (inp[1]) ? node326 : node313;
						assign node313 = (inp[0]) ? node321 : node314;
							assign node314 = (inp[3]) ? node316 : 11'b00001111111;
								assign node316 = (inp[10]) ? 11'b00000111111 : node317;
									assign node317 = (inp[2]) ? 11'b00001111111 : 11'b00000111111;
							assign node321 = (inp[2]) ? node323 : 11'b00000111111;
								assign node323 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node326 = (inp[2]) ? node336 : node327;
							assign node327 = (inp[7]) ? node331 : node328;
								assign node328 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
								assign node331 = (inp[0]) ? 11'b00000000111 : node332;
									assign node332 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
							assign node336 = (inp[10]) ? node342 : node337;
								assign node337 = (inp[3]) ? node339 : 11'b00000111111;
									assign node339 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node342 = (inp[3]) ? node346 : node343;
									assign node343 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
									assign node346 = (inp[0]) ? 11'b00000000011 : 11'b00000001111;
					assign node349 = (inp[7]) ? node379 : node350;
						assign node350 = (inp[2]) ? node364 : node351;
							assign node351 = (inp[8]) ? node359 : node352;
								assign node352 = (inp[0]) ? node356 : node353;
									assign node353 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
									assign node356 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
								assign node359 = (inp[1]) ? 11'b00000011111 : node360;
									assign node360 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node364 = (inp[8]) ? node372 : node365;
								assign node365 = (inp[1]) ? node369 : node366;
									assign node366 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node369 = (inp[10]) ? 11'b00000001111 : 11'b00000001111;
								assign node372 = (inp[0]) ? node376 : node373;
									assign node373 = (inp[10]) ? 11'b00000001111 : 11'b00000001111;
									assign node376 = (inp[1]) ? 11'b00000000111 : 11'b00000000111;
						assign node379 = (inp[0]) ? node389 : node380;
							assign node380 = (inp[1]) ? node384 : node381;
								assign node381 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
								assign node384 = (inp[2]) ? 11'b00000001111 : node385;
									assign node385 = (inp[8]) ? 11'b00000001111 : 11'b00000001111;
							assign node389 = (inp[3]) ? node393 : node390;
								assign node390 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node393 = (inp[8]) ? node397 : node394;
									assign node394 = (inp[1]) ? 11'b00000000111 : 11'b00000001111;
									assign node397 = (inp[10]) ? 11'b00000000011 : 11'b00000000111;
		assign node400 = (inp[3]) ? node600 : node401;
			assign node401 = (inp[2]) ? node509 : node402;
				assign node402 = (inp[10]) ? node454 : node403;
					assign node403 = (inp[7]) ? node431 : node404;
						assign node404 = (inp[0]) ? node416 : node405;
							assign node405 = (inp[5]) ? node411 : node406;
								assign node406 = (inp[4]) ? 11'b00011111111 : node407;
									assign node407 = (inp[1]) ? 11'b00111111111 : 11'b00011111111;
								assign node411 = (inp[1]) ? node413 : 11'b00011111111;
									assign node413 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node416 = (inp[9]) ? node424 : node417;
								assign node417 = (inp[1]) ? node421 : node418;
									assign node418 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node421 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
								assign node424 = (inp[8]) ? node428 : node425;
									assign node425 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node428 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
						assign node431 = (inp[8]) ? node443 : node432;
							assign node432 = (inp[4]) ? node438 : node433;
								assign node433 = (inp[1]) ? node435 : 11'b00011111111;
									assign node435 = (inp[0]) ? 11'b00000111111 : 11'b00001111111;
								assign node438 = (inp[5]) ? 11'b00000111111 : node439;
									assign node439 = (inp[0]) ? 11'b00000111111 : 11'b00001111111;
							assign node443 = (inp[9]) ? node451 : node444;
								assign node444 = (inp[1]) ? node448 : node445;
									assign node445 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
									assign node448 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node451 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
					assign node454 = (inp[1]) ? node482 : node455;
						assign node455 = (inp[7]) ? node469 : node456;
							assign node456 = (inp[4]) ? node462 : node457;
								assign node457 = (inp[0]) ? node459 : 11'b00001111111;
									assign node459 = (inp[5]) ? 11'b00000111111 : 11'b00001111111;
								assign node462 = (inp[8]) ? node466 : node463;
									assign node463 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
									assign node466 = (inp[5]) ? 11'b00000011111 : 11'b00000111111;
							assign node469 = (inp[5]) ? node477 : node470;
								assign node470 = (inp[9]) ? node474 : node471;
									assign node471 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node474 = (inp[0]) ? 11'b00000011111 : 11'b00000111111;
								assign node477 = (inp[8]) ? node479 : 11'b00000011111;
									assign node479 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
						assign node482 = (inp[4]) ? node494 : node483;
							assign node483 = (inp[7]) ? node491 : node484;
								assign node484 = (inp[0]) ? node488 : node485;
									assign node485 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node488 = (inp[8]) ? 11'b00000011111 : 11'b00000011111;
								assign node491 = (inp[5]) ? 11'b00000011111 : 11'b00000001111;
							assign node494 = (inp[9]) ? node502 : node495;
								assign node495 = (inp[8]) ? node499 : node496;
									assign node496 = (inp[5]) ? 11'b00000011111 : 11'b00000111111;
									assign node499 = (inp[5]) ? 11'b00000001111 : 11'b00000011111;
								assign node502 = (inp[5]) ? node506 : node503;
									assign node503 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
									assign node506 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
				assign node509 = (inp[0]) ? node553 : node510;
					assign node510 = (inp[1]) ? node532 : node511;
						assign node511 = (inp[10]) ? node523 : node512;
							assign node512 = (inp[9]) ? node516 : node513;
								assign node513 = (inp[5]) ? 11'b00011111111 : 11'b00001111111;
								assign node516 = (inp[4]) ? node520 : node517;
									assign node517 = (inp[5]) ? 11'b00000111111 : 11'b00011111111;
									assign node520 = (inp[5]) ? 11'b00000011111 : 11'b00000111111;
							assign node523 = (inp[7]) ? node527 : node524;
								assign node524 = (inp[5]) ? 11'b00000111111 : 11'b00001111111;
								assign node527 = (inp[5]) ? 11'b00000011111 : node528;
									assign node528 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
						assign node532 = (inp[5]) ? node548 : node533;
							assign node533 = (inp[10]) ? node541 : node534;
								assign node534 = (inp[4]) ? node538 : node535;
									assign node535 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node538 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node541 = (inp[9]) ? node545 : node542;
									assign node542 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
									assign node545 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
							assign node548 = (inp[9]) ? 11'b00000001111 : node549;
								assign node549 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
					assign node553 = (inp[4]) ? node575 : node554;
						assign node554 = (inp[1]) ? node568 : node555;
							assign node555 = (inp[5]) ? node561 : node556;
								assign node556 = (inp[7]) ? 11'b00000111111 : node557;
									assign node557 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node561 = (inp[10]) ? node565 : node562;
									assign node562 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
									assign node565 = (inp[8]) ? 11'b00000011111 : 11'b00000011111;
							assign node568 = (inp[9]) ? 11'b00000001111 : node569;
								assign node569 = (inp[8]) ? node571 : 11'b00000111111;
									assign node571 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
						assign node575 = (inp[9]) ? node585 : node576;
							assign node576 = (inp[7]) ? node580 : node577;
								assign node577 = (inp[5]) ? 11'b00000011111 : 11'b00000111111;
								assign node580 = (inp[1]) ? node582 : 11'b00000001111;
									assign node582 = (inp[5]) ? 11'b00000000111 : 11'b00000001111;
							assign node585 = (inp[10]) ? node593 : node586;
								assign node586 = (inp[1]) ? node590 : node587;
									assign node587 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
									assign node590 = (inp[5]) ? 11'b00000001111 : 11'b00000011111;
								assign node593 = (inp[5]) ? node597 : node594;
									assign node594 = (inp[1]) ? 11'b00000000111 : 11'b00000000111;
									assign node597 = (inp[7]) ? 11'b00000000001 : 11'b00000000111;
			assign node600 = (inp[5]) ? node698 : node601;
				assign node601 = (inp[0]) ? node647 : node602;
					assign node602 = (inp[9]) ? node624 : node603;
						assign node603 = (inp[8]) ? node615 : node604;
							assign node604 = (inp[1]) ? node612 : node605;
								assign node605 = (inp[2]) ? node609 : node606;
									assign node606 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
									assign node609 = (inp[7]) ? 11'b00001111111 : 11'b00001111111;
								assign node612 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
							assign node615 = (inp[2]) ? 11'b00000011111 : node616;
								assign node616 = (inp[7]) ? node620 : node617;
									assign node617 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
									assign node620 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node624 = (inp[1]) ? node634 : node625;
							assign node625 = (inp[10]) ? 11'b00000011111 : node626;
								assign node626 = (inp[2]) ? node630 : node627;
									assign node627 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
									assign node630 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node634 = (inp[2]) ? node642 : node635;
								assign node635 = (inp[8]) ? node639 : node636;
									assign node636 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
									assign node639 = (inp[7]) ? 11'b00000001111 : 11'b00000001111;
								assign node642 = (inp[10]) ? node644 : 11'b00000001111;
									assign node644 = (inp[4]) ? 11'b00000000111 : 11'b00000001111;
					assign node647 = (inp[9]) ? node673 : node648;
						assign node648 = (inp[2]) ? node660 : node649;
							assign node649 = (inp[7]) ? node655 : node650;
								assign node650 = (inp[8]) ? 11'b00000011111 : node651;
									assign node651 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
								assign node655 = (inp[10]) ? 11'b00000001111 : node656;
									assign node656 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
							assign node660 = (inp[7]) ? node668 : node661;
								assign node661 = (inp[1]) ? node665 : node662;
									assign node662 = (inp[8]) ? 11'b00000111111 : 11'b00000011111;
									assign node665 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node668 = (inp[4]) ? node670 : 11'b00000001111;
									assign node670 = (inp[10]) ? 11'b00000000111 : 11'b00000001111;
						assign node673 = (inp[4]) ? node683 : node674;
							assign node674 = (inp[8]) ? node676 : 11'b00000011111;
								assign node676 = (inp[2]) ? node680 : node677;
									assign node677 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
									assign node680 = (inp[7]) ? 11'b00000000111 : 11'b00000000111;
							assign node683 = (inp[1]) ? node691 : node684;
								assign node684 = (inp[7]) ? node688 : node685;
									assign node685 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
									assign node688 = (inp[8]) ? 11'b00000000111 : 11'b00000001111;
								assign node691 = (inp[10]) ? node695 : node692;
									assign node692 = (inp[8]) ? 11'b00000000111 : 11'b00000000111;
									assign node695 = (inp[8]) ? 11'b00000000011 : 11'b00000000111;
				assign node698 = (inp[1]) ? node750 : node699;
					assign node699 = (inp[4]) ? node721 : node700;
						assign node700 = (inp[9]) ? node710 : node701;
							assign node701 = (inp[10]) ? node707 : node702;
								assign node702 = (inp[7]) ? node704 : 11'b00001111111;
									assign node704 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
								assign node707 = (inp[0]) ? 11'b00000011111 : 11'b00000111111;
							assign node710 = (inp[7]) ? node714 : node711;
								assign node711 = (inp[2]) ? 11'b00000001111 : 11'b00000111111;
								assign node714 = (inp[0]) ? node718 : node715;
									assign node715 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
									assign node718 = (inp[10]) ? 11'b00000000111 : 11'b00000001111;
						assign node721 = (inp[2]) ? node737 : node722;
							assign node722 = (inp[7]) ? node730 : node723;
								assign node723 = (inp[10]) ? node727 : node724;
									assign node724 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node727 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node730 = (inp[8]) ? node734 : node731;
									assign node731 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
									assign node734 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
							assign node737 = (inp[10]) ? node743 : node738;
								assign node738 = (inp[0]) ? node740 : 11'b00000001111;
									assign node740 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
								assign node743 = (inp[8]) ? node747 : node744;
									assign node744 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
									assign node747 = (inp[9]) ? 11'b00000000011 : 11'b00000000111;
					assign node750 = (inp[9]) ? node780 : node751;
						assign node751 = (inp[4]) ? node765 : node752;
							assign node752 = (inp[10]) ? node758 : node753;
								assign node753 = (inp[7]) ? node755 : 11'b00000011111;
									assign node755 = (inp[0]) ? 11'b00000001111 : 11'b00000011111;
								assign node758 = (inp[7]) ? node762 : node759;
									assign node759 = (inp[0]) ? 11'b00000001111 : 11'b00000001111;
									assign node762 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
							assign node765 = (inp[2]) ? node773 : node766;
								assign node766 = (inp[0]) ? node770 : node767;
									assign node767 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
									assign node770 = (inp[8]) ? 11'b00000000111 : 11'b00000001111;
								assign node773 = (inp[8]) ? node777 : node774;
									assign node774 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
									assign node777 = (inp[10]) ? 11'b00000000011 : 11'b00000000011;
						assign node780 = (inp[10]) ? node796 : node781;
							assign node781 = (inp[8]) ? node789 : node782;
								assign node782 = (inp[4]) ? node786 : node783;
									assign node783 = (inp[7]) ? 11'b00000001111 : 11'b00000001111;
									assign node786 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node789 = (inp[0]) ? node793 : node790;
									assign node790 = (inp[4]) ? 11'b00000000111 : 11'b00000011111;
									assign node793 = (inp[7]) ? 11'b00000000011 : 11'b00000000111;
							assign node796 = (inp[2]) ? node804 : node797;
								assign node797 = (inp[8]) ? node801 : node798;
									assign node798 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
									assign node801 = (inp[7]) ? 11'b00000000011 : 11'b00000000111;
								assign node804 = (inp[8]) ? node808 : node805;
									assign node805 = (inp[4]) ? 11'b00000000011 : 11'b00000000011;
									assign node808 = (inp[4]) ? 11'b00000000001 : 11'b00000000001;

endmodule