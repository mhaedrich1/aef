module dtc_split75_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node288;

	assign outp = (inp[3]) ? node206 : node1;
		assign node1 = (inp[9]) ? node77 : node2;
			assign node2 = (inp[4]) ? node52 : node3;
				assign node3 = (inp[0]) ? node23 : node4;
					assign node4 = (inp[6]) ? node10 : node5;
						assign node5 = (inp[5]) ? node7 : 3'b001;
							assign node7 = (inp[1]) ? 3'b001 : 3'b000;
						assign node10 = (inp[5]) ? 3'b000 : node11;
							assign node11 = (inp[7]) ? node13 : 3'b000;
								assign node13 = (inp[2]) ? node15 : 3'b000;
									assign node15 = (inp[8]) ? node17 : 3'b000;
										assign node17 = (inp[10]) ? node19 : 3'b000;
											assign node19 = (inp[1]) ? 3'b000 : 3'b000;
					assign node23 = (inp[6]) ? 3'b001 : node24;
						assign node24 = (inp[5]) ? node38 : node25;
							assign node25 = (inp[1]) ? 3'b000 : node26;
								assign node26 = (inp[8]) ? node32 : node27;
									assign node27 = (inp[11]) ? node29 : 3'b000;
										assign node29 = (inp[2]) ? 3'b000 : 3'b001;
									assign node32 = (inp[2]) ? node34 : 3'b000;
										assign node34 = (inp[11]) ? 3'b000 : 3'b001;
							assign node38 = (inp[1]) ? 3'b001 : node39;
								assign node39 = (inp[11]) ? node45 : node40;
									assign node40 = (inp[2]) ? node42 : 3'b000;
										assign node42 = (inp[8]) ? 3'b001 : 3'b000;
									assign node45 = (inp[2]) ? 3'b000 : node46;
										assign node46 = (inp[8]) ? 3'b000 : 3'b001;
				assign node52 = (inp[0]) ? node54 : 3'b000;
					assign node54 = (inp[1]) ? node72 : node55;
						assign node55 = (inp[5]) ? node65 : node56;
							assign node56 = (inp[6]) ? 3'b000 : node57;
								assign node57 = (inp[10]) ? node59 : 3'b000;
									assign node59 = (inp[2]) ? node61 : 3'b000;
										assign node61 = (inp[7]) ? 3'b001 : 3'b000;
							assign node65 = (inp[6]) ? 3'b001 : node66;
								assign node66 = (inp[10]) ? node68 : 3'b000;
									assign node68 = (inp[7]) ? 3'b001 : 3'b000;
						assign node72 = (inp[5]) ? 3'b000 : node73;
							assign node73 = (inp[6]) ? 3'b000 : 3'b001;
			assign node77 = (inp[6]) ? node169 : node78;
				assign node78 = (inp[4]) ? node140 : node79;
					assign node79 = (inp[0]) ? node89 : node80;
						assign node80 = (inp[5]) ? node86 : node81;
							assign node81 = (inp[7]) ? 3'b110 : node82;
								assign node82 = (inp[1]) ? 3'b110 : 3'b010;
							assign node86 = (inp[1]) ? 3'b010 : 3'b100;
						assign node89 = (inp[5]) ? node119 : node90;
							assign node90 = (inp[7]) ? node104 : node91;
								assign node91 = (inp[1]) ? 3'b001 : node92;
									assign node92 = (inp[2]) ? node98 : node93;
										assign node93 = (inp[11]) ? node95 : 3'b001;
											assign node95 = (inp[8]) ? 3'b001 : 3'b110;
										assign node98 = (inp[8]) ? node100 : 3'b001;
											assign node100 = (inp[11]) ? 3'b001 : 3'b110;
								assign node104 = (inp[1]) ? 3'b101 : node105;
									assign node105 = (inp[10]) ? node111 : node106;
										assign node106 = (inp[11]) ? node108 : 3'b001;
											assign node108 = (inp[2]) ? 3'b001 : 3'b000;
										assign node111 = (inp[2]) ? node115 : node112;
											assign node112 = (inp[11]) ? 3'b110 : 3'b001;
											assign node115 = (inp[8]) ? 3'b000 : 3'b001;
							assign node119 = (inp[1]) ? 3'b110 : node120;
								assign node120 = (inp[10]) ? node128 : node121;
									assign node121 = (inp[11]) ? 3'b001 : node122;
										assign node122 = (inp[2]) ? node124 : 3'b001;
											assign node124 = (inp[8]) ? 3'b110 : 3'b001;
									assign node128 = (inp[8]) ? node134 : node129;
										assign node129 = (inp[11]) ? node131 : 3'b001;
											assign node131 = (inp[2]) ? 3'b001 : 3'b110;
										assign node134 = (inp[11]) ? 3'b001 : node135;
											assign node135 = (inp[2]) ? 3'b110 : 3'b001;
					assign node140 = (inp[0]) ? node152 : node141;
						assign node141 = (inp[5]) ? 3'b000 : node142;
							assign node142 = (inp[1]) ? node144 : 3'b000;
								assign node144 = (inp[10]) ? node146 : 3'b000;
									assign node146 = (inp[7]) ? 3'b000 : node147;
										assign node147 = (inp[2]) ? 3'b100 : 3'b000;
						assign node152 = (inp[5]) ? node162 : node153;
							assign node153 = (inp[1]) ? 3'b010 : node154;
								assign node154 = (inp[2]) ? node156 : 3'b100;
									assign node156 = (inp[7]) ? node158 : 3'b100;
										assign node158 = (inp[10]) ? 3'b010 : 3'b100;
							assign node162 = (inp[7]) ? node164 : 3'b100;
								assign node164 = (inp[1]) ? 3'b100 : node165;
									assign node165 = (inp[10]) ? 3'b010 : 3'b100;
				assign node169 = (inp[0]) ? node171 : 3'b001;
					assign node171 = (inp[4]) ? node189 : node172;
						assign node172 = (inp[5]) ? node182 : node173;
							assign node173 = (inp[1]) ? 3'b111 : node174;
								assign node174 = (inp[10]) ? node176 : 3'b011;
									assign node176 = (inp[2]) ? node178 : 3'b011;
										assign node178 = (inp[7]) ? 3'b111 : 3'b011;
							assign node182 = (inp[7]) ? node184 : 3'b011;
								assign node184 = (inp[10]) ? node186 : 3'b011;
									assign node186 = (inp[1]) ? 3'b011 : 3'b111;
						assign node189 = (inp[5]) ? node199 : node190;
							assign node190 = (inp[1]) ? 3'b101 : node191;
								assign node191 = (inp[7]) ? node193 : 3'b001;
									assign node193 = (inp[2]) ? node195 : 3'b001;
										assign node195 = (inp[10]) ? 3'b101 : 3'b001;
							assign node199 = (inp[1]) ? 3'b001 : node200;
								assign node200 = (inp[7]) ? node202 : 3'b010;
									assign node202 = (inp[10]) ? 3'b110 : 3'b010;
		assign node206 = (inp[6]) ? node208 : 3'b000;
			assign node208 = (inp[0]) ? node224 : node209;
				assign node209 = (inp[4]) ? node213 : node210;
					assign node210 = (inp[9]) ? 3'b100 : 3'b000;
					assign node213 = (inp[9]) ? 3'b000 : node214;
						assign node214 = (inp[10]) ? node216 : 3'b010;
							assign node216 = (inp[1]) ? node218 : 3'b010;
								assign node218 = (inp[2]) ? 3'b100 : node219;
									assign node219 = (inp[5]) ? 3'b100 : 3'b010;
				assign node224 = (inp[4]) ? node240 : node225;
					assign node225 = (inp[9]) ? node227 : 3'b001;
						assign node227 = (inp[7]) ? node229 : 3'b010;
							assign node229 = (inp[1]) ? node231 : 3'b010;
								assign node231 = (inp[10]) ? node233 : 3'b010;
									assign node233 = (inp[8]) ? node235 : 3'b010;
										assign node235 = (inp[5]) ? 3'b010 : node236;
											assign node236 = (inp[11]) ? 3'b110 : 3'b010;
					assign node240 = (inp[9]) ? node274 : node241;
						assign node241 = (inp[1]) ? node251 : node242;
							assign node242 = (inp[7]) ? node244 : 3'b010;
								assign node244 = (inp[10]) ? 3'b010 : node245;
									assign node245 = (inp[11]) ? node247 : 3'b110;
										assign node247 = (inp[2]) ? 3'b110 : 3'b010;
							assign node251 = (inp[7]) ? node253 : 3'b110;
								assign node253 = (inp[10]) ? node263 : node254;
									assign node254 = (inp[2]) ? node260 : node255;
										assign node255 = (inp[11]) ? node257 : 3'b110;
											assign node257 = (inp[8]) ? 3'b110 : 3'b010;
										assign node260 = (inp[11]) ? 3'b110 : 3'b001;
									assign node263 = (inp[8]) ? node269 : node264;
										assign node264 = (inp[11]) ? node266 : 3'b010;
											assign node266 = (inp[2]) ? 3'b010 : 3'b110;
										assign node269 = (inp[2]) ? node271 : 3'b010;
											assign node271 = (inp[11]) ? 3'b010 : 3'b110;
						assign node274 = (inp[7]) ? node276 : 3'b000;
							assign node276 = (inp[10]) ? 3'b000 : node277;
								assign node277 = (inp[11]) ? node285 : node278;
									assign node278 = (inp[8]) ? node280 : 3'b100;
										assign node280 = (inp[1]) ? node282 : 3'b100;
											assign node282 = (inp[2]) ? 3'b010 : 3'b100;
									assign node285 = (inp[1]) ? node287 : 3'b000;
										assign node287 = (inp[8]) ? 3'b100 : node288;
											assign node288 = (inp[2]) ? 3'b100 : 3'b000;

endmodule