module dtc_split75_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node887;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node947;
	wire [3-1:0] node949;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1074;
	wire [3-1:0] node1077;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1097;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1105;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1120;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1142;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1161;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1171;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1186;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1194;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1237;
	wire [3-1:0] node1239;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1246;
	wire [3-1:0] node1249;
	wire [3-1:0] node1251;
	wire [3-1:0] node1254;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1265;
	wire [3-1:0] node1267;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1280;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1292;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1320;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;

	assign outp = (inp[6]) ? node798 : node1;
		assign node1 = (inp[3]) ? node363 : node2;
			assign node2 = (inp[7]) ? node90 : node3;
				assign node3 = (inp[9]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node30 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[5]) ? node22 : node7;
								assign node7 = (inp[11]) ? node15 : node8;
									assign node8 = (inp[0]) ? node10 : 3'b101;
										assign node10 = (inp[1]) ? node12 : 3'b101;
											assign node12 = (inp[8]) ? 3'b011 : 3'b101;
									assign node15 = (inp[8]) ? 3'b011 : node16;
										assign node16 = (inp[0]) ? node18 : 3'b101;
											assign node18 = (inp[2]) ? 3'b011 : 3'b101;
								assign node22 = (inp[11]) ? node24 : 3'b011;
									assign node24 = (inp[8]) ? 3'b101 : node25;
										assign node25 = (inp[2]) ? 3'b101 : 3'b011;
						assign node30 = (inp[10]) ? node50 : node31;
							assign node31 = (inp[8]) ? node41 : node32;
								assign node32 = (inp[11]) ? node34 : 3'b010;
									assign node34 = (inp[2]) ? 3'b110 : node35;
										assign node35 = (inp[1]) ? 3'b110 : node36;
											assign node36 = (inp[0]) ? 3'b110 : 3'b001;
								assign node41 = (inp[11]) ? node43 : 3'b100;
									assign node43 = (inp[1]) ? 3'b010 : node44;
										assign node44 = (inp[0]) ? 3'b110 : node45;
											assign node45 = (inp[2]) ? 3'b110 : 3'b101;
							assign node50 = (inp[11]) ? node78 : node51;
								assign node51 = (inp[8]) ? node67 : node52;
									assign node52 = (inp[1]) ? node60 : node53;
										assign node53 = (inp[2]) ? 3'b101 : node54;
											assign node54 = (inp[0]) ? node56 : 3'b101;
												assign node56 = (inp[5]) ? 3'b001 : 3'b101;
										assign node60 = (inp[2]) ? 3'b001 : node61;
											assign node61 = (inp[5]) ? node63 : 3'b101;
												assign node63 = (inp[0]) ? 3'b001 : 3'b101;
									assign node67 = (inp[0]) ? node73 : node68;
										assign node68 = (inp[1]) ? node70 : 3'b001;
											assign node70 = (inp[2]) ? 3'b110 : 3'b001;
										assign node73 = (inp[5]) ? 3'b110 : node74;
											assign node74 = (inp[2]) ? 3'b110 : 3'b001;
								assign node78 = (inp[8]) ? node84 : node79;
									assign node79 = (inp[5]) ? node81 : 3'b011;
										assign node81 = (inp[0]) ? 3'b101 : 3'b011;
									assign node84 = (inp[0]) ? node86 : 3'b101;
										assign node86 = (inp[5]) ? 3'b001 : 3'b101;
				assign node90 = (inp[10]) ? node238 : node91;
					assign node91 = (inp[4]) ? node173 : node92;
						assign node92 = (inp[9]) ? node142 : node93;
							assign node93 = (inp[11]) ? node115 : node94;
								assign node94 = (inp[8]) ? node104 : node95;
									assign node95 = (inp[1]) ? node97 : 3'b110;
										assign node97 = (inp[0]) ? node101 : node98;
											assign node98 = (inp[5]) ? 3'b110 : 3'b010;
											assign node101 = (inp[5]) ? 3'b010 : 3'b110;
									assign node104 = (inp[5]) ? node108 : node105;
										assign node105 = (inp[2]) ? 3'b010 : 3'b110;
										assign node108 = (inp[2]) ? node110 : 3'b000;
											assign node110 = (inp[1]) ? node112 : 3'b000;
												assign node112 = (inp[0]) ? 3'b100 : 3'b000;
								assign node115 = (inp[8]) ? node133 : node116;
									assign node116 = (inp[5]) ? node122 : node117;
										assign node117 = (inp[0]) ? node119 : 3'b111;
											assign node119 = (inp[2]) ? 3'b001 : 3'b011;
										assign node122 = (inp[2]) ? node128 : node123;
											assign node123 = (inp[0]) ? node125 : 3'b001;
												assign node125 = (inp[1]) ? 3'b100 : 3'b001;
											assign node128 = (inp[0]) ? node130 : 3'b011;
												assign node130 = (inp[1]) ? 3'b110 : 3'b011;
									assign node133 = (inp[5]) ? 3'b110 : node134;
										assign node134 = (inp[2]) ? node136 : 3'b001;
											assign node136 = (inp[0]) ? node138 : 3'b101;
												assign node138 = (inp[1]) ? 3'b110 : 3'b101;
							assign node142 = (inp[5]) ? node166 : node143;
								assign node143 = (inp[8]) ? node153 : node144;
									assign node144 = (inp[11]) ? node146 : 3'b110;
										assign node146 = (inp[1]) ? node148 : 3'b110;
											assign node148 = (inp[0]) ? node150 : 3'b110;
												assign node150 = (inp[2]) ? 3'b000 : 3'b110;
									assign node153 = (inp[11]) ? node159 : node154;
										assign node154 = (inp[0]) ? node156 : 3'b110;
											assign node156 = (inp[1]) ? 3'b000 : 3'b110;
										assign node159 = (inp[0]) ? node161 : 3'b000;
											assign node161 = (inp[2]) ? node163 : 3'b000;
												assign node163 = (inp[1]) ? 3'b110 : 3'b000;
								assign node166 = (inp[11]) ? node168 : 3'b000;
									assign node168 = (inp[2]) ? 3'b110 : node169;
										assign node169 = (inp[8]) ? 3'b110 : 3'b000;
						assign node173 = (inp[9]) ? node201 : node174;
							assign node174 = (inp[11]) ? node182 : node175;
								assign node175 = (inp[5]) ? 3'b000 : node176;
									assign node176 = (inp[8]) ? node178 : 3'b100;
										assign node178 = (inp[1]) ? 3'b000 : 3'b100;
								assign node182 = (inp[8]) ? node192 : node183;
									assign node183 = (inp[2]) ? node187 : node184;
										assign node184 = (inp[1]) ? 3'b010 : 3'b100;
										assign node187 = (inp[5]) ? node189 : 3'b010;
											assign node189 = (inp[1]) ? 3'b100 : 3'b010;
									assign node192 = (inp[1]) ? node196 : node193;
										assign node193 = (inp[2]) ? 3'b100 : 3'b000;
										assign node196 = (inp[5]) ? node198 : 3'b100;
											assign node198 = (inp[2]) ? 3'b000 : 3'b100;
							assign node201 = (inp[8]) ? node221 : node202;
								assign node202 = (inp[11]) ? node204 : 3'b001;
									assign node204 = (inp[1]) ? node212 : node205;
										assign node205 = (inp[2]) ? node209 : node206;
											assign node206 = (inp[5]) ? 3'b010 : 3'b011;
											assign node209 = (inp[0]) ? 3'b100 : 3'b101;
										assign node212 = (inp[2]) ? node216 : node213;
											assign node213 = (inp[5]) ? 3'b100 : 3'b101;
											assign node216 = (inp[0]) ? node218 : 3'b101;
												assign node218 = (inp[5]) ? 3'b101 : 3'b100;
								assign node221 = (inp[11]) ? node225 : node222;
									assign node222 = (inp[5]) ? 3'b110 : 3'b111;
									assign node225 = (inp[1]) ? node233 : node226;
										assign node226 = (inp[5]) ? 3'b101 : node227;
											assign node227 = (inp[0]) ? 3'b100 : node228;
												assign node228 = (inp[2]) ? 3'b100 : 3'b110;
										assign node233 = (inp[2]) ? 3'b001 : node234;
											assign node234 = (inp[5]) ? 3'b001 : 3'b000;
					assign node238 = (inp[4]) ? node290 : node239;
						assign node239 = (inp[9]) ? 3'b100 : node240;
							assign node240 = (inp[8]) ? node262 : node241;
								assign node241 = (inp[11]) ? node251 : node242;
									assign node242 = (inp[5]) ? node246 : node243;
										assign node243 = (inp[0]) ? 3'b101 : 3'b001;
										assign node246 = (inp[0]) ? node248 : 3'b101;
											assign node248 = (inp[1]) ? 3'b001 : 3'b101;
									assign node251 = (inp[0]) ? node255 : node252;
										assign node252 = (inp[5]) ? 3'b011 : 3'b101;
										assign node255 = (inp[5]) ? node259 : node256;
											assign node256 = (inp[2]) ? 3'b011 : 3'b001;
											assign node259 = (inp[2]) ? 3'b101 : 3'b111;
								assign node262 = (inp[11]) ? node274 : node263;
									assign node263 = (inp[5]) ? node267 : node264;
										assign node264 = (inp[2]) ? 3'b001 : 3'b101;
										assign node267 = (inp[0]) ? node269 : 3'b010;
											assign node269 = (inp[2]) ? node271 : 3'b010;
												assign node271 = (inp[1]) ? 3'b110 : 3'b010;
									assign node274 = (inp[5]) ? node282 : node275;
										assign node275 = (inp[2]) ? node277 : 3'b011;
											assign node277 = (inp[1]) ? node279 : 3'b111;
												assign node279 = (inp[0]) ? 3'b101 : 3'b111;
										assign node282 = (inp[2]) ? node284 : 3'b101;
											assign node284 = (inp[0]) ? node286 : 3'b101;
												assign node286 = (inp[1]) ? 3'b001 : 3'b101;
						assign node290 = (inp[9]) ? node324 : node291;
							assign node291 = (inp[11]) ? node303 : node292;
								assign node292 = (inp[8]) ? node298 : node293;
									assign node293 = (inp[5]) ? node295 : 3'b110;
										assign node295 = (inp[0]) ? 3'b010 : 3'b110;
									assign node298 = (inp[0]) ? node300 : 3'b010;
										assign node300 = (inp[5]) ? 3'b100 : 3'b010;
								assign node303 = (inp[2]) ? node317 : node304;
									assign node304 = (inp[5]) ? node310 : node305;
										assign node305 = (inp[0]) ? node307 : 3'b001;
											assign node307 = (inp[8]) ? 3'b101 : 3'b001;
										assign node310 = (inp[8]) ? 3'b110 : node311;
											assign node311 = (inp[1]) ? node313 : 3'b001;
												assign node313 = (inp[0]) ? 3'b110 : 3'b001;
									assign node317 = (inp[5]) ? 3'b110 : node318;
										assign node318 = (inp[8]) ? node320 : 3'b001;
											assign node320 = (inp[0]) ? 3'b110 : 3'b010;
							assign node324 = (inp[11]) ? node348 : node325;
								assign node325 = (inp[8]) ? node339 : node326;
									assign node326 = (inp[1]) ? node332 : node327;
										assign node327 = (inp[5]) ? node329 : 3'b111;
											assign node329 = (inp[0]) ? 3'b011 : 3'b111;
										assign node332 = (inp[2]) ? 3'b011 : node333;
											assign node333 = (inp[0]) ? node335 : 3'b111;
												assign node335 = (inp[5]) ? 3'b011 : 3'b111;
									assign node339 = (inp[2]) ? node345 : node340;
										assign node340 = (inp[0]) ? node342 : 3'b011;
											assign node342 = (inp[5]) ? 3'b101 : 3'b011;
										assign node345 = (inp[1]) ? 3'b101 : 3'b011;
								assign node348 = (inp[8]) ? node358 : node349;
									assign node349 = (inp[1]) ? node351 : 3'b001;
										assign node351 = (inp[2]) ? node353 : 3'b111;
											assign node353 = (inp[5]) ? node355 : 3'b001;
												assign node355 = (inp[0]) ? 3'b111 : 3'b001;
									assign node358 = (inp[5]) ? node360 : 3'b111;
										assign node360 = (inp[0]) ? 3'b011 : 3'b111;
			assign node363 = (inp[9]) ? node515 : node364;
				assign node364 = (inp[4]) ? node504 : node365;
					assign node365 = (inp[7]) ? node465 : node366;
						assign node366 = (inp[10]) ? node412 : node367;
							assign node367 = (inp[11]) ? node379 : node368;
								assign node368 = (inp[8]) ? 3'b000 : node369;
									assign node369 = (inp[0]) ? node371 : 3'b100;
										assign node371 = (inp[2]) ? 3'b000 : node372;
											assign node372 = (inp[5]) ? node374 : 3'b100;
												assign node374 = (inp[1]) ? 3'b000 : 3'b100;
								assign node379 = (inp[8]) ? node397 : node380;
									assign node380 = (inp[1]) ? node386 : node381;
										assign node381 = (inp[5]) ? 3'b010 : node382;
											assign node382 = (inp[0]) ? 3'b010 : 3'b110;
										assign node386 = (inp[2]) ? node392 : node387;
											assign node387 = (inp[0]) ? 3'b010 : node388;
												assign node388 = (inp[5]) ? 3'b010 : 3'b110;
											assign node392 = (inp[0]) ? 3'b100 : node393;
												assign node393 = (inp[5]) ? 3'b010 : 3'b110;
									assign node397 = (inp[5]) ? node405 : node398;
										assign node398 = (inp[2]) ? node400 : 3'b010;
											assign node400 = (inp[0]) ? node402 : 3'b110;
												assign node402 = (inp[1]) ? 3'b100 : 3'b110;
										assign node405 = (inp[1]) ? node407 : 3'b100;
											assign node407 = (inp[0]) ? node409 : 3'b100;
												assign node409 = (inp[2]) ? 3'b000 : 3'b100;
							assign node412 = (inp[11]) ? node434 : node413;
								assign node413 = (inp[8]) ? node423 : node414;
									assign node414 = (inp[5]) ? node418 : node415;
										assign node415 = (inp[0]) ? 3'b110 : 3'b010;
										assign node418 = (inp[0]) ? node420 : 3'b110;
											assign node420 = (inp[1]) ? 3'b010 : 3'b110;
									assign node423 = (inp[5]) ? node427 : node424;
										assign node424 = (inp[2]) ? 3'b010 : 3'b110;
										assign node427 = (inp[1]) ? node429 : 3'b000;
											assign node429 = (inp[2]) ? node431 : 3'b000;
												assign node431 = (inp[0]) ? 3'b100 : 3'b000;
								assign node434 = (inp[5]) ? node448 : node435;
									assign node435 = (inp[0]) ? node441 : node436;
										assign node436 = (inp[8]) ? node438 : 3'b111;
											assign node438 = (inp[2]) ? 3'b101 : 3'b001;
										assign node441 = (inp[8]) ? node445 : node442;
											assign node442 = (inp[2]) ? 3'b001 : 3'b011;
											assign node445 = (inp[2]) ? 3'b110 : 3'b001;
									assign node448 = (inp[8]) ? node460 : node449;
										assign node449 = (inp[2]) ? node455 : node450;
											assign node450 = (inp[1]) ? node452 : 3'b001;
												assign node452 = (inp[0]) ? 3'b100 : 3'b001;
											assign node455 = (inp[0]) ? node457 : 3'b011;
												assign node457 = (inp[1]) ? 3'b110 : 3'b011;
										assign node460 = (inp[1]) ? node462 : 3'b110;
											assign node462 = (inp[2]) ? 3'b010 : 3'b110;
						assign node465 = (inp[10]) ? node467 : 3'b000;
							assign node467 = (inp[11]) ? node475 : node468;
								assign node468 = (inp[8]) ? 3'b000 : node469;
									assign node469 = (inp[5]) ? node471 : 3'b100;
										assign node471 = (inp[0]) ? 3'b000 : 3'b100;
								assign node475 = (inp[8]) ? node495 : node476;
									assign node476 = (inp[0]) ? node486 : node477;
										assign node477 = (inp[5]) ? node481 : node478;
											assign node478 = (inp[2]) ? 3'b010 : 3'b000;
											assign node481 = (inp[2]) ? node483 : 3'b010;
												assign node483 = (inp[1]) ? 3'b000 : 3'b010;
										assign node486 = (inp[5]) ? node488 : 3'b010;
											assign node488 = (inp[2]) ? node492 : node489;
												assign node489 = (inp[1]) ? 3'b110 : 3'b000;
												assign node492 = (inp[1]) ? 3'b100 : 3'b110;
									assign node495 = (inp[5]) ? node499 : node496;
										assign node496 = (inp[0]) ? 3'b100 : 3'b000;
										assign node499 = (inp[1]) ? node501 : 3'b100;
											assign node501 = (inp[0]) ? 3'b000 : 3'b100;
					assign node504 = (inp[7]) ? 3'b000 : node505;
						assign node505 = (inp[11]) ? node507 : 3'b000;
							assign node507 = (inp[10]) ? node509 : 3'b000;
								assign node509 = (inp[5]) ? node511 : 3'b100;
									assign node511 = (inp[8]) ? 3'b000 : 3'b100;
				assign node515 = (inp[4]) ? node661 : node516;
					assign node516 = (inp[7]) ? node542 : node517;
						assign node517 = (inp[10]) ? 3'b111 : node518;
							assign node518 = (inp[11]) ? node526 : node519;
								assign node519 = (inp[5]) ? 3'b011 : node520;
									assign node520 = (inp[8]) ? node522 : 3'b101;
										assign node522 = (inp[1]) ? 3'b011 : 3'b101;
								assign node526 = (inp[5]) ? node536 : node527;
									assign node527 = (inp[8]) ? node529 : 3'b101;
										assign node529 = (inp[0]) ? node531 : 3'b011;
											assign node531 = (inp[2]) ? node533 : 3'b011;
												assign node533 = (inp[1]) ? 3'b101 : 3'b011;
									assign node536 = (inp[8]) ? 3'b101 : node537;
										assign node537 = (inp[2]) ? 3'b101 : 3'b011;
						assign node542 = (inp[10]) ? node604 : node543;
							assign node543 = (inp[11]) ? node577 : node544;
								assign node544 = (inp[8]) ? node566 : node545;
									assign node545 = (inp[1]) ? node551 : node546;
										assign node546 = (inp[5]) ? 3'b110 : node547;
											assign node547 = (inp[0]) ? 3'b110 : 3'b010;
										assign node551 = (inp[2]) ? node559 : node552;
											assign node552 = (inp[5]) ? node556 : node553;
												assign node553 = (inp[0]) ? 3'b110 : 3'b010;
												assign node556 = (inp[0]) ? 3'b010 : 3'b110;
											assign node559 = (inp[5]) ? node563 : node560;
												assign node560 = (inp[0]) ? 3'b110 : 3'b010;
												assign node563 = (inp[0]) ? 3'b010 : 3'b110;
									assign node566 = (inp[5]) ? node570 : node567;
										assign node567 = (inp[2]) ? 3'b010 : 3'b110;
										assign node570 = (inp[0]) ? node572 : 3'b000;
											assign node572 = (inp[1]) ? node574 : 3'b000;
												assign node574 = (inp[2]) ? 3'b100 : 3'b000;
								assign node577 = (inp[8]) ? node595 : node578;
									assign node578 = (inp[5]) ? node584 : node579;
										assign node579 = (inp[0]) ? node581 : 3'b111;
											assign node581 = (inp[2]) ? 3'b001 : 3'b011;
										assign node584 = (inp[2]) ? node590 : node585;
											assign node585 = (inp[1]) ? node587 : 3'b001;
												assign node587 = (inp[0]) ? 3'b100 : 3'b001;
											assign node590 = (inp[1]) ? node592 : 3'b011;
												assign node592 = (inp[0]) ? 3'b110 : 3'b011;
									assign node595 = (inp[5]) ? 3'b110 : node596;
										assign node596 = (inp[2]) ? node598 : 3'b001;
											assign node598 = (inp[1]) ? node600 : 3'b101;
												assign node600 = (inp[0]) ? 3'b110 : 3'b101;
							assign node604 = (inp[8]) ? node638 : node605;
								assign node605 = (inp[11]) ? node623 : node606;
									assign node606 = (inp[1]) ? node610 : node607;
										assign node607 = (inp[0]) ? 3'b101 : 3'b001;
										assign node610 = (inp[2]) ? node618 : node611;
											assign node611 = (inp[0]) ? node615 : node612;
												assign node612 = (inp[5]) ? 3'b101 : 3'b001;
												assign node615 = (inp[5]) ? 3'b001 : 3'b101;
											assign node618 = (inp[5]) ? node620 : 3'b001;
												assign node620 = (inp[0]) ? 3'b001 : 3'b101;
									assign node623 = (inp[0]) ? node629 : node624;
										assign node624 = (inp[5]) ? node626 : 3'b101;
											assign node626 = (inp[2]) ? 3'b001 : 3'b011;
										assign node629 = (inp[5]) ? node633 : node630;
											assign node630 = (inp[2]) ? 3'b011 : 3'b001;
											assign node633 = (inp[1]) ? node635 : 3'b001;
												assign node635 = (inp[2]) ? 3'b101 : 3'b111;
								assign node638 = (inp[11]) ? node648 : node639;
									assign node639 = (inp[5]) ? node643 : node640;
										assign node640 = (inp[2]) ? 3'b001 : 3'b101;
										assign node643 = (inp[0]) ? node645 : 3'b010;
											assign node645 = (inp[2]) ? 3'b110 : 3'b010;
									assign node648 = (inp[5]) ? node656 : node649;
										assign node649 = (inp[2]) ? node651 : 3'b011;
											assign node651 = (inp[0]) ? node653 : 3'b111;
												assign node653 = (inp[1]) ? 3'b101 : 3'b111;
										assign node656 = (inp[0]) ? node658 : 3'b101;
											assign node658 = (inp[2]) ? 3'b001 : 3'b101;
					assign node661 = (inp[10]) ? node729 : node662;
						assign node662 = (inp[7]) ? node682 : node663;
							assign node663 = (inp[8]) ? node673 : node664;
								assign node664 = (inp[11]) ? node666 : 3'b010;
									assign node666 = (inp[0]) ? 3'b110 : node667;
										assign node667 = (inp[1]) ? 3'b110 : node668;
											assign node668 = (inp[2]) ? 3'b110 : 3'b001;
								assign node673 = (inp[11]) ? node675 : 3'b100;
									assign node675 = (inp[1]) ? 3'b010 : node676;
										assign node676 = (inp[0]) ? 3'b110 : node677;
											assign node677 = (inp[2]) ? 3'b110 : 3'b101;
							assign node682 = (inp[5]) ? node702 : node683;
								assign node683 = (inp[11]) ? node691 : node684;
									assign node684 = (inp[1]) ? node686 : 3'b100;
										assign node686 = (inp[0]) ? node688 : 3'b100;
											assign node688 = (inp[8]) ? 3'b000 : 3'b100;
									assign node691 = (inp[8]) ? node697 : node692;
										assign node692 = (inp[1]) ? 3'b010 : node693;
											assign node693 = (inp[2]) ? 3'b010 : 3'b100;
										assign node697 = (inp[2]) ? 3'b100 : node698;
											assign node698 = (inp[1]) ? 3'b100 : 3'b000;
								assign node702 = (inp[11]) ? node704 : 3'b000;
									assign node704 = (inp[8]) ? node718 : node705;
										assign node705 = (inp[0]) ? node713 : node706;
											assign node706 = (inp[1]) ? node710 : node707;
												assign node707 = (inp[2]) ? 3'b010 : 3'b100;
												assign node710 = (inp[2]) ? 3'b100 : 3'b010;
											assign node713 = (inp[2]) ? node715 : 3'b010;
												assign node715 = (inp[1]) ? 3'b100 : 3'b010;
										assign node718 = (inp[0]) ? node724 : node719;
											assign node719 = (inp[1]) ? node721 : 3'b100;
												assign node721 = (inp[2]) ? 3'b000 : 3'b100;
											assign node724 = (inp[2]) ? 3'b100 : node725;
												assign node725 = (inp[1]) ? 3'b100 : 3'b000;
						assign node729 = (inp[7]) ? node763 : node730;
							assign node730 = (inp[11]) ? node752 : node731;
								assign node731 = (inp[8]) ? node747 : node732;
									assign node732 = (inp[1]) ? node740 : node733;
										assign node733 = (inp[0]) ? node735 : 3'b101;
											assign node735 = (inp[2]) ? 3'b101 : node736;
												assign node736 = (inp[5]) ? 3'b001 : 3'b101;
										assign node740 = (inp[2]) ? 3'b001 : node741;
											assign node741 = (inp[0]) ? node743 : 3'b101;
												assign node743 = (inp[5]) ? 3'b001 : 3'b101;
									assign node747 = (inp[0]) ? node749 : 3'b001;
										assign node749 = (inp[5]) ? 3'b110 : 3'b001;
								assign node752 = (inp[8]) ? node758 : node753;
									assign node753 = (inp[5]) ? node755 : 3'b011;
										assign node755 = (inp[0]) ? 3'b101 : 3'b011;
									assign node758 = (inp[0]) ? node760 : 3'b101;
										assign node760 = (inp[5]) ? 3'b001 : 3'b101;
							assign node763 = (inp[11]) ? node775 : node764;
								assign node764 = (inp[8]) ? node770 : node765;
									assign node765 = (inp[0]) ? node767 : 3'b110;
										assign node767 = (inp[5]) ? 3'b010 : 3'b110;
									assign node770 = (inp[0]) ? node772 : 3'b010;
										assign node772 = (inp[5]) ? 3'b100 : 3'b010;
								assign node775 = (inp[8]) ? node781 : node776;
									assign node776 = (inp[0]) ? node778 : 3'b001;
										assign node778 = (inp[5]) ? 3'b110 : 3'b001;
									assign node781 = (inp[2]) ? node789 : node782;
										assign node782 = (inp[5]) ? node786 : node783;
											assign node783 = (inp[0]) ? 3'b101 : 3'b001;
											assign node786 = (inp[0]) ? 3'b010 : 3'b110;
										assign node789 = (inp[0]) ? node793 : node790;
											assign node790 = (inp[5]) ? 3'b110 : 3'b010;
											assign node793 = (inp[5]) ? node795 : 3'b110;
												assign node795 = (inp[1]) ? 3'b010 : 3'b110;
		assign node798 = (inp[9]) ? node954 : node799;
			assign node799 = (inp[3]) ? 3'b000 : node800;
				assign node800 = (inp[4]) ? node916 : node801;
					assign node801 = (inp[7]) ? node879 : node802;
						assign node802 = (inp[10]) ? node838 : node803;
							assign node803 = (inp[11]) ? node813 : node804;
								assign node804 = (inp[8]) ? 3'b000 : node805;
									assign node805 = (inp[0]) ? node807 : 3'b100;
										assign node807 = (inp[5]) ? node809 : 3'b100;
											assign node809 = (inp[2]) ? 3'b000 : 3'b100;
								assign node813 = (inp[5]) ? node829 : node814;
									assign node814 = (inp[2]) ? node820 : node815;
										assign node815 = (inp[0]) ? 3'b010 : node816;
											assign node816 = (inp[8]) ? 3'b010 : 3'b110;
										assign node820 = (inp[8]) ? node824 : node821;
											assign node821 = (inp[0]) ? 3'b010 : 3'b110;
											assign node824 = (inp[0]) ? node826 : 3'b110;
												assign node826 = (inp[1]) ? 3'b100 : 3'b110;
									assign node829 = (inp[8]) ? node833 : node830;
										assign node830 = (inp[1]) ? 3'b100 : 3'b010;
										assign node833 = (inp[1]) ? node835 : 3'b100;
											assign node835 = (inp[2]) ? 3'b000 : 3'b100;
							assign node838 = (inp[11]) ? node858 : node839;
								assign node839 = (inp[8]) ? node853 : node840;
									assign node840 = (inp[1]) ? node846 : node841;
										assign node841 = (inp[5]) ? 3'b110 : node842;
											assign node842 = (inp[0]) ? 3'b110 : 3'b010;
										assign node846 = (inp[5]) ? node850 : node847;
											assign node847 = (inp[0]) ? 3'b110 : 3'b010;
											assign node850 = (inp[0]) ? 3'b010 : 3'b110;
									assign node853 = (inp[5]) ? 3'b000 : node854;
										assign node854 = (inp[2]) ? 3'b010 : 3'b110;
								assign node858 = (inp[5]) ? node868 : node859;
									assign node859 = (inp[8]) ? node865 : node860;
										assign node860 = (inp[0]) ? node862 : 3'b111;
											assign node862 = (inp[1]) ? 3'b001 : 3'b011;
										assign node865 = (inp[2]) ? 3'b101 : 3'b001;
									assign node868 = (inp[8]) ? node874 : node869;
										assign node869 = (inp[2]) ? node871 : 3'b001;
											assign node871 = (inp[0]) ? 3'b110 : 3'b011;
										assign node874 = (inp[1]) ? node876 : 3'b110;
											assign node876 = (inp[0]) ? 3'b010 : 3'b110;
						assign node879 = (inp[10]) ? node881 : 3'b000;
							assign node881 = (inp[11]) ? node891 : node882;
								assign node882 = (inp[8]) ? 3'b000 : node883;
									assign node883 = (inp[0]) ? node885 : 3'b100;
										assign node885 = (inp[2]) ? node887 : 3'b100;
											assign node887 = (inp[5]) ? 3'b000 : 3'b100;
								assign node891 = (inp[5]) ? node903 : node892;
									assign node892 = (inp[2]) ? node898 : node893;
										assign node893 = (inp[8]) ? 3'b010 : node894;
											assign node894 = (inp[0]) ? 3'b010 : 3'b110;
										assign node898 = (inp[1]) ? node900 : 3'b110;
											assign node900 = (inp[0]) ? 3'b100 : 3'b110;
									assign node903 = (inp[8]) ? node909 : node904;
										assign node904 = (inp[0]) ? node906 : 3'b010;
											assign node906 = (inp[1]) ? 3'b100 : 3'b010;
										assign node909 = (inp[1]) ? node911 : 3'b100;
											assign node911 = (inp[2]) ? node913 : 3'b100;
												assign node913 = (inp[0]) ? 3'b000 : 3'b100;
					assign node916 = (inp[10]) ? node918 : 3'b000;
						assign node918 = (inp[7]) ? 3'b000 : node919;
							assign node919 = (inp[11]) ? node927 : node920;
								assign node920 = (inp[8]) ? 3'b000 : node921;
									assign node921 = (inp[0]) ? node923 : 3'b100;
										assign node923 = (inp[5]) ? 3'b000 : 3'b100;
								assign node927 = (inp[5]) ? node939 : node928;
									assign node928 = (inp[0]) ? node934 : node929;
										assign node929 = (inp[2]) ? 3'b110 : node930;
											assign node930 = (inp[8]) ? 3'b010 : 3'b110;
										assign node934 = (inp[8]) ? node936 : 3'b010;
											assign node936 = (inp[1]) ? 3'b100 : 3'b010;
									assign node939 = (inp[8]) ? node945 : node940;
										assign node940 = (inp[0]) ? node942 : 3'b010;
											assign node942 = (inp[1]) ? 3'b100 : 3'b010;
										assign node945 = (inp[0]) ? node947 : 3'b100;
											assign node947 = (inp[1]) ? node949 : 3'b100;
												assign node949 = (inp[2]) ? 3'b000 : 3'b100;
			assign node954 = (inp[3]) ? node1164 : node955;
				assign node955 = (inp[4]) ? node1053 : node956;
					assign node956 = (inp[7]) ? node988 : node957;
						assign node957 = (inp[10]) ? 3'b011 : node958;
							assign node958 = (inp[5]) ? node980 : node959;
								assign node959 = (inp[11]) ? node967 : node960;
									assign node960 = (inp[8]) ? node962 : 3'b001;
										assign node962 = (inp[1]) ? node964 : 3'b001;
											assign node964 = (inp[0]) ? 3'b011 : 3'b001;
									assign node967 = (inp[8]) ? node973 : node968;
										assign node968 = (inp[0]) ? node970 : 3'b001;
											assign node970 = (inp[2]) ? 3'b011 : 3'b001;
										assign node973 = (inp[1]) ? node975 : 3'b011;
											assign node975 = (inp[0]) ? node977 : 3'b011;
												assign node977 = (inp[2]) ? 3'b001 : 3'b011;
								assign node980 = (inp[11]) ? node982 : 3'b011;
									assign node982 = (inp[2]) ? 3'b001 : node983;
										assign node983 = (inp[8]) ? 3'b001 : 3'b011;
						assign node988 = (inp[10]) ? node1036 : node989;
							assign node989 = (inp[11]) ? node1013 : node990;
								assign node990 = (inp[5]) ? node1002 : node991;
									assign node991 = (inp[0]) ? node997 : node992;
										assign node992 = (inp[2]) ? 3'b010 : node993;
											assign node993 = (inp[8]) ? 3'b110 : 3'b010;
										assign node997 = (inp[2]) ? node999 : 3'b110;
											assign node999 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1002 = (inp[8]) ? node1008 : node1003;
										assign node1003 = (inp[1]) ? node1005 : 3'b110;
											assign node1005 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1008 = (inp[0]) ? node1010 : 3'b000;
											assign node1010 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1013 = (inp[5]) ? node1027 : node1014;
									assign node1014 = (inp[2]) ? node1020 : node1015;
										assign node1015 = (inp[8]) ? 3'b001 : node1016;
											assign node1016 = (inp[0]) ? 3'b011 : 3'b111;
										assign node1020 = (inp[8]) ? node1022 : 3'b111;
											assign node1022 = (inp[0]) ? node1024 : 3'b101;
												assign node1024 = (inp[1]) ? 3'b110 : 3'b101;
									assign node1027 = (inp[8]) ? 3'b110 : node1028;
										assign node1028 = (inp[0]) ? node1032 : node1029;
											assign node1029 = (inp[2]) ? 3'b011 : 3'b001;
											assign node1032 = (inp[2]) ? 3'b110 : 3'b100;
							assign node1036 = (inp[5]) ? node1044 : node1037;
								assign node1037 = (inp[11]) ? node1039 : 3'b001;
									assign node1039 = (inp[8]) ? node1041 : 3'b011;
										assign node1041 = (inp[1]) ? 3'b101 : 3'b011;
								assign node1044 = (inp[11]) ? node1048 : node1045;
									assign node1045 = (inp[8]) ? 3'b110 : 3'b111;
									assign node1048 = (inp[1]) ? node1050 : 3'b101;
										assign node1050 = (inp[8]) ? 3'b001 : 3'b101;
					assign node1053 = (inp[10]) ? node1091 : node1054;
						assign node1054 = (inp[7]) ? node1068 : node1055;
							assign node1055 = (inp[8]) ? node1059 : node1056;
								assign node1056 = (inp[11]) ? 3'b110 : 3'b010;
								assign node1059 = (inp[11]) ? node1061 : 3'b100;
									assign node1061 = (inp[1]) ? 3'b010 : node1062;
										assign node1062 = (inp[2]) ? 3'b110 : node1063;
											assign node1063 = (inp[0]) ? 3'b110 : 3'b101;
							assign node1068 = (inp[5]) ? node1082 : node1069;
								assign node1069 = (inp[8]) ? node1071 : 3'b010;
									assign node1071 = (inp[11]) ? node1077 : node1072;
										assign node1072 = (inp[0]) ? node1074 : 3'b010;
											assign node1074 = (inp[1]) ? 3'b000 : 3'b010;
										assign node1077 = (inp[1]) ? node1079 : 3'b110;
											assign node1079 = (inp[0]) ? 3'b100 : 3'b110;
								assign node1082 = (inp[11]) ? node1084 : 3'b000;
									assign node1084 = (inp[0]) ? node1088 : node1085;
										assign node1085 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1088 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1091 = (inp[7]) ? node1125 : node1092;
							assign node1092 = (inp[8]) ? node1110 : node1093;
								assign node1093 = (inp[11]) ? node1105 : node1094;
									assign node1094 = (inp[5]) ? node1100 : node1095;
										assign node1095 = (inp[2]) ? node1097 : 3'b101;
											assign node1097 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1100 = (inp[1]) ? 3'b001 : node1101;
											assign node1101 = (inp[0]) ? 3'b001 : 3'b101;
									assign node1105 = (inp[5]) ? node1107 : 3'b011;
										assign node1107 = (inp[0]) ? 3'b101 : 3'b011;
								assign node1110 = (inp[11]) ? node1120 : node1111;
									assign node1111 = (inp[2]) ? node1117 : node1112;
										assign node1112 = (inp[5]) ? node1114 : 3'b001;
											assign node1114 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1117 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1120 = (inp[0]) ? node1122 : 3'b101;
										assign node1122 = (inp[5]) ? 3'b001 : 3'b101;
							assign node1125 = (inp[11]) ? node1145 : node1126;
								assign node1126 = (inp[8]) ? node1132 : node1127;
									assign node1127 = (inp[0]) ? node1129 : 3'b110;
										assign node1129 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1132 = (inp[1]) ? node1138 : node1133;
										assign node1133 = (inp[5]) ? 3'b010 : node1134;
											assign node1134 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1138 = (inp[5]) ? node1142 : node1139;
											assign node1139 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1142 = (inp[2]) ? 3'b010 : 3'b100;
								assign node1145 = (inp[5]) ? node1153 : node1146;
									assign node1146 = (inp[0]) ? node1148 : 3'b001;
										assign node1148 = (inp[8]) ? node1150 : 3'b001;
											assign node1150 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1153 = (inp[8]) ? node1159 : node1154;
										assign node1154 = (inp[0]) ? node1156 : 3'b101;
											assign node1156 = (inp[1]) ? 3'b110 : 3'b101;
										assign node1159 = (inp[0]) ? node1161 : 3'b110;
											assign node1161 = (inp[1]) ? 3'b010 : 3'b110;
				assign node1164 = (inp[10]) ? node1204 : node1165;
					assign node1165 = (inp[4]) ? 3'b000 : node1166;
						assign node1166 = (inp[7]) ? 3'b000 : node1167;
							assign node1167 = (inp[11]) ? node1175 : node1168;
								assign node1168 = (inp[8]) ? 3'b000 : node1169;
									assign node1169 = (inp[5]) ? node1171 : 3'b100;
										assign node1171 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1175 = (inp[5]) ? node1191 : node1176;
									assign node1176 = (inp[2]) ? node1182 : node1177;
										assign node1177 = (inp[0]) ? 3'b010 : node1178;
											assign node1178 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1182 = (inp[8]) ? node1186 : node1183;
											assign node1183 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1186 = (inp[0]) ? node1188 : 3'b110;
												assign node1188 = (inp[1]) ? 3'b100 : 3'b110;
									assign node1191 = (inp[8]) ? node1197 : node1192;
										assign node1192 = (inp[1]) ? node1194 : 3'b010;
											assign node1194 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1197 = (inp[2]) ? node1199 : 3'b100;
											assign node1199 = (inp[1]) ? 3'b000 : 3'b100;
					assign node1204 = (inp[4]) ? node1296 : node1205;
						assign node1205 = (inp[7]) ? node1261 : node1206;
							assign node1206 = (inp[11]) ? node1226 : node1207;
								assign node1207 = (inp[8]) ? node1217 : node1208;
									assign node1208 = (inp[5]) ? node1212 : node1209;
										assign node1209 = (inp[0]) ? 3'b110 : 3'b010;
										assign node1212 = (inp[0]) ? node1214 : 3'b110;
											assign node1214 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1217 = (inp[5]) ? node1221 : node1218;
										assign node1218 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1221 = (inp[1]) ? node1223 : 3'b000;
											assign node1223 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1226 = (inp[5]) ? node1242 : node1227;
									assign node1227 = (inp[2]) ? node1233 : node1228;
										assign node1228 = (inp[8]) ? 3'b001 : node1229;
											assign node1229 = (inp[0]) ? 3'b011 : 3'b111;
										assign node1233 = (inp[0]) ? node1237 : node1234;
											assign node1234 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1237 = (inp[8]) ? node1239 : 3'b001;
												assign node1239 = (inp[1]) ? 3'b110 : 3'b101;
									assign node1242 = (inp[8]) ? node1254 : node1243;
										assign node1243 = (inp[2]) ? node1249 : node1244;
											assign node1244 = (inp[1]) ? node1246 : 3'b001;
												assign node1246 = (inp[0]) ? 3'b100 : 3'b001;
											assign node1249 = (inp[1]) ? node1251 : 3'b011;
												assign node1251 = (inp[0]) ? 3'b110 : 3'b011;
										assign node1254 = (inp[2]) ? node1256 : 3'b110;
											assign node1256 = (inp[1]) ? node1258 : 3'b110;
												assign node1258 = (inp[0]) ? 3'b010 : 3'b110;
							assign node1261 = (inp[11]) ? node1271 : node1262;
								assign node1262 = (inp[5]) ? 3'b000 : node1263;
									assign node1263 = (inp[0]) ? node1265 : 3'b100;
										assign node1265 = (inp[8]) ? node1267 : 3'b100;
											assign node1267 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1271 = (inp[5]) ? node1283 : node1272;
									assign node1272 = (inp[8]) ? node1278 : node1273;
										assign node1273 = (inp[2]) ? node1275 : 3'b110;
											assign node1275 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1278 = (inp[1]) ? node1280 : 3'b010;
											assign node1280 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1283 = (inp[8]) ? 3'b100 : node1284;
										assign node1284 = (inp[2]) ? node1290 : node1285;
											assign node1285 = (inp[1]) ? node1287 : 3'b010;
												assign node1287 = (inp[0]) ? 3'b000 : 3'b010;
											assign node1290 = (inp[0]) ? node1292 : 3'b110;
												assign node1292 = (inp[1]) ? 3'b100 : 3'b110;
						assign node1296 = (inp[7]) ? node1320 : node1297;
							assign node1297 = (inp[11]) ? node1305 : node1298;
								assign node1298 = (inp[8]) ? 3'b000 : node1299;
									assign node1299 = (inp[5]) ? node1301 : 3'b100;
										assign node1301 = (inp[2]) ? 3'b000 : 3'b100;
								assign node1305 = (inp[8]) ? node1315 : node1306;
									assign node1306 = (inp[0]) ? node1310 : node1307;
										assign node1307 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1310 = (inp[2]) ? 3'b010 : node1311;
											assign node1311 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1315 = (inp[5]) ? 3'b100 : node1316;
										assign node1316 = (inp[2]) ? 3'b100 : 3'b010;
							assign node1320 = (inp[11]) ? node1322 : 3'b000;
								assign node1322 = (inp[2]) ? 3'b000 : node1323;
									assign node1323 = (inp[8]) ? 3'b000 : node1324;
										assign node1324 = (inp[5]) ? 3'b000 : 3'b100;

endmodule