module dtc_split33_bm21 (
	input  wire [10-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node7;
	wire [10-1:0] node9;
	wire [10-1:0] node12;
	wire [10-1:0] node13;
	wire [10-1:0] node17;
	wire [10-1:0] node19;
	wire [10-1:0] node20;
	wire [10-1:0] node24;
	wire [10-1:0] node25;
	wire [10-1:0] node26;
	wire [10-1:0] node27;
	wire [10-1:0] node29;
	wire [10-1:0] node33;
	wire [10-1:0] node36;
	wire [10-1:0] node37;
	wire [10-1:0] node40;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node45;
	wire [10-1:0] node48;
	wire [10-1:0] node49;
	wire [10-1:0] node53;
	wire [10-1:0] node54;
	wire [10-1:0] node55;
	wire [10-1:0] node58;
	wire [10-1:0] node60;
	wire [10-1:0] node63;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node67;
	wire [10-1:0] node72;
	wire [10-1:0] node73;
	wire [10-1:0] node74;
	wire [10-1:0] node75;
	wire [10-1:0] node76;
	wire [10-1:0] node80;
	wire [10-1:0] node81;
	wire [10-1:0] node84;
	wire [10-1:0] node87;
	wire [10-1:0] node88;
	wire [10-1:0] node89;
	wire [10-1:0] node92;
	wire [10-1:0] node93;
	wire [10-1:0] node94;
	wire [10-1:0] node99;
	wire [10-1:0] node100;
	wire [10-1:0] node101;
	wire [10-1:0] node103;
	wire [10-1:0] node107;
	wire [10-1:0] node110;
	wire [10-1:0] node111;
	wire [10-1:0] node113;
	wire [10-1:0] node114;
	wire [10-1:0] node115;
	wire [10-1:0] node117;
	wire [10-1:0] node121;
	wire [10-1:0] node124;
	wire [10-1:0] node126;
	wire [10-1:0] node129;
	wire [10-1:0] node130;
	wire [10-1:0] node131;
	wire [10-1:0] node132;
	wire [10-1:0] node133;
	wire [10-1:0] node134;
	wire [10-1:0] node138;
	wire [10-1:0] node139;
	wire [10-1:0] node143;
	wire [10-1:0] node144;
	wire [10-1:0] node145;
	wire [10-1:0] node146;
	wire [10-1:0] node147;
	wire [10-1:0] node152;
	wire [10-1:0] node154;
	wire [10-1:0] node155;
	wire [10-1:0] node159;
	wire [10-1:0] node161;
	wire [10-1:0] node162;
	wire [10-1:0] node164;
	wire [10-1:0] node168;
	wire [10-1:0] node169;
	wire [10-1:0] node171;
	wire [10-1:0] node172;
	wire [10-1:0] node173;
	wire [10-1:0] node177;
	wire [10-1:0] node180;
	wire [10-1:0] node181;
	wire [10-1:0] node183;
	wire [10-1:0] node186;
	wire [10-1:0] node187;
	wire [10-1:0] node189;
	wire [10-1:0] node193;
	wire [10-1:0] node194;
	wire [10-1:0] node195;
	wire [10-1:0] node196;
	wire [10-1:0] node198;
	wire [10-1:0] node201;
	wire [10-1:0] node203;
	wire [10-1:0] node206;
	wire [10-1:0] node207;
	wire [10-1:0] node208;
	wire [10-1:0] node212;
	wire [10-1:0] node213;
	wire [10-1:0] node216;
	wire [10-1:0] node219;
	wire [10-1:0] node220;
	wire [10-1:0] node221;
	wire [10-1:0] node223;
	wire [10-1:0] node226;
	wire [10-1:0] node227;
	wire [10-1:0] node231;
	wire [10-1:0] node232;
	wire [10-1:0] node233;
	wire [10-1:0] node236;
	wire [10-1:0] node239;
	wire [10-1:0] node240;
	wire [10-1:0] node243;
	wire [10-1:0] node244;
	wire [10-1:0] node248;
	wire [10-1:0] node249;
	wire [10-1:0] node250;
	wire [10-1:0] node251;
	wire [10-1:0] node252;
	wire [10-1:0] node253;
	wire [10-1:0] node254;
	wire [10-1:0] node255;
	wire [10-1:0] node260;
	wire [10-1:0] node261;
	wire [10-1:0] node263;
	wire [10-1:0] node266;
	wire [10-1:0] node267;
	wire [10-1:0] node269;
	wire [10-1:0] node273;
	wire [10-1:0] node274;
	wire [10-1:0] node277;
	wire [10-1:0] node280;
	wire [10-1:0] node281;
	wire [10-1:0] node282;
	wire [10-1:0] node283;
	wire [10-1:0] node286;
	wire [10-1:0] node287;
	wire [10-1:0] node289;
	wire [10-1:0] node292;
	wire [10-1:0] node293;
	wire [10-1:0] node296;
	wire [10-1:0] node300;
	wire [10-1:0] node301;
	wire [10-1:0] node303;
	wire [10-1:0] node306;
	wire [10-1:0] node307;
	wire [10-1:0] node311;
	wire [10-1:0] node312;
	wire [10-1:0] node313;
	wire [10-1:0] node314;
	wire [10-1:0] node315;
	wire [10-1:0] node319;
	wire [10-1:0] node321;
	wire [10-1:0] node324;
	wire [10-1:0] node325;
	wire [10-1:0] node326;
	wire [10-1:0] node327;
	wire [10-1:0] node331;
	wire [10-1:0] node332;
	wire [10-1:0] node334;
	wire [10-1:0] node338;
	wire [10-1:0] node340;
	wire [10-1:0] node343;
	wire [10-1:0] node344;
	wire [10-1:0] node345;
	wire [10-1:0] node347;
	wire [10-1:0] node350;
	wire [10-1:0] node352;
	wire [10-1:0] node353;
	wire [10-1:0] node357;
	wire [10-1:0] node358;
	wire [10-1:0] node359;
	wire [10-1:0] node360;
	wire [10-1:0] node362;
	wire [10-1:0] node366;
	wire [10-1:0] node367;
	wire [10-1:0] node371;
	wire [10-1:0] node372;
	wire [10-1:0] node373;
	wire [10-1:0] node377;
	wire [10-1:0] node380;
	wire [10-1:0] node381;
	wire [10-1:0] node382;
	wire [10-1:0] node383;
	wire [10-1:0] node384;
	wire [10-1:0] node386;
	wire [10-1:0] node387;
	wire [10-1:0] node391;
	wire [10-1:0] node392;
	wire [10-1:0] node394;
	wire [10-1:0] node398;
	wire [10-1:0] node399;
	wire [10-1:0] node402;
	wire [10-1:0] node405;
	wire [10-1:0] node406;
	wire [10-1:0] node407;
	wire [10-1:0] node408;
	wire [10-1:0] node411;
	wire [10-1:0] node413;
	wire [10-1:0] node416;
	wire [10-1:0] node417;
	wire [10-1:0] node420;
	wire [10-1:0] node422;
	wire [10-1:0] node423;
	wire [10-1:0] node427;
	wire [10-1:0] node428;
	wire [10-1:0] node429;
	wire [10-1:0] node430;
	wire [10-1:0] node434;
	wire [10-1:0] node435;
	wire [10-1:0] node439;
	wire [10-1:0] node440;
	wire [10-1:0] node441;
	wire [10-1:0] node445;
	wire [10-1:0] node448;
	wire [10-1:0] node449;
	wire [10-1:0] node450;
	wire [10-1:0] node451;
	wire [10-1:0] node452;
	wire [10-1:0] node456;
	wire [10-1:0] node457;
	wire [10-1:0] node458;
	wire [10-1:0] node463;
	wire [10-1:0] node464;
	wire [10-1:0] node465;
	wire [10-1:0] node466;
	wire [10-1:0] node470;
	wire [10-1:0] node471;
	wire [10-1:0] node473;
	wire [10-1:0] node476;
	wire [10-1:0] node479;
	wire [10-1:0] node480;
	wire [10-1:0] node483;
	wire [10-1:0] node486;
	wire [10-1:0] node487;
	wire [10-1:0] node488;
	wire [10-1:0] node490;
	wire [10-1:0] node493;
	wire [10-1:0] node494;
	wire [10-1:0] node497;
	wire [10-1:0] node499;
	wire [10-1:0] node502;
	wire [10-1:0] node503;
	wire [10-1:0] node504;
	wire [10-1:0] node507;
	wire [10-1:0] node509;
	wire [10-1:0] node510;
	wire [10-1:0] node514;
	wire [10-1:0] node515;
	wire [10-1:0] node517;
	wire [10-1:0] node518;
	wire [10-1:0] node522;
	wire [10-1:0] node523;
	wire [10-1:0] node526;
	wire [10-1:0] node528;

	assign outp = (inp[2]) ? node248 : node1;
		assign node1 = (inp[4]) ? node129 : node2;
			assign node2 = (inp[7]) ? node72 : node3;
				assign node3 = (inp[1]) ? node43 : node4;
					assign node4 = (inp[8]) ? node24 : node5;
						assign node5 = (inp[5]) ? node17 : node6;
							assign node6 = (inp[9]) ? node12 : node7;
								assign node7 = (inp[3]) ? node9 : 10'b0111111111;
									assign node9 = (inp[6]) ? 10'b0011111111 : 10'b0111111111;
								assign node12 = (inp[3]) ? 10'b0011111111 : node13;
									assign node13 = (inp[6]) ? 10'b0011111111 : 10'b0111111111;
							assign node17 = (inp[9]) ? node19 : 10'b0011111111;
								assign node19 = (inp[0]) ? 10'b0001111111 : node20;
									assign node20 = (inp[6]) ? 10'b0001111111 : 10'b0011111111;
						assign node24 = (inp[0]) ? node36 : node25;
							assign node25 = (inp[3]) ? node33 : node26;
								assign node26 = (inp[9]) ? 10'b0001111111 : node27;
									assign node27 = (inp[6]) ? node29 : 10'b0111111111;
										assign node29 = (inp[5]) ? 10'b0001111111 : 10'b0011111111;
								assign node33 = (inp[5]) ? 10'b0000111111 : 10'b0001111111;
							assign node36 = (inp[6]) ? node40 : node37;
								assign node37 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
								assign node40 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
					assign node43 = (inp[6]) ? node53 : node44;
						assign node44 = (inp[8]) ? node48 : node45;
							assign node45 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
							assign node48 = (inp[0]) ? 10'b0000111111 : node49;
								assign node49 = (inp[5]) ? 10'b0000111111 : 10'b0001111111;
						assign node53 = (inp[8]) ? node63 : node54;
							assign node54 = (inp[0]) ? node58 : node55;
								assign node55 = (inp[5]) ? 10'b0000111111 : 10'b0001111111;
								assign node58 = (inp[9]) ? node60 : 10'b0000111111;
									assign node60 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
							assign node63 = (inp[3]) ? 10'b0000011111 : node64;
								assign node64 = (inp[5]) ? 10'b0000011111 : node65;
									assign node65 = (inp[9]) ? node67 : 10'b0000111111;
										assign node67 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
				assign node72 = (inp[9]) ? node110 : node73;
					assign node73 = (inp[8]) ? node87 : node74;
						assign node74 = (inp[6]) ? node80 : node75;
							assign node75 = (inp[5]) ? 10'b0001111111 : node76;
								assign node76 = (inp[1]) ? 10'b0001111111 : 10'b0011111111;
							assign node80 = (inp[3]) ? node84 : node81;
								assign node81 = (inp[1]) ? 10'b0000111111 : 10'b0001111111;
								assign node84 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
						assign node87 = (inp[3]) ? node99 : node88;
							assign node88 = (inp[1]) ? node92 : node89;
								assign node89 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
								assign node92 = (inp[0]) ? 10'b0000011111 : node93;
									assign node93 = (inp[6]) ? 10'b0000011111 : node94;
										assign node94 = (inp[5]) ? 10'b0000111111 : 10'b0001111111;
							assign node99 = (inp[5]) ? node107 : node100;
								assign node100 = (inp[1]) ? 10'b0000011111 : node101;
									assign node101 = (inp[0]) ? node103 : 10'b0000111111;
										assign node103 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
								assign node107 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
					assign node110 = (inp[0]) ? node124 : node111;
						assign node111 = (inp[5]) ? node113 : 10'b0000111111;
							assign node113 = (inp[1]) ? node121 : node114;
								assign node114 = (inp[6]) ? 10'b0000001111 : node115;
									assign node115 = (inp[8]) ? node117 : 10'b0000111111;
										assign node117 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
								assign node121 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
						assign node124 = (inp[1]) ? node126 : 10'b0000011111;
							assign node126 = (inp[3]) ? 10'b0000011111 : 10'b0000001111;
			assign node129 = (inp[5]) ? node193 : node130;
				assign node130 = (inp[3]) ? node168 : node131;
					assign node131 = (inp[8]) ? node143 : node132;
						assign node132 = (inp[6]) ? node138 : node133;
							assign node133 = (inp[0]) ? 10'b0001111111 : node134;
								assign node134 = (inp[9]) ? 10'b0011111111 : 10'b0111111111;
							assign node138 = (inp[9]) ? 10'b0000111111 : node139;
								assign node139 = (inp[0]) ? 10'b0000111111 : 10'b0001111111;
						assign node143 = (inp[6]) ? node159 : node144;
							assign node144 = (inp[0]) ? node152 : node145;
								assign node145 = (inp[7]) ? 10'b0000011111 : node146;
									assign node146 = (inp[1]) ? 10'b0001111111 : node147;
										assign node147 = (inp[9]) ? 10'b0001111111 : 10'b0011111111;
								assign node152 = (inp[1]) ? node154 : 10'b0000111111;
									assign node154 = (inp[9]) ? 10'b0000011111 : node155;
										assign node155 = (inp[7]) ? 10'b0000011111 : 10'b0000111111;
							assign node159 = (inp[7]) ? node161 : 10'b0000011111;
								assign node161 = (inp[1]) ? 10'b0000001111 : node162;
									assign node162 = (inp[9]) ? node164 : 10'b0000011111;
										assign node164 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
					assign node168 = (inp[0]) ? node180 : node169;
						assign node169 = (inp[1]) ? node171 : 10'b0000111111;
							assign node171 = (inp[6]) ? node177 : node172;
								assign node172 = (inp[9]) ? 10'b0000011111 : node173;
									assign node173 = (inp[7]) ? 10'b0000011111 : 10'b0000111111;
								assign node177 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
						assign node180 = (inp[9]) ? node186 : node181;
							assign node181 = (inp[8]) ? node183 : 10'b0000011111;
								assign node183 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
							assign node186 = (inp[7]) ? 10'b0000001111 : node187;
								assign node187 = (inp[6]) ? node189 : 10'b0000011111;
									assign node189 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
				assign node193 = (inp[9]) ? node219 : node194;
					assign node194 = (inp[3]) ? node206 : node195;
						assign node195 = (inp[1]) ? node201 : node196;
							assign node196 = (inp[8]) ? node198 : 10'b0000111111;
								assign node198 = (inp[0]) ? 10'b0000111111 : 10'b0000011111;
							assign node201 = (inp[6]) ? node203 : 10'b0000011111;
								assign node203 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
						assign node206 = (inp[6]) ? node212 : node207;
							assign node207 = (inp[8]) ? 10'b0000011111 : node208;
								assign node208 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
							assign node212 = (inp[1]) ? node216 : node213;
								assign node213 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
								assign node216 = (inp[0]) ? 10'b0000000111 : 10'b0000011111;
					assign node219 = (inp[1]) ? node231 : node220;
						assign node220 = (inp[8]) ? node226 : node221;
							assign node221 = (inp[7]) ? node223 : 10'b0000011111;
								assign node223 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
							assign node226 = (inp[0]) ? 10'b0000001111 : node227;
								assign node227 = (inp[3]) ? 10'b0000001111 : 10'b0000011111;
						assign node231 = (inp[0]) ? node239 : node232;
							assign node232 = (inp[8]) ? node236 : node233;
								assign node233 = (inp[3]) ? 10'b0000001111 : 10'b0000011111;
								assign node236 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
							assign node239 = (inp[7]) ? node243 : node240;
								assign node240 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
								assign node243 = (inp[6]) ? 10'b0000000001 : node244;
									assign node244 = (inp[8]) ? 10'b0000000011 : 10'b0000000111;
		assign node248 = (inp[1]) ? node380 : node249;
			assign node249 = (inp[5]) ? node311 : node250;
				assign node250 = (inp[7]) ? node280 : node251;
					assign node251 = (inp[9]) ? node273 : node252;
						assign node252 = (inp[0]) ? node260 : node253;
							assign node253 = (inp[3]) ? 10'b0001111111 : node254;
								assign node254 = (inp[4]) ? 10'b0011111111 : node255;
									assign node255 = (inp[8]) ? 10'b0011111111 : 10'b0111111111;
							assign node260 = (inp[4]) ? node266 : node261;
								assign node261 = (inp[3]) ? node263 : 10'b0001111111;
									assign node263 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
								assign node266 = (inp[3]) ? 10'b0000011111 : node267;
									assign node267 = (inp[6]) ? node269 : 10'b0000111111;
										assign node269 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
						assign node273 = (inp[0]) ? node277 : node274;
							assign node274 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
							assign node277 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
					assign node280 = (inp[3]) ? node300 : node281;
						assign node281 = (inp[0]) ? 10'b0000011111 : node282;
							assign node282 = (inp[6]) ? node286 : node283;
								assign node283 = (inp[8]) ? 10'b0000111111 : 10'b0001111111;
								assign node286 = (inp[4]) ? node292 : node287;
									assign node287 = (inp[9]) ? node289 : 10'b0000111111;
										assign node289 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
									assign node292 = (inp[9]) ? node296 : node293;
										assign node293 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
										assign node296 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
						assign node300 = (inp[8]) ? node306 : node301;
							assign node301 = (inp[9]) ? node303 : 10'b0000011111;
								assign node303 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
							assign node306 = (inp[0]) ? 10'b0000000111 : node307;
								assign node307 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
				assign node311 = (inp[4]) ? node343 : node312;
					assign node312 = (inp[0]) ? node324 : node313;
						assign node313 = (inp[8]) ? node319 : node314;
							assign node314 = (inp[6]) ? 10'b0000111111 : node315;
								assign node315 = (inp[7]) ? 10'b0000111111 : 10'b0011111111;
							assign node319 = (inp[7]) ? node321 : 10'b0000111111;
								assign node321 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
						assign node324 = (inp[7]) ? node338 : node325;
							assign node325 = (inp[8]) ? node331 : node326;
								assign node326 = (inp[6]) ? 10'b0000011111 : node327;
									assign node327 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
								assign node331 = (inp[3]) ? 10'b0000001111 : node332;
									assign node332 = (inp[6]) ? node334 : 10'b0000011111;
										assign node334 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
							assign node338 = (inp[8]) ? node340 : 10'b0000001111;
								assign node340 = (inp[6]) ? 10'b0000000011 : 10'b0000000111;
					assign node343 = (inp[6]) ? node357 : node344;
						assign node344 = (inp[8]) ? node350 : node345;
							assign node345 = (inp[0]) ? node347 : 10'b0000011111;
								assign node347 = (inp[3]) ? 10'b0000001111 : 10'b0000011111;
							assign node350 = (inp[7]) ? node352 : 10'b0000001111;
								assign node352 = (inp[3]) ? 10'b0000001111 : node353;
									assign node353 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
						assign node357 = (inp[3]) ? node371 : node358;
							assign node358 = (inp[9]) ? node366 : node359;
								assign node359 = (inp[7]) ? 10'b0000001111 : node360;
									assign node360 = (inp[8]) ? node362 : 10'b0000011111;
										assign node362 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
								assign node366 = (inp[7]) ? 10'b0000000111 : node367;
									assign node367 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
							assign node371 = (inp[0]) ? node377 : node372;
								assign node372 = (inp[8]) ? 10'b0000000111 : node373;
									assign node373 = (inp[7]) ? 10'b0000000111 : 10'b0000001111;
								assign node377 = (inp[8]) ? 10'b0000000001 : 10'b0000000011;
			assign node380 = (inp[3]) ? node448 : node381;
				assign node381 = (inp[7]) ? node405 : node382;
					assign node382 = (inp[5]) ? node398 : node383;
						assign node383 = (inp[4]) ? node391 : node384;
							assign node384 = (inp[6]) ? node386 : 10'b0001111111;
								assign node386 = (inp[8]) ? 10'b0000111111 : node387;
									assign node387 = (inp[0]) ? 10'b0000111111 : 10'b0001111111;
							assign node391 = (inp[9]) ? 10'b0000001111 : node392;
								assign node392 = (inp[6]) ? node394 : 10'b0000111111;
									assign node394 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
						assign node398 = (inp[0]) ? node402 : node399;
							assign node399 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
							assign node402 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
					assign node405 = (inp[6]) ? node427 : node406;
						assign node406 = (inp[0]) ? node416 : node407;
							assign node407 = (inp[5]) ? node411 : node408;
								assign node408 = (inp[4]) ? 10'b0000111111 : 10'b0000011111;
								assign node411 = (inp[4]) ? node413 : 10'b0000011111;
									assign node413 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
							assign node416 = (inp[5]) ? node420 : node417;
								assign node417 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
								assign node420 = (inp[9]) ? node422 : 10'b0000001111;
									assign node422 = (inp[4]) ? 10'b0000000111 : node423;
										assign node423 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
						assign node427 = (inp[8]) ? node439 : node428;
							assign node428 = (inp[9]) ? node434 : node429;
								assign node429 = (inp[0]) ? 10'b0000001111 : node430;
									assign node430 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
								assign node434 = (inp[5]) ? 10'b0000000111 : node435;
									assign node435 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
							assign node439 = (inp[0]) ? node445 : node440;
								assign node440 = (inp[9]) ? 10'b0000000111 : node441;
									assign node441 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
								assign node445 = (inp[5]) ? 10'b0000000001 : 10'b0000000111;
				assign node448 = (inp[0]) ? node486 : node449;
					assign node449 = (inp[6]) ? node463 : node450;
						assign node450 = (inp[8]) ? node456 : node451;
							assign node451 = (inp[4]) ? 10'b0000011111 : node452;
								assign node452 = (inp[7]) ? 10'b0000111111 : 10'b0000011111;
							assign node456 = (inp[4]) ? 10'b0000001111 : node457;
								assign node457 = (inp[9]) ? 10'b0000001111 : node458;
									assign node458 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
						assign node463 = (inp[8]) ? node479 : node464;
							assign node464 = (inp[9]) ? node470 : node465;
								assign node465 = (inp[5]) ? 10'b0000001111 : node466;
									assign node466 = (inp[4]) ? 10'b0000011111 : 10'b0000111111;
								assign node470 = (inp[5]) ? node476 : node471;
									assign node471 = (inp[4]) ? node473 : 10'b0000001111;
										assign node473 = (inp[7]) ? 10'b0000000111 : 10'b0000001111;
									assign node476 = (inp[7]) ? 10'b0000000011 : 10'b0000000111;
							assign node479 = (inp[7]) ? node483 : node480;
								assign node480 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
								assign node483 = (inp[4]) ? 10'b0000000011 : 10'b0000000111;
					assign node486 = (inp[9]) ? node502 : node487;
						assign node487 = (inp[8]) ? node493 : node488;
							assign node488 = (inp[5]) ? node490 : 10'b0000001111;
								assign node490 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
							assign node493 = (inp[4]) ? node497 : node494;
								assign node494 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
								assign node497 = (inp[7]) ? node499 : 10'b0000000111;
									assign node499 = (inp[5]) ? 10'b0000000011 : 10'b0000000111;
						assign node502 = (inp[5]) ? node514 : node503;
							assign node503 = (inp[7]) ? node507 : node504;
								assign node504 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
								assign node507 = (inp[4]) ? node509 : 10'b0000000111;
									assign node509 = (inp[6]) ? 10'b0000000011 : node510;
										assign node510 = (inp[8]) ? 10'b0000000011 : 10'b0000000111;
							assign node514 = (inp[6]) ? node522 : node515;
								assign node515 = (inp[4]) ? node517 : 10'b0000000111;
									assign node517 = (inp[7]) ? 10'b0000000011 : node518;
										assign node518 = (inp[8]) ? 10'b0000000011 : 10'b0000000111;
								assign node522 = (inp[8]) ? node526 : node523;
									assign node523 = (inp[7]) ? 10'b0000000001 : 10'b0000000011;
									assign node526 = (inp[7]) ? node528 : 10'b0000000001;
										assign node528 = (inp[4]) ? 10'b0000000000 : 10'b0000000001;

endmodule